module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40);
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    reg [485:0] src16;
    reg [485:0] src17;
    reg [485:0] src18;
    reg [485:0] src19;
    reg [485:0] src20;
    reg [485:0] src21;
    reg [485:0] src22;
    reg [485:0] src23;
    reg [485:0] src24;
    reg [485:0] src25;
    reg [485:0] src26;
    reg [485:0] src27;
    reg [485:0] src28;
    reg [485:0] src29;
    reg [485:0] src30;
    reg [485:0] src31;
    compressor_CLA486_32 compressor_CLA486_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40));
    initial begin
        src0 <= 486'h0;
        src1 <= 486'h0;
        src2 <= 486'h0;
        src3 <= 486'h0;
        src4 <= 486'h0;
        src5 <= 486'h0;
        src6 <= 486'h0;
        src7 <= 486'h0;
        src8 <= 486'h0;
        src9 <= 486'h0;
        src10 <= 486'h0;
        src11 <= 486'h0;
        src12 <= 486'h0;
        src13 <= 486'h0;
        src14 <= 486'h0;
        src15 <= 486'h0;
        src16 <= 486'h0;
        src17 <= 486'h0;
        src18 <= 486'h0;
        src19 <= 486'h0;
        src20 <= 486'h0;
        src21 <= 486'h0;
        src22 <= 486'h0;
        src23 <= 486'h0;
        src24 <= 486'h0;
        src25 <= 486'h0;
        src26 <= 486'h0;
        src27 <= 486'h0;
        src28 <= 486'h0;
        src29 <= 486'h0;
        src30 <= 486'h0;
        src31 <= 486'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA486_32(
    input [485:0]src0,
    input [485:0]src1,
    input [485:0]src2,
    input [485:0]src3,
    input [485:0]src4,
    input [485:0]src5,
    input [485:0]src6,
    input [485:0]src7,
    input [485:0]src8,
    input [485:0]src9,
    input [485:0]src10,
    input [485:0]src11,
    input [485:0]src12,
    input [485:0]src13,
    input [485:0]src14,
    input [485:0]src15,
    input [485:0]src16,
    input [485:0]src17,
    input [485:0]src18,
    input [485:0]src19,
    input [485:0]src20,
    input [485:0]src21,
    input [485:0]src22,
    input [485:0]src23,
    input [485:0]src24,
    input [485:0]src25,
    input [485:0]src26,
    input [485:0]src27,
    input [485:0]src28,
    input [485:0]src29,
    input [485:0]src30,
    input [485:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [0:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [0:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [0:0] comp_out39;
    wire [0:0] comp_out40;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], 1'h0, comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], 1'h0, comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], 1'h0}),
        .dst({dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [485:0] src0,
      input wire [485:0] src1,
      input wire [485:0] src2,
      input wire [485:0] src3,
      input wire [485:0] src4,
      input wire [485:0] src5,
      input wire [485:0] src6,
      input wire [485:0] src7,
      input wire [485:0] src8,
      input wire [485:0] src9,
      input wire [485:0] src10,
      input wire [485:0] src11,
      input wire [485:0] src12,
      input wire [485:0] src13,
      input wire [485:0] src14,
      input wire [485:0] src15,
      input wire [485:0] src16,
      input wire [485:0] src17,
      input wire [485:0] src18,
      input wire [485:0] src19,
      input wire [485:0] src20,
      input wire [485:0] src21,
      input wire [485:0] src22,
      input wire [485:0] src23,
      input wire [485:0] src24,
      input wire [485:0] src25,
      input wire [485:0] src26,
      input wire [485:0] src27,
      input wire [485:0] src28,
      input wire [485:0] src29,
      input wire [485:0] src30,
      input wire [485:0] src31,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [0:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [0:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [0:0] dst39,
      output wire [0:0] dst40);

   wire [485:0] stage0_0;
   wire [485:0] stage0_1;
   wire [485:0] stage0_2;
   wire [485:0] stage0_3;
   wire [485:0] stage0_4;
   wire [485:0] stage0_5;
   wire [485:0] stage0_6;
   wire [485:0] stage0_7;
   wire [485:0] stage0_8;
   wire [485:0] stage0_9;
   wire [485:0] stage0_10;
   wire [485:0] stage0_11;
   wire [485:0] stage0_12;
   wire [485:0] stage0_13;
   wire [485:0] stage0_14;
   wire [485:0] stage0_15;
   wire [485:0] stage0_16;
   wire [485:0] stage0_17;
   wire [485:0] stage0_18;
   wire [485:0] stage0_19;
   wire [485:0] stage0_20;
   wire [485:0] stage0_21;
   wire [485:0] stage0_22;
   wire [485:0] stage0_23;
   wire [485:0] stage0_24;
   wire [485:0] stage0_25;
   wire [485:0] stage0_26;
   wire [485:0] stage0_27;
   wire [485:0] stage0_28;
   wire [485:0] stage0_29;
   wire [485:0] stage0_30;
   wire [485:0] stage0_31;
   wire [126:0] stage1_0;
   wire [137:0] stage1_1;
   wire [227:0] stage1_2;
   wire [187:0] stage1_3;
   wire [225:0] stage1_4;
   wire [217:0] stage1_5;
   wire [246:0] stage1_6;
   wire [223:0] stage1_7;
   wire [205:0] stage1_8;
   wire [213:0] stage1_9;
   wire [187:0] stage1_10;
   wire [219:0] stage1_11;
   wire [281:0] stage1_12;
   wire [204:0] stage1_13;
   wire [296:0] stage1_14;
   wire [171:0] stage1_15;
   wire [264:0] stage1_16;
   wire [270:0] stage1_17;
   wire [200:0] stage1_18;
   wire [299:0] stage1_19;
   wire [188:0] stage1_20;
   wire [198:0] stage1_21;
   wire [250:0] stage1_22;
   wire [177:0] stage1_23;
   wire [211:0] stage1_24;
   wire [234:0] stage1_25;
   wire [214:0] stage1_26;
   wire [158:0] stage1_27;
   wire [251:0] stage1_28;
   wire [235:0] stage1_29;
   wire [171:0] stage1_30;
   wire [160:0] stage1_31;
   wire [150:0] stage1_32;
   wire [80:0] stage1_33;
   wire [21:0] stage2_0;
   wire [106:0] stage2_1;
   wire [50:0] stage2_2;
   wire [87:0] stage2_3;
   wire [90:0] stage2_4;
   wire [83:0] stage2_5;
   wire [93:0] stage2_6;
   wire [109:0] stage2_7;
   wire [107:0] stage2_8;
   wire [74:0] stage2_9;
   wire [88:0] stage2_10;
   wire [91:0] stage2_11;
   wire [102:0] stage2_12;
   wire [101:0] stage2_13;
   wire [138:0] stage2_14;
   wire [135:0] stage2_15;
   wire [103:0] stage2_16;
   wire [121:0] stage2_17;
   wire [81:0] stage2_18;
   wire [109:0] stage2_19;
   wire [127:0] stage2_20;
   wire [78:0] stage2_21;
   wire [78:0] stage2_22;
   wire [109:0] stage2_23;
   wire [99:0] stage2_24;
   wire [87:0] stage2_25;
   wire [98:0] stage2_26;
   wire [96:0] stage2_27;
   wire [74:0] stage2_28;
   wire [120:0] stage2_29;
   wire [129:0] stage2_30;
   wire [83:0] stage2_31;
   wire [64:0] stage2_32;
   wire [45:0] stage2_33;
   wire [35:0] stage2_34;
   wire [13:0] stage2_35;
   wire [7:0] stage3_0;
   wire [17:0] stage3_1;
   wire [31:0] stage3_2;
   wire [26:0] stage3_3;
   wire [43:0] stage3_4;
   wire [48:0] stage3_5;
   wire [42:0] stage3_6;
   wire [68:0] stage3_7;
   wire [37:0] stage3_8;
   wire [69:0] stage3_9;
   wire [28:0] stage3_10;
   wire [43:0] stage3_11;
   wire [41:0] stage3_12;
   wire [40:0] stage3_13;
   wire [50:0] stage3_14;
   wire [89:0] stage3_15;
   wire [61:0] stage3_16;
   wire [49:0] stage3_17;
   wire [49:0] stage3_18;
   wire [49:0] stage3_19;
   wire [45:0] stage3_20;
   wire [58:0] stage3_21;
   wire [46:0] stage3_22;
   wire [47:0] stage3_23;
   wire [40:0] stage3_24;
   wire [39:0] stage3_25;
   wire [31:0] stage3_26;
   wire [66:0] stage3_27;
   wire [42:0] stage3_28;
   wire [38:0] stage3_29;
   wire [59:0] stage3_30;
   wire [39:0] stage3_31;
   wire [35:0] stage3_32;
   wire [39:0] stage3_33;
   wire [21:0] stage3_34;
   wire [12:0] stage3_35;
   wire [6:0] stage3_36;
   wire [1:0] stage3_37;
   wire [2:0] stage4_0;
   wire [8:0] stage4_1;
   wire [8:0] stage4_2;
   wire [9:0] stage4_3;
   wire [16:0] stage4_4;
   wire [22:0] stage4_5;
   wire [20:0] stage4_6;
   wire [26:0] stage4_7;
   wire [22:0] stage4_8;
   wire [26:0] stage4_9;
   wire [28:0] stage4_10;
   wire [20:0] stage4_11;
   wire [13:0] stage4_12;
   wire [27:0] stage4_13;
   wire [12:0] stage4_14;
   wire [47:0] stage4_15;
   wire [28:0] stage4_16;
   wire [34:0] stage4_17;
   wire [18:0] stage4_18;
   wire [28:0] stage4_19;
   wire [25:0] stage4_20;
   wire [21:0] stage4_21;
   wire [22:0] stage4_22;
   wire [21:0] stage4_23;
   wire [30:0] stage4_24;
   wire [16:0] stage4_25;
   wire [23:0] stage4_26;
   wire [27:0] stage4_27;
   wire [17:0] stage4_28;
   wire [20:0] stage4_29;
   wire [22:0] stage4_30;
   wire [20:0] stage4_31;
   wire [18:0] stage4_32;
   wire [13:0] stage4_33;
   wire [16:0] stage4_34;
   wire [13:0] stage4_35;
   wire [9:0] stage4_36;
   wire [1:0] stage4_37;
   wire [0:0] stage4_38;
   wire [2:0] stage5_0;
   wire [8:0] stage5_1;
   wire [4:0] stage5_2;
   wire [7:0] stage5_3;
   wire [3:0] stage5_4;
   wire [8:0] stage5_5;
   wire [9:0] stage5_6;
   wire [10:0] stage5_7;
   wire [12:0] stage5_8;
   wire [11:0] stage5_9;
   wire [22:0] stage5_10;
   wire [8:0] stage5_11;
   wire [10:0] stage5_12;
   wire [15:0] stage5_13;
   wire [7:0] stage5_14;
   wire [10:0] stage5_15;
   wire [21:0] stage5_16;
   wire [14:0] stage5_17;
   wire [12:0] stage5_18;
   wire [12:0] stage5_19;
   wire [9:0] stage5_20;
   wire [10:0] stage5_21;
   wire [11:0] stage5_22;
   wire [13:0] stage5_23;
   wire [7:0] stage5_24;
   wire [7:0] stage5_25;
   wire [13:0] stage5_26;
   wire [13:0] stage5_27;
   wire [6:0] stage5_28;
   wire [12:0] stage5_29;
   wire [11:0] stage5_30;
   wire [10:0] stage5_31;
   wire [10:0] stage5_32;
   wire [8:0] stage5_33;
   wire [7:0] stage5_34;
   wire [14:0] stage5_35;
   wire [3:0] stage5_36;
   wire [5:0] stage5_37;
   wire [1:0] stage5_38;
   wire [2:0] stage6_0;
   wire [6:0] stage6_1;
   wire [0:0] stage6_2;
   wire [3:0] stage6_3;
   wire [1:0] stage6_4;
   wire [5:0] stage6_5;
   wire [4:0] stage6_6;
   wire [2:0] stage6_7;
   wire [5:0] stage6_8;
   wire [4:0] stage6_9;
   wire [6:0] stage6_10;
   wire [5:0] stage6_11;
   wire [6:0] stage6_12;
   wire [8:0] stage6_13;
   wire [5:0] stage6_14;
   wire [5:0] stage6_15;
   wire [4:0] stage6_16;
   wire [9:0] stage6_17;
   wire [5:0] stage6_18;
   wire [4:0] stage6_19;
   wire [5:0] stage6_20;
   wire [5:0] stage6_21;
   wire [4:0] stage6_22;
   wire [8:0] stage6_23;
   wire [3:0] stage6_24;
   wire [4:0] stage6_25;
   wire [11:0] stage6_26;
   wire [8:0] stage6_27;
   wire [6:0] stage6_28;
   wire [3:0] stage6_29;
   wire [4:0] stage6_30;
   wire [7:0] stage6_31;
   wire [3:0] stage6_32;
   wire [5:0] stage6_33;
   wire [10:0] stage6_34;
   wire [4:0] stage6_35;
   wire [5:0] stage6_36;
   wire [1:0] stage6_37;
   wire [2:0] stage6_38;
   wire [0:0] stage6_39;
   wire [2:0] stage7_0;
   wire [6:0] stage7_1;
   wire [0:0] stage7_2;
   wire [3:0] stage7_3;
   wire [1:0] stage7_4;
   wire [3:0] stage7_5;
   wire [3:0] stage7_6;
   wire [1:0] stage7_7;
   wire [6:0] stage7_8;
   wire [0:0] stage7_9;
   wire [4:0] stage7_10;
   wire [1:0] stage7_11;
   wire [3:0] stage7_12;
   wire [1:0] stage7_13;
   wire [6:0] stage7_14;
   wire [5:0] stage7_15;
   wire [1:0] stage7_16;
   wire [3:0] stage7_17;
   wire [1:0] stage7_18;
   wire [2:0] stage7_19;
   wire [6:0] stage7_20;
   wire [0:0] stage7_21;
   wire [5:0] stage7_22;
   wire [5:0] stage7_23;
   wire [3:0] stage7_24;
   wire [0:0] stage7_25;
   wire [2:0] stage7_26;
   wire [5:0] stage7_27;
   wire [5:0] stage7_28;
   wire [3:0] stage7_29;
   wire [2:0] stage7_30;
   wire [1:0] stage7_31;
   wire [5:0] stage7_32;
   wire [1:0] stage7_33;
   wire [6:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [3:0] stage7_37;
   wire [3:0] stage7_38;
   wire [0:0] stage7_39;
   wire [0:0] stage8_0;
   wire [1:0] stage8_1;
   wire [0:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [0:0] stage8_5;
   wire [1:0] stage8_6;
   wire [1:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [0:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [1:0] stage8_24;
   wire [1:0] stage8_25;
   wire [1:0] stage8_26;
   wire [1:0] stage8_27;
   wire [1:0] stage8_28;
   wire [1:0] stage8_29;
   wire [1:0] stage8_30;
   wire [1:0] stage8_31;
   wire [1:0] stage8_32;
   wire [1:0] stage8_33;
   wire [1:0] stage8_34;
   wire [1:0] stage8_35;
   wire [1:0] stage8_36;
   wire [1:0] stage8_37;
   wire [1:0] stage8_38;
   wire [0:0] stage8_39;
   wire [0:0] stage8_40;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;
   assign dst25 = stage8_25;
   assign dst26 = stage8_26;
   assign dst27 = stage8_27;
   assign dst28 = stage8_28;
   assign dst29 = stage8_29;
   assign dst30 = stage8_30;
   assign dst31 = stage8_31;
   assign dst32 = stage8_32;
   assign dst33 = stage8_33;
   assign dst34 = stage8_34;
   assign dst35 = stage8_35;
   assign dst36 = stage8_36;
   assign dst37 = stage8_37;
   assign dst38 = stage8_38;
   assign dst39 = stage8_39;
   assign dst40 = stage8_40;

   gpc1343_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3]},
      {stage0_2[0], stage0_2[1], stage0_2[2]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[4]},
      {stage0_2[3]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_1[5]},
      {stage0_2[4]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_1[6]},
      {stage0_2[5]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30]},
      {stage0_1[7]},
      {stage0_2[6]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc117_4 gpc5 (
      {stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_1[8]},
      {stage0_2[7]},
      {stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc117_4 gpc6 (
      {stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[9]},
      {stage0_2[8]},
      {stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc117_4 gpc7 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51]},
      {stage0_1[10]},
      {stage0_2[9]},
      {stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc117_4 gpc8 (
      {stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58]},
      {stage0_1[11]},
      {stage0_2[10]},
      {stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc117_4 gpc9 (
      {stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63], stage0_0[64], stage0_0[65]},
      {stage0_1[12]},
      {stage0_2[11]},
      {stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc117_4 gpc10 (
      {stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72]},
      {stage0_1[13]},
      {stage0_2[12]},
      {stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc117_4 gpc11 (
      {stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79]},
      {stage0_1[14]},
      {stage0_2[13]},
      {stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc117_4 gpc12 (
      {stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_1[15]},
      {stage0_2[14]},
      {stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc117_4 gpc13 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_1[16]},
      {stage0_2[15]},
      {stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc117_4 gpc14 (
      {stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100]},
      {stage0_1[17]},
      {stage0_2[16]},
      {stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc117_4 gpc15 (
      {stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107]},
      {stage0_1[18]},
      {stage0_2[17]},
      {stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc117_4 gpc16 (
      {stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[19]},
      {stage0_2[18]},
      {stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_2[19]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_2[20]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37]},
      {stage0_2[21]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43]},
      {stage0_2[22]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49]},
      {stage0_2[23]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55]},
      {stage0_2[24]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61]},
      {stage0_2[25]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67]},
      {stage0_2[26]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73]},
      {stage0_2[27]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79]},
      {stage0_2[28]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85]},
      {stage0_2[29]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[148], stage0_0[149], stage0_0[150]},
      {stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91]},
      {stage0_2[30]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97]},
      {stage0_2[31]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103]},
      {stage0_2[32]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109]},
      {stage0_2[33]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[160], stage0_0[161], stage0_0[162]},
      {stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115]},
      {stage0_2[34]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121]},
      {stage0_2[35]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[166], stage0_0[167], stage0_0[168]},
      {stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127]},
      {stage0_2[36]},
      {stage0_3[18]},
      {stage1_4[18],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133]},
      {stage0_2[37]},
      {stage0_3[19]},
      {stage1_4[19],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[172], stage0_0[173], stage0_0[174]},
      {stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139]},
      {stage0_2[38]},
      {stage0_3[20]},
      {stage1_4[20],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145]},
      {stage0_2[39]},
      {stage0_3[21]},
      {stage1_4[21],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[178], stage0_0[179], stage0_0[180]},
      {stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151]},
      {stage0_2[40]},
      {stage0_3[22]},
      {stage1_4[22],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157]},
      {stage0_2[41]},
      {stage0_3[23]},
      {stage1_4[23],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[184], stage0_0[185], stage0_0[186]},
      {stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163]},
      {stage0_2[42]},
      {stage0_3[24]},
      {stage1_4[24],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169]},
      {stage0_2[43]},
      {stage0_3[25]},
      {stage1_4[25],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc1163_5 gpc42 (
      {stage0_0[190], stage0_0[191], stage0_0[192]},
      {stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175]},
      {stage0_2[44]},
      {stage0_3[26]},
      {stage1_4[26],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[193], stage0_0[194], stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[27],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[28],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[29],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[30],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[31],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226], stage0_0[227], stage0_0[228]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[32],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232], stage0_0[233], stage0_0[234]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[33],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[235], stage0_0[236], stage0_0[237], stage0_0[238], stage0_0[239], stage0_0[240]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[34],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[241], stage0_0[242], stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[35],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[247], stage0_0[248], stage0_0[249], stage0_0[250], stage0_0[251], stage0_0[252]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[36],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[253], stage0_0[254], stage0_0[255], stage0_0[256], stage0_0[257], stage0_0[258]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[37],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[259], stage0_0[260], stage0_0[261], stage0_0[262], stage0_0[263], stage0_0[264]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[38],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[265], stage0_0[266], stage0_0[267], stage0_0[268], stage0_0[269], stage0_0[270]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[39],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[271], stage0_0[272], stage0_0[273], stage0_0[274], stage0_0[275], stage0_0[276]},
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128]},
      {stage1_4[40],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[277], stage0_0[278], stage0_0[279], stage0_0[280], stage0_0[281], stage0_0[282]},
      {stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage1_4[41],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[283], stage0_0[284], stage0_0[285], stage0_0[286], stage0_0[287], stage0_0[288]},
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140]},
      {stage1_4[42],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[289], stage0_0[290], stage0_0[291], stage0_0[292], stage0_0[293], stage0_0[294]},
      {stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage1_4[43],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[295], stage0_0[296], stage0_0[297], stage0_0[298], stage0_0[299], stage0_0[300]},
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152]},
      {stage1_4[44],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[301], stage0_0[302], stage0_0[303], stage0_0[304], stage0_0[305], stage0_0[306]},
      {stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage1_4[45],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[307], stage0_0[308], stage0_0[309], stage0_0[310], stage0_0[311], stage0_0[312]},
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164]},
      {stage1_4[46],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[313], stage0_0[314], stage0_0[315], stage0_0[316], stage0_0[317], stage0_0[318]},
      {stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage1_4[47],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[319], stage0_0[320], stage0_0[321], stage0_0[322], stage0_0[323], stage0_0[324]},
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176]},
      {stage1_4[48],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[325], stage0_0[326], stage0_0[327], stage0_0[328], stage0_0[329], stage0_0[330]},
      {stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage1_4[49],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[331], stage0_0[332], stage0_0[333], stage0_0[334], stage0_0[335], stage0_0[336]},
      {stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage1_4[50],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[337], stage0_0[338], stage0_0[339], stage0_0[340], stage0_0[341], stage0_0[342]},
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194]},
      {stage1_4[51],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[343], stage0_0[344], stage0_0[345], stage0_0[346], stage0_0[347], stage0_0[348]},
      {stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage1_4[52],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[349], stage0_0[350], stage0_0[351], stage0_0[352], stage0_0[353], stage0_0[354]},
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205], stage0_2[206]},
      {stage1_4[53],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[355], stage0_0[356], stage0_0[357], stage0_0[358], stage0_0[359], stage0_0[360]},
      {stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210], stage0_2[211], stage0_2[212]},
      {stage1_4[54],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[361], stage0_0[362], stage0_0[363], stage0_0[364], stage0_0[365], stage0_0[366]},
      {stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216], stage0_2[217], stage0_2[218]},
      {stage1_4[55],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[367], stage0_0[368], stage0_0[369], stage0_0[370], stage0_0[371], stage0_0[372]},
      {stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224]},
      {stage1_4[56],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[373], stage0_0[374], stage0_0[375], stage0_0[376], stage0_0[377], stage0_0[378]},
      {stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage1_4[57],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[379], stage0_0[380], stage0_0[381], stage0_0[382], stage0_0[383], stage0_0[384]},
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235], stage0_2[236]},
      {stage1_4[58],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[385], stage0_0[386], stage0_0[387], stage0_0[388], stage0_0[389], stage0_0[390]},
      {stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240], stage0_2[241], stage0_2[242]},
      {stage1_4[59],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[391], stage0_0[392], stage0_0[393], stage0_0[394], stage0_0[395], stage0_0[396]},
      {stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246], stage0_2[247], stage0_2[248]},
      {stage1_4[60],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[397], stage0_0[398], stage0_0[399], stage0_0[400], stage0_0[401], stage0_0[402]},
      {stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252], stage0_2[253], stage0_2[254]},
      {stage1_4[61],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[403], stage0_0[404], stage0_0[405], stage0_0[406], stage0_0[407], stage0_0[408]},
      {stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258], stage0_2[259], stage0_2[260]},
      {stage1_4[62],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[409], stage0_0[410], stage0_0[411], stage0_0[412], stage0_0[413], stage0_0[414]},
      {stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264], stage0_2[265], stage0_2[266]},
      {stage1_4[63],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[415], stage0_0[416], stage0_0[417], stage0_0[418], stage0_0[419], stage0_0[420]},
      {stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270], stage0_2[271], stage0_2[272]},
      {stage1_4[64],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[421], stage0_0[422], stage0_0[423], stage0_0[424], stage0_0[425], stage0_0[426]},
      {stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276], stage0_2[277], stage0_2[278]},
      {stage1_4[65],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[427], stage0_0[428], stage0_0[429], stage0_0[430], stage0_0[431], stage0_0[432]},
      {stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282], stage0_2[283], stage0_2[284]},
      {stage1_4[66],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[433], stage0_0[434], stage0_0[435], stage0_0[436], stage0_0[437], stage0_0[438]},
      {stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288], stage0_2[289], stage0_2[290]},
      {stage1_4[67],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc1325_5 gpc84 (
      {stage0_0[439], stage0_0[440], stage0_0[441], stage0_0[442], stage0_0[443]},
      {stage0_1[176], stage0_1[177]},
      {stage0_2[291], stage0_2[292], stage0_2[293]},
      {stage0_3[27]},
      {stage1_4[68],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183]},
      {stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33]},
      {stage1_5[0],stage1_4[69],stage1_3[85],stage1_2[85],stage1_1[85]}
   );
   gpc606_5 gpc86 (
      {stage0_1[184], stage0_1[185], stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189]},
      {stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage1_5[1],stage1_4[70],stage1_3[86],stage1_2[86],stage1_1[86]}
   );
   gpc606_5 gpc87 (
      {stage0_1[190], stage0_1[191], stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195]},
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45]},
      {stage1_5[2],stage1_4[71],stage1_3[87],stage1_2[87],stage1_1[87]}
   );
   gpc606_5 gpc88 (
      {stage0_1[196], stage0_1[197], stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201]},
      {stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage1_5[3],stage1_4[72],stage1_3[88],stage1_2[88],stage1_1[88]}
   );
   gpc606_5 gpc89 (
      {stage0_1[202], stage0_1[203], stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207]},
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57]},
      {stage1_5[4],stage1_4[73],stage1_3[89],stage1_2[89],stage1_1[89]}
   );
   gpc606_5 gpc90 (
      {stage0_1[208], stage0_1[209], stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213]},
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage1_5[5],stage1_4[74],stage1_3[90],stage1_2[90],stage1_1[90]}
   );
   gpc606_5 gpc91 (
      {stage0_1[214], stage0_1[215], stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219]},
      {stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69]},
      {stage1_5[6],stage1_4[75],stage1_3[91],stage1_2[91],stage1_1[91]}
   );
   gpc606_5 gpc92 (
      {stage0_1[220], stage0_1[221], stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225]},
      {stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75]},
      {stage1_5[7],stage1_4[76],stage1_3[92],stage1_2[92],stage1_1[92]}
   );
   gpc606_5 gpc93 (
      {stage0_1[226], stage0_1[227], stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231]},
      {stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81]},
      {stage1_5[8],stage1_4[77],stage1_3[93],stage1_2[93],stage1_1[93]}
   );
   gpc606_5 gpc94 (
      {stage0_1[232], stage0_1[233], stage0_1[234], stage0_1[235], stage0_1[236], stage0_1[237]},
      {stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87]},
      {stage1_5[9],stage1_4[78],stage1_3[94],stage1_2[94],stage1_1[94]}
   );
   gpc606_5 gpc95 (
      {stage0_1[238], stage0_1[239], stage0_1[240], stage0_1[241], stage0_1[242], stage0_1[243]},
      {stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93]},
      {stage1_5[10],stage1_4[79],stage1_3[95],stage1_2[95],stage1_1[95]}
   );
   gpc606_5 gpc96 (
      {stage0_1[244], stage0_1[245], stage0_1[246], stage0_1[247], stage0_1[248], stage0_1[249]},
      {stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage1_5[11],stage1_4[80],stage1_3[96],stage1_2[96],stage1_1[96]}
   );
   gpc606_5 gpc97 (
      {stage0_1[250], stage0_1[251], stage0_1[252], stage0_1[253], stage0_1[254], stage0_1[255]},
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105]},
      {stage1_5[12],stage1_4[81],stage1_3[97],stage1_2[97],stage1_1[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[256], stage0_1[257], stage0_1[258], stage0_1[259], stage0_1[260], stage0_1[261]},
      {stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage1_5[13],stage1_4[82],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[262], stage0_1[263], stage0_1[264], stage0_1[265], stage0_1[266], stage0_1[267]},
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117]},
      {stage1_5[14],stage1_4[83],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[268], stage0_1[269], stage0_1[270], stage0_1[271], stage0_1[272], stage0_1[273]},
      {stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage1_5[15],stage1_4[84],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[274], stage0_1[275], stage0_1[276], stage0_1[277], stage0_1[278], stage0_1[279]},
      {stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129]},
      {stage1_5[16],stage1_4[85],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[280], stage0_1[281], stage0_1[282], stage0_1[283], stage0_1[284], stage0_1[285]},
      {stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134], stage0_3[135]},
      {stage1_5[17],stage1_4[86],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[286], stage0_1[287], stage0_1[288], stage0_1[289], stage0_1[290], stage0_1[291]},
      {stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140], stage0_3[141]},
      {stage1_5[18],stage1_4[87],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[292], stage0_1[293], stage0_1[294], stage0_1[295], stage0_1[296], stage0_1[297]},
      {stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146], stage0_3[147]},
      {stage1_5[19],stage1_4[88],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[298], stage0_1[299], stage0_1[300], stage0_1[301], stage0_1[302], stage0_1[303]},
      {stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153]},
      {stage1_5[20],stage1_4[89],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[304], stage0_1[305], stage0_1[306], stage0_1[307], stage0_1[308], stage0_1[309]},
      {stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159]},
      {stage1_5[21],stage1_4[90],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[310], stage0_1[311], stage0_1[312], stage0_1[313], stage0_1[314], stage0_1[315]},
      {stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165]},
      {stage1_5[22],stage1_4[91],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[316], stage0_1[317], stage0_1[318], stage0_1[319], stage0_1[320], stage0_1[321]},
      {stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170], stage0_3[171]},
      {stage1_5[23],stage1_4[92],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[322], stage0_1[323], stage0_1[324], stage0_1[325], stage0_1[326], stage0_1[327]},
      {stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176], stage0_3[177]},
      {stage1_5[24],stage1_4[93],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[328], stage0_1[329], stage0_1[330], stage0_1[331], stage0_1[332], stage0_1[333]},
      {stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182], stage0_3[183]},
      {stage1_5[25],stage1_4[94],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[334], stage0_1[335], stage0_1[336], stage0_1[337], stage0_1[338], stage0_1[339]},
      {stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188], stage0_3[189]},
      {stage1_5[26],stage1_4[95],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[340], stage0_1[341], stage0_1[342], stage0_1[343], stage0_1[344], stage0_1[345]},
      {stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195]},
      {stage1_5[27],stage1_4[96],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[346], stage0_1[347], stage0_1[348], stage0_1[349], stage0_1[350], stage0_1[351]},
      {stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201]},
      {stage1_5[28],stage1_4[97],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[352], stage0_1[353], stage0_1[354], stage0_1[355], stage0_1[356], stage0_1[357]},
      {stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206], stage0_3[207]},
      {stage1_5[29],stage1_4[98],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[358], stage0_1[359], stage0_1[360], stage0_1[361], stage0_1[362], stage0_1[363]},
      {stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212], stage0_3[213]},
      {stage1_5[30],stage1_4[99],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[364], stage0_1[365], stage0_1[366], stage0_1[367], stage0_1[368], stage0_1[369]},
      {stage0_3[214], stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218], stage0_3[219]},
      {stage1_5[31],stage1_4[100],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[370], stage0_1[371], stage0_1[372], stage0_1[373], stage0_1[374], stage0_1[375]},
      {stage0_3[220], stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225]},
      {stage1_5[32],stage1_4[101],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[376], stage0_1[377], stage0_1[378], stage0_1[379], stage0_1[380], stage0_1[381]},
      {stage0_3[226], stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231]},
      {stage1_5[33],stage1_4[102],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[382], stage0_1[383], stage0_1[384], stage0_1[385], stage0_1[386], stage0_1[387]},
      {stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236], stage0_3[237]},
      {stage1_5[34],stage1_4[103],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[388], stage0_1[389], stage0_1[390], stage0_1[391], stage0_1[392], stage0_1[393]},
      {stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242], stage0_3[243]},
      {stage1_5[35],stage1_4[104],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[394], stage0_1[395], stage0_1[396], stage0_1[397], stage0_1[398], stage0_1[399]},
      {stage0_3[244], stage0_3[245], stage0_3[246], stage0_3[247], stage0_3[248], stage0_3[249]},
      {stage1_5[36],stage1_4[105],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[400], stage0_1[401], stage0_1[402], stage0_1[403], stage0_1[404], stage0_1[405]},
      {stage0_3[250], stage0_3[251], stage0_3[252], stage0_3[253], stage0_3[254], stage0_3[255]},
      {stage1_5[37],stage1_4[106],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[406], stage0_1[407], stage0_1[408], stage0_1[409], stage0_1[410], stage0_1[411]},
      {stage0_3[256], stage0_3[257], stage0_3[258], stage0_3[259], stage0_3[260], stage0_3[261]},
      {stage1_5[38],stage1_4[107],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[412], stage0_1[413], stage0_1[414], stage0_1[415], stage0_1[416], stage0_1[417]},
      {stage0_3[262], stage0_3[263], stage0_3[264], stage0_3[265], stage0_3[266], stage0_3[267]},
      {stage1_5[39],stage1_4[108],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[418], stage0_1[419], stage0_1[420], stage0_1[421], stage0_1[422], stage0_1[423]},
      {stage0_3[268], stage0_3[269], stage0_3[270], stage0_3[271], stage0_3[272], stage0_3[273]},
      {stage1_5[40],stage1_4[109],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[424], stage0_1[425], stage0_1[426], stage0_1[427], stage0_1[428], stage0_1[429]},
      {stage0_3[274], stage0_3[275], stage0_3[276], stage0_3[277], stage0_3[278], stage0_3[279]},
      {stage1_5[41],stage1_4[110],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[430], stage0_1[431], stage0_1[432], stage0_1[433], stage0_1[434], stage0_1[435]},
      {stage0_3[280], stage0_3[281], stage0_3[282], stage0_3[283], stage0_3[284], stage0_3[285]},
      {stage1_5[42],stage1_4[111],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[436], stage0_1[437], stage0_1[438], stage0_1[439], stage0_1[440], stage0_1[441]},
      {stage0_3[286], stage0_3[287], stage0_3[288], stage0_3[289], stage0_3[290], stage0_3[291]},
      {stage1_5[43],stage1_4[112],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[442], stage0_1[443], stage0_1[444], stage0_1[445], stage0_1[446], stage0_1[447]},
      {stage0_3[292], stage0_3[293], stage0_3[294], stage0_3[295], stage0_3[296], stage0_3[297]},
      {stage1_5[44],stage1_4[113],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[448], stage0_1[449], stage0_1[450], stage0_1[451], stage0_1[452], stage0_1[453]},
      {stage0_3[298], stage0_3[299], stage0_3[300], stage0_3[301], stage0_3[302], stage0_3[303]},
      {stage1_5[45],stage1_4[114],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[454], stage0_1[455], stage0_1[456], stage0_1[457], stage0_1[458], stage0_1[459]},
      {stage0_3[304], stage0_3[305], stage0_3[306], stage0_3[307], stage0_3[308], stage0_3[309]},
      {stage1_5[46],stage1_4[115],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[460], stage0_1[461], stage0_1[462], stage0_1[463], stage0_1[464], stage0_1[465]},
      {stage0_3[310], stage0_3[311], stage0_3[312], stage0_3[313], stage0_3[314], stage0_3[315]},
      {stage1_5[47],stage1_4[116],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[466], stage0_1[467], stage0_1[468], stage0_1[469], stage0_1[470], stage0_1[471]},
      {stage0_3[316], stage0_3[317], stage0_3[318], stage0_3[319], stage0_3[320], stage0_3[321]},
      {stage1_5[48],stage1_4[117],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[472], stage0_1[473], stage0_1[474], stage0_1[475], stage0_1[476], stage0_1[477]},
      {stage0_3[322], stage0_3[323], stage0_3[324], stage0_3[325], stage0_3[326], stage0_3[327]},
      {stage1_5[49],stage1_4[118],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[478], stage0_1[479], stage0_1[480], stage0_1[481], stage0_1[482], stage0_1[483]},
      {stage0_3[328], stage0_3[329], stage0_3[330], stage0_3[331], stage0_3[332], stage0_3[333]},
      {stage1_5[50],stage1_4[119],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_2[294], stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[51],stage1_4[120],stage1_3[136],stage1_2[136]}
   );
   gpc606_5 gpc137 (
      {stage0_2[300], stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[52],stage1_4[121],stage1_3[137],stage1_2[137]}
   );
   gpc606_5 gpc138 (
      {stage0_2[306], stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[53],stage1_4[122],stage1_3[138],stage1_2[138]}
   );
   gpc606_5 gpc139 (
      {stage0_2[312], stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[54],stage1_4[123],stage1_3[139],stage1_2[139]}
   );
   gpc606_5 gpc140 (
      {stage0_2[318], stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[55],stage1_4[124],stage1_3[140],stage1_2[140]}
   );
   gpc606_5 gpc141 (
      {stage0_2[324], stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[56],stage1_4[125],stage1_3[141],stage1_2[141]}
   );
   gpc606_5 gpc142 (
      {stage0_2[330], stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[57],stage1_4[126],stage1_3[142],stage1_2[142]}
   );
   gpc606_5 gpc143 (
      {stage0_2[336], stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[58],stage1_4[127],stage1_3[143],stage1_2[143]}
   );
   gpc606_5 gpc144 (
      {stage0_2[342], stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[59],stage1_4[128],stage1_3[144],stage1_2[144]}
   );
   gpc606_5 gpc145 (
      {stage0_2[348], stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[60],stage1_4[129],stage1_3[145],stage1_2[145]}
   );
   gpc606_5 gpc146 (
      {stage0_2[354], stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358], stage0_2[359]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[61],stage1_4[130],stage1_3[146],stage1_2[146]}
   );
   gpc606_5 gpc147 (
      {stage0_2[360], stage0_2[361], stage0_2[362], stage0_2[363], stage0_2[364], stage0_2[365]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[62],stage1_4[131],stage1_3[147],stage1_2[147]}
   );
   gpc606_5 gpc148 (
      {stage0_2[366], stage0_2[367], stage0_2[368], stage0_2[369], stage0_2[370], stage0_2[371]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[63],stage1_4[132],stage1_3[148],stage1_2[148]}
   );
   gpc606_5 gpc149 (
      {stage0_2[372], stage0_2[373], stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[64],stage1_4[133],stage1_3[149],stage1_2[149]}
   );
   gpc606_5 gpc150 (
      {stage0_2[378], stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[65],stage1_4[134],stage1_3[150],stage1_2[150]}
   );
   gpc606_5 gpc151 (
      {stage0_2[384], stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388], stage0_2[389]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[66],stage1_4[135],stage1_3[151],stage1_2[151]}
   );
   gpc615_5 gpc152 (
      {stage0_2[390], stage0_2[391], stage0_2[392], stage0_2[393], stage0_2[394]},
      {stage0_3[334]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[67],stage1_4[136],stage1_3[152],stage1_2[152]}
   );
   gpc615_5 gpc153 (
      {stage0_2[395], stage0_2[396], stage0_2[397], stage0_2[398], stage0_2[399]},
      {stage0_3[335]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[68],stage1_4[137],stage1_3[153],stage1_2[153]}
   );
   gpc615_5 gpc154 (
      {stage0_2[400], stage0_2[401], stage0_2[402], stage0_2[403], stage0_2[404]},
      {stage0_3[336]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage1_6[18],stage1_5[69],stage1_4[138],stage1_3[154],stage1_2[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[405], stage0_2[406], stage0_2[407], stage0_2[408], stage0_2[409]},
      {stage0_3[337]},
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage1_6[19],stage1_5[70],stage1_4[139],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[410], stage0_2[411], stage0_2[412], stage0_2[413], stage0_2[414]},
      {stage0_3[338]},
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage1_6[20],stage1_5[71],stage1_4[140],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_3[339], stage0_3[340], stage0_3[341], stage0_3[342], stage0_3[343]},
      {stage0_4[126]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[21],stage1_5[72],stage1_4[141],stage1_3[157]}
   );
   gpc615_5 gpc158 (
      {stage0_3[344], stage0_3[345], stage0_3[346], stage0_3[347], stage0_3[348]},
      {stage0_4[127]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[22],stage1_5[73],stage1_4[142],stage1_3[158]}
   );
   gpc615_5 gpc159 (
      {stage0_3[349], stage0_3[350], stage0_3[351], stage0_3[352], stage0_3[353]},
      {stage0_4[128]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[23],stage1_5[74],stage1_4[143],stage1_3[159]}
   );
   gpc615_5 gpc160 (
      {stage0_3[354], stage0_3[355], stage0_3[356], stage0_3[357], stage0_3[358]},
      {stage0_4[129]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[24],stage1_5[75],stage1_4[144],stage1_3[160]}
   );
   gpc615_5 gpc161 (
      {stage0_3[359], stage0_3[360], stage0_3[361], stage0_3[362], stage0_3[363]},
      {stage0_4[130]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[25],stage1_5[76],stage1_4[145],stage1_3[161]}
   );
   gpc615_5 gpc162 (
      {stage0_3[364], stage0_3[365], stage0_3[366], stage0_3[367], stage0_3[368]},
      {stage0_4[131]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[26],stage1_5[77],stage1_4[146],stage1_3[162]}
   );
   gpc615_5 gpc163 (
      {stage0_3[369], stage0_3[370], stage0_3[371], stage0_3[372], stage0_3[373]},
      {stage0_4[132]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[27],stage1_5[78],stage1_4[147],stage1_3[163]}
   );
   gpc615_5 gpc164 (
      {stage0_3[374], stage0_3[375], stage0_3[376], stage0_3[377], stage0_3[378]},
      {stage0_4[133]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[28],stage1_5[79],stage1_4[148],stage1_3[164]}
   );
   gpc615_5 gpc165 (
      {stage0_3[379], stage0_3[380], stage0_3[381], stage0_3[382], stage0_3[383]},
      {stage0_4[134]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[29],stage1_5[80],stage1_4[149],stage1_3[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[384], stage0_3[385], stage0_3[386], stage0_3[387], stage0_3[388]},
      {stage0_4[135]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[30],stage1_5[81],stage1_4[150],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[389], stage0_3[390], stage0_3[391], stage0_3[392], stage0_3[393]},
      {stage0_4[136]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[31],stage1_5[82],stage1_4[151],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[394], stage0_3[395], stage0_3[396], stage0_3[397], stage0_3[398]},
      {stage0_4[137]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[32],stage1_5[83],stage1_4[152],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[399], stage0_3[400], stage0_3[401], stage0_3[402], stage0_3[403]},
      {stage0_4[138]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[33],stage1_5[84],stage1_4[153],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[404], stage0_3[405], stage0_3[406], stage0_3[407], stage0_3[408]},
      {stage0_4[139]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[34],stage1_5[85],stage1_4[154],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[409], stage0_3[410], stage0_3[411], stage0_3[412], stage0_3[413]},
      {stage0_4[140]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[35],stage1_5[86],stage1_4[155],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[414], stage0_3[415], stage0_3[416], stage0_3[417], stage0_3[418]},
      {stage0_4[141]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[36],stage1_5[87],stage1_4[156],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[419], stage0_3[420], stage0_3[421], stage0_3[422], stage0_3[423]},
      {stage0_4[142]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[37],stage1_5[88],stage1_4[157],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[424], stage0_3[425], stage0_3[426], stage0_3[427], stage0_3[428]},
      {stage0_4[143]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[38],stage1_5[89],stage1_4[158],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[429], stage0_3[430], stage0_3[431], stage0_3[432], stage0_3[433]},
      {stage0_4[144]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[39],stage1_5[90],stage1_4[159],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[434], stage0_3[435], stage0_3[436], stage0_3[437], stage0_3[438]},
      {stage0_4[145]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[40],stage1_5[91],stage1_4[160],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[439], stage0_3[440], stage0_3[441], stage0_3[442], stage0_3[443]},
      {stage0_4[146]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[41],stage1_5[92],stage1_4[161],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[444], stage0_3[445], stage0_3[446], stage0_3[447], stage0_3[448]},
      {stage0_4[147]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[42],stage1_5[93],stage1_4[162],stage1_3[178]}
   );
   gpc615_5 gpc179 (
      {stage0_3[449], stage0_3[450], stage0_3[451], stage0_3[452], stage0_3[453]},
      {stage0_4[148]},
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage1_7[22],stage1_6[43],stage1_5[94],stage1_4[163],stage1_3[179]}
   );
   gpc615_5 gpc180 (
      {stage0_3[454], stage0_3[455], stage0_3[456], stage0_3[457], stage0_3[458]},
      {stage0_4[149]},
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage1_7[23],stage1_6[44],stage1_5[95],stage1_4[164],stage1_3[180]}
   );
   gpc615_5 gpc181 (
      {stage0_3[459], stage0_3[460], stage0_3[461], stage0_3[462], stage0_3[463]},
      {stage0_4[150]},
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage1_7[24],stage1_6[45],stage1_5[96],stage1_4[165],stage1_3[181]}
   );
   gpc615_5 gpc182 (
      {stage0_3[464], stage0_3[465], stage0_3[466], stage0_3[467], stage0_3[468]},
      {stage0_4[151]},
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage1_7[25],stage1_6[46],stage1_5[97],stage1_4[166],stage1_3[182]}
   );
   gpc615_5 gpc183 (
      {stage0_3[469], stage0_3[470], stage0_3[471], stage0_3[472], stage0_3[473]},
      {stage0_4[152]},
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage1_7[26],stage1_6[47],stage1_5[98],stage1_4[167],stage1_3[183]}
   );
   gpc615_5 gpc184 (
      {stage0_3[474], stage0_3[475], stage0_3[476], stage0_3[477], stage0_3[478]},
      {stage0_4[153]},
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage1_7[27],stage1_6[48],stage1_5[99],stage1_4[168],stage1_3[184]}
   );
   gpc615_5 gpc185 (
      {stage0_3[479], stage0_3[480], stage0_3[481], stage0_3[482], stage0_3[483]},
      {stage0_4[154]},
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage1_7[28],stage1_6[49],stage1_5[100],stage1_4[169],stage1_3[185]}
   );
   gpc606_5 gpc186 (
      {stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[29],stage1_6[50],stage1_5[101],stage1_4[170]}
   );
   gpc606_5 gpc187 (
      {stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[30],stage1_6[51],stage1_5[102],stage1_4[171]}
   );
   gpc606_5 gpc188 (
      {stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[31],stage1_6[52],stage1_5[103],stage1_4[172]}
   );
   gpc606_5 gpc189 (
      {stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[32],stage1_6[53],stage1_5[104],stage1_4[173]}
   );
   gpc606_5 gpc190 (
      {stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[33],stage1_6[54],stage1_5[105],stage1_4[174]}
   );
   gpc606_5 gpc191 (
      {stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188], stage0_4[189], stage0_4[190]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[34],stage1_6[55],stage1_5[106],stage1_4[175]}
   );
   gpc606_5 gpc192 (
      {stage0_4[191], stage0_4[192], stage0_4[193], stage0_4[194], stage0_4[195], stage0_4[196]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[35],stage1_6[56],stage1_5[107],stage1_4[176]}
   );
   gpc606_5 gpc193 (
      {stage0_4[197], stage0_4[198], stage0_4[199], stage0_4[200], stage0_4[201], stage0_4[202]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[36],stage1_6[57],stage1_5[108],stage1_4[177]}
   );
   gpc606_5 gpc194 (
      {stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207], stage0_4[208]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[37],stage1_6[58],stage1_5[109],stage1_4[178]}
   );
   gpc606_5 gpc195 (
      {stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213], stage0_4[214]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[38],stage1_6[59],stage1_5[110],stage1_4[179]}
   );
   gpc606_5 gpc196 (
      {stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218], stage0_4[219], stage0_4[220]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[39],stage1_6[60],stage1_5[111],stage1_4[180]}
   );
   gpc606_5 gpc197 (
      {stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224], stage0_4[225], stage0_4[226]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[40],stage1_6[61],stage1_5[112],stage1_4[181]}
   );
   gpc606_5 gpc198 (
      {stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[41],stage1_6[62],stage1_5[113],stage1_4[182]}
   );
   gpc606_5 gpc199 (
      {stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[42],stage1_6[63],stage1_5[114],stage1_4[183]}
   );
   gpc606_5 gpc200 (
      {stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243], stage0_4[244]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[43],stage1_6[64],stage1_5[115],stage1_4[184]}
   );
   gpc606_5 gpc201 (
      {stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248], stage0_4[249], stage0_4[250]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[44],stage1_6[65],stage1_5[116],stage1_4[185]}
   );
   gpc606_5 gpc202 (
      {stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254], stage0_4[255], stage0_4[256]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[45],stage1_6[66],stage1_5[117],stage1_4[186]}
   );
   gpc606_5 gpc203 (
      {stage0_4[257], stage0_4[258], stage0_4[259], stage0_4[260], stage0_4[261], stage0_4[262]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[46],stage1_6[67],stage1_5[118],stage1_4[187]}
   );
   gpc606_5 gpc204 (
      {stage0_4[263], stage0_4[264], stage0_4[265], stage0_4[266], stage0_4[267], stage0_4[268]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[47],stage1_6[68],stage1_5[119],stage1_4[188]}
   );
   gpc606_5 gpc205 (
      {stage0_4[269], stage0_4[270], stage0_4[271], stage0_4[272], stage0_4[273], stage0_4[274]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[48],stage1_6[69],stage1_5[120],stage1_4[189]}
   );
   gpc606_5 gpc206 (
      {stage0_4[275], stage0_4[276], stage0_4[277], stage0_4[278], stage0_4[279], stage0_4[280]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[49],stage1_6[70],stage1_5[121],stage1_4[190]}
   );
   gpc606_5 gpc207 (
      {stage0_4[281], stage0_4[282], stage0_4[283], stage0_4[284], stage0_4[285], stage0_4[286]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[50],stage1_6[71],stage1_5[122],stage1_4[191]}
   );
   gpc606_5 gpc208 (
      {stage0_4[287], stage0_4[288], stage0_4[289], stage0_4[290], stage0_4[291], stage0_4[292]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[51],stage1_6[72],stage1_5[123],stage1_4[192]}
   );
   gpc606_5 gpc209 (
      {stage0_4[293], stage0_4[294], stage0_4[295], stage0_4[296], stage0_4[297], stage0_4[298]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[52],stage1_6[73],stage1_5[124],stage1_4[193]}
   );
   gpc606_5 gpc210 (
      {stage0_4[299], stage0_4[300], stage0_4[301], stage0_4[302], stage0_4[303], stage0_4[304]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[53],stage1_6[74],stage1_5[125],stage1_4[194]}
   );
   gpc606_5 gpc211 (
      {stage0_4[305], stage0_4[306], stage0_4[307], stage0_4[308], stage0_4[309], stage0_4[310]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[54],stage1_6[75],stage1_5[126],stage1_4[195]}
   );
   gpc606_5 gpc212 (
      {stage0_4[311], stage0_4[312], stage0_4[313], stage0_4[314], stage0_4[315], stage0_4[316]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[55],stage1_6[76],stage1_5[127],stage1_4[196]}
   );
   gpc606_5 gpc213 (
      {stage0_4[317], stage0_4[318], stage0_4[319], stage0_4[320], stage0_4[321], stage0_4[322]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[56],stage1_6[77],stage1_5[128],stage1_4[197]}
   );
   gpc606_5 gpc214 (
      {stage0_4[323], stage0_4[324], stage0_4[325], stage0_4[326], stage0_4[327], stage0_4[328]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[57],stage1_6[78],stage1_5[129],stage1_4[198]}
   );
   gpc606_5 gpc215 (
      {stage0_4[329], stage0_4[330], stage0_4[331], stage0_4[332], stage0_4[333], stage0_4[334]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[58],stage1_6[79],stage1_5[130],stage1_4[199]}
   );
   gpc606_5 gpc216 (
      {stage0_4[335], stage0_4[336], stage0_4[337], stage0_4[338], stage0_4[339], stage0_4[340]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[59],stage1_6[80],stage1_5[131],stage1_4[200]}
   );
   gpc606_5 gpc217 (
      {stage0_4[341], stage0_4[342], stage0_4[343], stage0_4[344], stage0_4[345], stage0_4[346]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[60],stage1_6[81],stage1_5[132],stage1_4[201]}
   );
   gpc606_5 gpc218 (
      {stage0_4[347], stage0_4[348], stage0_4[349], stage0_4[350], stage0_4[351], stage0_4[352]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[61],stage1_6[82],stage1_5[133],stage1_4[202]}
   );
   gpc606_5 gpc219 (
      {stage0_4[353], stage0_4[354], stage0_4[355], stage0_4[356], stage0_4[357], stage0_4[358]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[62],stage1_6[83],stage1_5[134],stage1_4[203]}
   );
   gpc606_5 gpc220 (
      {stage0_4[359], stage0_4[360], stage0_4[361], stage0_4[362], stage0_4[363], stage0_4[364]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[63],stage1_6[84],stage1_5[135],stage1_4[204]}
   );
   gpc606_5 gpc221 (
      {stage0_4[365], stage0_4[366], stage0_4[367], stage0_4[368], stage0_4[369], stage0_4[370]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[64],stage1_6[85],stage1_5[136],stage1_4[205]}
   );
   gpc606_5 gpc222 (
      {stage0_4[371], stage0_4[372], stage0_4[373], stage0_4[374], stage0_4[375], stage0_4[376]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[65],stage1_6[86],stage1_5[137],stage1_4[206]}
   );
   gpc606_5 gpc223 (
      {stage0_4[377], stage0_4[378], stage0_4[379], stage0_4[380], stage0_4[381], stage0_4[382]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[66],stage1_6[87],stage1_5[138],stage1_4[207]}
   );
   gpc606_5 gpc224 (
      {stage0_4[383], stage0_4[384], stage0_4[385], stage0_4[386], stage0_4[387], stage0_4[388]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[67],stage1_6[88],stage1_5[139],stage1_4[208]}
   );
   gpc606_5 gpc225 (
      {stage0_4[389], stage0_4[390], stage0_4[391], stage0_4[392], stage0_4[393], stage0_4[394]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[68],stage1_6[89],stage1_5[140],stage1_4[209]}
   );
   gpc606_5 gpc226 (
      {stage0_4[395], stage0_4[396], stage0_4[397], stage0_4[398], stage0_4[399], stage0_4[400]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[69],stage1_6[90],stage1_5[141],stage1_4[210]}
   );
   gpc606_5 gpc227 (
      {stage0_4[401], stage0_4[402], stage0_4[403], stage0_4[404], stage0_4[405], stage0_4[406]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[70],stage1_6[91],stage1_5[142],stage1_4[211]}
   );
   gpc606_5 gpc228 (
      {stage0_4[407], stage0_4[408], stage0_4[409], stage0_4[410], stage0_4[411], stage0_4[412]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[71],stage1_6[92],stage1_5[143],stage1_4[212]}
   );
   gpc606_5 gpc229 (
      {stage0_4[413], stage0_4[414], stage0_4[415], stage0_4[416], stage0_4[417], stage0_4[418]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[72],stage1_6[93],stage1_5[144],stage1_4[213]}
   );
   gpc606_5 gpc230 (
      {stage0_4[419], stage0_4[420], stage0_4[421], stage0_4[422], stage0_4[423], stage0_4[424]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[73],stage1_6[94],stage1_5[145],stage1_4[214]}
   );
   gpc606_5 gpc231 (
      {stage0_4[425], stage0_4[426], stage0_4[427], stage0_4[428], stage0_4[429], stage0_4[430]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[74],stage1_6[95],stage1_5[146],stage1_4[215]}
   );
   gpc606_5 gpc232 (
      {stage0_4[431], stage0_4[432], stage0_4[433], stage0_4[434], stage0_4[435], stage0_4[436]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[75],stage1_6[96],stage1_5[147],stage1_4[216]}
   );
   gpc606_5 gpc233 (
      {stage0_4[437], stage0_4[438], stage0_4[439], stage0_4[440], stage0_4[441], stage0_4[442]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[76],stage1_6[97],stage1_5[148],stage1_4[217]}
   );
   gpc606_5 gpc234 (
      {stage0_4[443], stage0_4[444], stage0_4[445], stage0_4[446], stage0_4[447], stage0_4[448]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[77],stage1_6[98],stage1_5[149],stage1_4[218]}
   );
   gpc606_5 gpc235 (
      {stage0_4[449], stage0_4[450], stage0_4[451], stage0_4[452], stage0_4[453], stage0_4[454]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[78],stage1_6[99],stage1_5[150],stage1_4[219]}
   );
   gpc606_5 gpc236 (
      {stage0_4[455], stage0_4[456], stage0_4[457], stage0_4[458], stage0_4[459], stage0_4[460]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[79],stage1_6[100],stage1_5[151],stage1_4[220]}
   );
   gpc606_5 gpc237 (
      {stage0_4[461], stage0_4[462], stage0_4[463], stage0_4[464], stage0_4[465], stage0_4[466]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[80],stage1_6[101],stage1_5[152],stage1_4[221]}
   );
   gpc606_5 gpc238 (
      {stage0_4[467], stage0_4[468], stage0_4[469], stage0_4[470], stage0_4[471], stage0_4[472]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[81],stage1_6[102],stage1_5[153],stage1_4[222]}
   );
   gpc606_5 gpc239 (
      {stage0_4[473], stage0_4[474], stage0_4[475], stage0_4[476], stage0_4[477], stage0_4[478]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[82],stage1_6[103],stage1_5[154],stage1_4[223]}
   );
   gpc606_5 gpc240 (
      {stage0_4[479], stage0_4[480], stage0_4[481], stage0_4[482], stage0_4[483], stage0_4[484]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[83],stage1_6[104],stage1_5[155],stage1_4[224]}
   );
   gpc606_5 gpc241 (
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[55],stage1_7[84],stage1_6[105],stage1_5[156]}
   );
   gpc606_5 gpc242 (
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[56],stage1_7[85],stage1_6[106],stage1_5[157]}
   );
   gpc606_5 gpc243 (
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[57],stage1_7[86],stage1_6[107],stage1_5[158]}
   );
   gpc606_5 gpc244 (
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[58],stage1_7[87],stage1_6[108],stage1_5[159]}
   );
   gpc606_5 gpc245 (
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[59],stage1_7[88],stage1_6[109],stage1_5[160]}
   );
   gpc606_5 gpc246 (
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[60],stage1_7[89],stage1_6[110],stage1_5[161]}
   );
   gpc606_5 gpc247 (
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[61],stage1_7[90],stage1_6[111],stage1_5[162]}
   );
   gpc606_5 gpc248 (
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[62],stage1_7[91],stage1_6[112],stage1_5[163]}
   );
   gpc606_5 gpc249 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[63],stage1_7[92],stage1_6[113],stage1_5[164]}
   );
   gpc606_5 gpc250 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[64],stage1_7[93],stage1_6[114],stage1_5[165]}
   );
   gpc606_5 gpc251 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[65],stage1_7[94],stage1_6[115],stage1_5[166]}
   );
   gpc606_5 gpc252 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[66],stage1_7[95],stage1_6[116],stage1_5[167]}
   );
   gpc606_5 gpc253 (
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[67],stage1_7[96],stage1_6[117],stage1_5[168]}
   );
   gpc606_5 gpc254 (
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[68],stage1_7[97],stage1_6[118],stage1_5[169]}
   );
   gpc606_5 gpc255 (
      {stage0_5[258], stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[69],stage1_7[98],stage1_6[119],stage1_5[170]}
   );
   gpc606_5 gpc256 (
      {stage0_5[264], stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[70],stage1_7[99],stage1_6[120],stage1_5[171]}
   );
   gpc606_5 gpc257 (
      {stage0_5[270], stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[71],stage1_7[100],stage1_6[121],stage1_5[172]}
   );
   gpc606_5 gpc258 (
      {stage0_5[276], stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[72],stage1_7[101],stage1_6[122],stage1_5[173]}
   );
   gpc606_5 gpc259 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[73],stage1_7[102],stage1_6[123],stage1_5[174]}
   );
   gpc606_5 gpc260 (
      {stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[74],stage1_7[103],stage1_6[124],stage1_5[175]}
   );
   gpc606_5 gpc261 (
      {stage0_5[294], stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[75],stage1_7[104],stage1_6[125],stage1_5[176]}
   );
   gpc606_5 gpc262 (
      {stage0_5[300], stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[76],stage1_7[105],stage1_6[126],stage1_5[177]}
   );
   gpc606_5 gpc263 (
      {stage0_5[306], stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[77],stage1_7[106],stage1_6[127],stage1_5[178]}
   );
   gpc606_5 gpc264 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[78],stage1_7[107],stage1_6[128],stage1_5[179]}
   );
   gpc606_5 gpc265 (
      {stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[79],stage1_7[108],stage1_6[129],stage1_5[180]}
   );
   gpc606_5 gpc266 (
      {stage0_5[324], stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[80],stage1_7[109],stage1_6[130],stage1_5[181]}
   );
   gpc606_5 gpc267 (
      {stage0_5[330], stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[81],stage1_7[110],stage1_6[131],stage1_5[182]}
   );
   gpc606_5 gpc268 (
      {stage0_5[336], stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[82],stage1_7[111],stage1_6[132],stage1_5[183]}
   );
   gpc606_5 gpc269 (
      {stage0_5[342], stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[83],stage1_7[112],stage1_6[133],stage1_5[184]}
   );
   gpc606_5 gpc270 (
      {stage0_5[348], stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[84],stage1_7[113],stage1_6[134],stage1_5[185]}
   );
   gpc606_5 gpc271 (
      {stage0_5[354], stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[85],stage1_7[114],stage1_6[135],stage1_5[186]}
   );
   gpc606_5 gpc272 (
      {stage0_5[360], stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[86],stage1_7[115],stage1_6[136],stage1_5[187]}
   );
   gpc606_5 gpc273 (
      {stage0_5[366], stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[87],stage1_7[116],stage1_6[137],stage1_5[188]}
   );
   gpc606_5 gpc274 (
      {stage0_5[372], stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[88],stage1_7[117],stage1_6[138],stage1_5[189]}
   );
   gpc606_5 gpc275 (
      {stage0_5[378], stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[89],stage1_7[118],stage1_6[139],stage1_5[190]}
   );
   gpc606_5 gpc276 (
      {stage0_5[384], stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[90],stage1_7[119],stage1_6[140],stage1_5[191]}
   );
   gpc606_5 gpc277 (
      {stage0_5[390], stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[91],stage1_7[120],stage1_6[141],stage1_5[192]}
   );
   gpc606_5 gpc278 (
      {stage0_5[396], stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[92],stage1_7[121],stage1_6[142],stage1_5[193]}
   );
   gpc606_5 gpc279 (
      {stage0_5[402], stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[93],stage1_7[122],stage1_6[143],stage1_5[194]}
   );
   gpc606_5 gpc280 (
      {stage0_5[408], stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[94],stage1_7[123],stage1_6[144],stage1_5[195]}
   );
   gpc606_5 gpc281 (
      {stage0_5[414], stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[95],stage1_7[124],stage1_6[145],stage1_5[196]}
   );
   gpc606_5 gpc282 (
      {stage0_5[420], stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[96],stage1_7[125],stage1_6[146],stage1_5[197]}
   );
   gpc606_5 gpc283 (
      {stage0_5[426], stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[97],stage1_7[126],stage1_6[147],stage1_5[198]}
   );
   gpc606_5 gpc284 (
      {stage0_5[432], stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[98],stage1_7[127],stage1_6[148],stage1_5[199]}
   );
   gpc606_5 gpc285 (
      {stage0_5[438], stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[99],stage1_7[128],stage1_6[149],stage1_5[200]}
   );
   gpc606_5 gpc286 (
      {stage0_5[444], stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[100],stage1_7[129],stage1_6[150],stage1_5[201]}
   );
   gpc606_5 gpc287 (
      {stage0_5[450], stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[101],stage1_7[130],stage1_6[151],stage1_5[202]}
   );
   gpc606_5 gpc288 (
      {stage0_5[456], stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[102],stage1_7[131],stage1_6[152],stage1_5[203]}
   );
   gpc606_5 gpc289 (
      {stage0_5[462], stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[103],stage1_7[132],stage1_6[153],stage1_5[204]}
   );
   gpc606_5 gpc290 (
      {stage0_5[468], stage0_5[469], stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[104],stage1_7[133],stage1_6[154],stage1_5[205]}
   );
   gpc615_5 gpc291 (
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334]},
      {stage0_7[300]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[50],stage1_8[105],stage1_7[134],stage1_6[155]}
   );
   gpc615_5 gpc292 (
      {stage0_6[335], stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339]},
      {stage0_7[301]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[51],stage1_8[106],stage1_7[135],stage1_6[156]}
   );
   gpc615_5 gpc293 (
      {stage0_6[340], stage0_6[341], stage0_6[342], stage0_6[343], stage0_6[344]},
      {stage0_7[302]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[52],stage1_8[107],stage1_7[136],stage1_6[157]}
   );
   gpc615_5 gpc294 (
      {stage0_6[345], stage0_6[346], stage0_6[347], stage0_6[348], stage0_6[349]},
      {stage0_7[303]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[53],stage1_8[108],stage1_7[137],stage1_6[158]}
   );
   gpc615_5 gpc295 (
      {stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353], stage0_6[354]},
      {stage0_7[304]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[54],stage1_8[109],stage1_7[138],stage1_6[159]}
   );
   gpc615_5 gpc296 (
      {stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage0_7[305]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[55],stage1_8[110],stage1_7[139],stage1_6[160]}
   );
   gpc615_5 gpc297 (
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364]},
      {stage0_7[306]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[56],stage1_8[111],stage1_7[140],stage1_6[161]}
   );
   gpc615_5 gpc298 (
      {stage0_6[365], stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369]},
      {stage0_7[307]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[57],stage1_8[112],stage1_7[141],stage1_6[162]}
   );
   gpc615_5 gpc299 (
      {stage0_6[370], stage0_6[371], stage0_6[372], stage0_6[373], stage0_6[374]},
      {stage0_7[308]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[58],stage1_8[113],stage1_7[142],stage1_6[163]}
   );
   gpc615_5 gpc300 (
      {stage0_6[375], stage0_6[376], stage0_6[377], stage0_6[378], stage0_6[379]},
      {stage0_7[309]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[59],stage1_8[114],stage1_7[143],stage1_6[164]}
   );
   gpc615_5 gpc301 (
      {stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383], stage0_6[384]},
      {stage0_7[310]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[60],stage1_8[115],stage1_7[144],stage1_6[165]}
   );
   gpc615_5 gpc302 (
      {stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage0_7[311]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[61],stage1_8[116],stage1_7[145],stage1_6[166]}
   );
   gpc615_5 gpc303 (
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394]},
      {stage0_7[312]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[62],stage1_8[117],stage1_7[146],stage1_6[167]}
   );
   gpc615_5 gpc304 (
      {stage0_6[395], stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399]},
      {stage0_7[313]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[63],stage1_8[118],stage1_7[147],stage1_6[168]}
   );
   gpc615_5 gpc305 (
      {stage0_6[400], stage0_6[401], stage0_6[402], stage0_6[403], stage0_6[404]},
      {stage0_7[314]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[64],stage1_8[119],stage1_7[148],stage1_6[169]}
   );
   gpc615_5 gpc306 (
      {stage0_6[405], stage0_6[406], stage0_6[407], stage0_6[408], stage0_6[409]},
      {stage0_7[315]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[65],stage1_8[120],stage1_7[149],stage1_6[170]}
   );
   gpc615_5 gpc307 (
      {stage0_7[316], stage0_7[317], stage0_7[318], stage0_7[319], stage0_7[320]},
      {stage0_8[96]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[16],stage1_9[66],stage1_8[121],stage1_7[150]}
   );
   gpc615_5 gpc308 (
      {stage0_7[321], stage0_7[322], stage0_7[323], stage0_7[324], stage0_7[325]},
      {stage0_8[97]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[17],stage1_9[67],stage1_8[122],stage1_7[151]}
   );
   gpc615_5 gpc309 (
      {stage0_7[326], stage0_7[327], stage0_7[328], stage0_7[329], stage0_7[330]},
      {stage0_8[98]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[18],stage1_9[68],stage1_8[123],stage1_7[152]}
   );
   gpc615_5 gpc310 (
      {stage0_7[331], stage0_7[332], stage0_7[333], stage0_7[334], stage0_7[335]},
      {stage0_8[99]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[19],stage1_9[69],stage1_8[124],stage1_7[153]}
   );
   gpc615_5 gpc311 (
      {stage0_7[336], stage0_7[337], stage0_7[338], stage0_7[339], stage0_7[340]},
      {stage0_8[100]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[20],stage1_9[70],stage1_8[125],stage1_7[154]}
   );
   gpc615_5 gpc312 (
      {stage0_7[341], stage0_7[342], stage0_7[343], stage0_7[344], stage0_7[345]},
      {stage0_8[101]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[21],stage1_9[71],stage1_8[126],stage1_7[155]}
   );
   gpc615_5 gpc313 (
      {stage0_7[346], stage0_7[347], stage0_7[348], stage0_7[349], stage0_7[350]},
      {stage0_8[102]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[22],stage1_9[72],stage1_8[127],stage1_7[156]}
   );
   gpc615_5 gpc314 (
      {stage0_7[351], stage0_7[352], stage0_7[353], stage0_7[354], stage0_7[355]},
      {stage0_8[103]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[23],stage1_9[73],stage1_8[128],stage1_7[157]}
   );
   gpc615_5 gpc315 (
      {stage0_7[356], stage0_7[357], stage0_7[358], stage0_7[359], stage0_7[360]},
      {stage0_8[104]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[24],stage1_9[74],stage1_8[129],stage1_7[158]}
   );
   gpc615_5 gpc316 (
      {stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364], stage0_7[365]},
      {stage0_8[105]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[25],stage1_9[75],stage1_8[130],stage1_7[159]}
   );
   gpc615_5 gpc317 (
      {stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370]},
      {stage0_8[106]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[26],stage1_9[76],stage1_8[131],stage1_7[160]}
   );
   gpc615_5 gpc318 (
      {stage0_7[371], stage0_7[372], stage0_7[373], stage0_7[374], stage0_7[375]},
      {stage0_8[107]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[27],stage1_9[77],stage1_8[132],stage1_7[161]}
   );
   gpc615_5 gpc319 (
      {stage0_7[376], stage0_7[377], stage0_7[378], stage0_7[379], stage0_7[380]},
      {stage0_8[108]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[28],stage1_9[78],stage1_8[133],stage1_7[162]}
   );
   gpc615_5 gpc320 (
      {stage0_7[381], stage0_7[382], stage0_7[383], stage0_7[384], stage0_7[385]},
      {stage0_8[109]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[29],stage1_9[79],stage1_8[134],stage1_7[163]}
   );
   gpc615_5 gpc321 (
      {stage0_7[386], stage0_7[387], stage0_7[388], stage0_7[389], stage0_7[390]},
      {stage0_8[110]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[30],stage1_9[80],stage1_8[135],stage1_7[164]}
   );
   gpc615_5 gpc322 (
      {stage0_7[391], stage0_7[392], stage0_7[393], stage0_7[394], stage0_7[395]},
      {stage0_8[111]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[31],stage1_9[81],stage1_8[136],stage1_7[165]}
   );
   gpc615_5 gpc323 (
      {stage0_7[396], stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400]},
      {stage0_8[112]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[32],stage1_9[82],stage1_8[137],stage1_7[166]}
   );
   gpc615_5 gpc324 (
      {stage0_7[401], stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405]},
      {stage0_8[113]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[33],stage1_9[83],stage1_8[138],stage1_7[167]}
   );
   gpc615_5 gpc325 (
      {stage0_7[406], stage0_7[407], stage0_7[408], stage0_7[409], stage0_7[410]},
      {stage0_8[114]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[34],stage1_9[84],stage1_8[139],stage1_7[168]}
   );
   gpc615_5 gpc326 (
      {stage0_7[411], stage0_7[412], stage0_7[413], stage0_7[414], stage0_7[415]},
      {stage0_8[115]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[35],stage1_9[85],stage1_8[140],stage1_7[169]}
   );
   gpc615_5 gpc327 (
      {stage0_7[416], stage0_7[417], stage0_7[418], stage0_7[419], stage0_7[420]},
      {stage0_8[116]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[36],stage1_9[86],stage1_8[141],stage1_7[170]}
   );
   gpc615_5 gpc328 (
      {stage0_7[421], stage0_7[422], stage0_7[423], stage0_7[424], stage0_7[425]},
      {stage0_8[117]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[37],stage1_9[87],stage1_8[142],stage1_7[171]}
   );
   gpc615_5 gpc329 (
      {stage0_7[426], stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430]},
      {stage0_8[118]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[38],stage1_9[88],stage1_8[143],stage1_7[172]}
   );
   gpc615_5 gpc330 (
      {stage0_7[431], stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435]},
      {stage0_8[119]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[39],stage1_9[89],stage1_8[144],stage1_7[173]}
   );
   gpc606_5 gpc331 (
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[24],stage1_10[40],stage1_9[90],stage1_8[145]}
   );
   gpc606_5 gpc332 (
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[25],stage1_10[41],stage1_9[91],stage1_8[146]}
   );
   gpc606_5 gpc333 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[26],stage1_10[42],stage1_9[92],stage1_8[147]}
   );
   gpc606_5 gpc334 (
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[27],stage1_10[43],stage1_9[93],stage1_8[148]}
   );
   gpc606_5 gpc335 (
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[28],stage1_10[44],stage1_9[94],stage1_8[149]}
   );
   gpc606_5 gpc336 (
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[29],stage1_10[45],stage1_9[95],stage1_8[150]}
   );
   gpc606_5 gpc337 (
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[30],stage1_10[46],stage1_9[96],stage1_8[151]}
   );
   gpc606_5 gpc338 (
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[31],stage1_10[47],stage1_9[97],stage1_8[152]}
   );
   gpc606_5 gpc339 (
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[32],stage1_10[48],stage1_9[98],stage1_8[153]}
   );
   gpc606_5 gpc340 (
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[33],stage1_10[49],stage1_9[99],stage1_8[154]}
   );
   gpc606_5 gpc341 (
      {stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[34],stage1_10[50],stage1_9[100],stage1_8[155]}
   );
   gpc606_5 gpc342 (
      {stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[35],stage1_10[51],stage1_9[101],stage1_8[156]}
   );
   gpc606_5 gpc343 (
      {stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[36],stage1_10[52],stage1_9[102],stage1_8[157]}
   );
   gpc606_5 gpc344 (
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[37],stage1_10[53],stage1_9[103],stage1_8[158]}
   );
   gpc606_5 gpc345 (
      {stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[38],stage1_10[54],stage1_9[104],stage1_8[159]}
   );
   gpc606_5 gpc346 (
      {stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[39],stage1_10[55],stage1_9[105],stage1_8[160]}
   );
   gpc606_5 gpc347 (
      {stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[40],stage1_10[56],stage1_9[106],stage1_8[161]}
   );
   gpc606_5 gpc348 (
      {stage0_8[222], stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[41],stage1_10[57],stage1_9[107],stage1_8[162]}
   );
   gpc606_5 gpc349 (
      {stage0_8[228], stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[42],stage1_10[58],stage1_9[108],stage1_8[163]}
   );
   gpc606_5 gpc350 (
      {stage0_8[234], stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[43],stage1_10[59],stage1_9[109],stage1_8[164]}
   );
   gpc606_5 gpc351 (
      {stage0_8[240], stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[44],stage1_10[60],stage1_9[110],stage1_8[165]}
   );
   gpc606_5 gpc352 (
      {stage0_8[246], stage0_8[247], stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[45],stage1_10[61],stage1_9[111],stage1_8[166]}
   );
   gpc606_5 gpc353 (
      {stage0_8[252], stage0_8[253], stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[46],stage1_10[62],stage1_9[112],stage1_8[167]}
   );
   gpc606_5 gpc354 (
      {stage0_8[258], stage0_8[259], stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[47],stage1_10[63],stage1_9[113],stage1_8[168]}
   );
   gpc606_5 gpc355 (
      {stage0_8[264], stage0_8[265], stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[48],stage1_10[64],stage1_9[114],stage1_8[169]}
   );
   gpc606_5 gpc356 (
      {stage0_8[270], stage0_8[271], stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[49],stage1_10[65],stage1_9[115],stage1_8[170]}
   );
   gpc606_5 gpc357 (
      {stage0_8[276], stage0_8[277], stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[50],stage1_10[66],stage1_9[116],stage1_8[171]}
   );
   gpc606_5 gpc358 (
      {stage0_8[282], stage0_8[283], stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[51],stage1_10[67],stage1_9[117],stage1_8[172]}
   );
   gpc606_5 gpc359 (
      {stage0_8[288], stage0_8[289], stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[52],stage1_10[68],stage1_9[118],stage1_8[173]}
   );
   gpc606_5 gpc360 (
      {stage0_8[294], stage0_8[295], stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[53],stage1_10[69],stage1_9[119],stage1_8[174]}
   );
   gpc606_5 gpc361 (
      {stage0_8[300], stage0_8[301], stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[54],stage1_10[70],stage1_9[120],stage1_8[175]}
   );
   gpc606_5 gpc362 (
      {stage0_8[306], stage0_8[307], stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[55],stage1_10[71],stage1_9[121],stage1_8[176]}
   );
   gpc606_5 gpc363 (
      {stage0_8[312], stage0_8[313], stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[56],stage1_10[72],stage1_9[122],stage1_8[177]}
   );
   gpc606_5 gpc364 (
      {stage0_8[318], stage0_8[319], stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[57],stage1_10[73],stage1_9[123],stage1_8[178]}
   );
   gpc606_5 gpc365 (
      {stage0_8[324], stage0_8[325], stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[58],stage1_10[74],stage1_9[124],stage1_8[179]}
   );
   gpc606_5 gpc366 (
      {stage0_8[330], stage0_8[331], stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[59],stage1_10[75],stage1_9[125],stage1_8[180]}
   );
   gpc606_5 gpc367 (
      {stage0_8[336], stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[60],stage1_10[76],stage1_9[126],stage1_8[181]}
   );
   gpc606_5 gpc368 (
      {stage0_8[342], stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[61],stage1_10[77],stage1_9[127],stage1_8[182]}
   );
   gpc606_5 gpc369 (
      {stage0_8[348], stage0_8[349], stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[62],stage1_10[78],stage1_9[128],stage1_8[183]}
   );
   gpc606_5 gpc370 (
      {stage0_8[354], stage0_8[355], stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[63],stage1_10[79],stage1_9[129],stage1_8[184]}
   );
   gpc606_5 gpc371 (
      {stage0_8[360], stage0_8[361], stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[64],stage1_10[80],stage1_9[130],stage1_8[185]}
   );
   gpc606_5 gpc372 (
      {stage0_8[366], stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[65],stage1_10[81],stage1_9[131],stage1_8[186]}
   );
   gpc606_5 gpc373 (
      {stage0_8[372], stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[66],stage1_10[82],stage1_9[132],stage1_8[187]}
   );
   gpc606_5 gpc374 (
      {stage0_8[378], stage0_8[379], stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[67],stage1_10[83],stage1_9[133],stage1_8[188]}
   );
   gpc606_5 gpc375 (
      {stage0_8[384], stage0_8[385], stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[68],stage1_10[84],stage1_9[134],stage1_8[189]}
   );
   gpc606_5 gpc376 (
      {stage0_8[390], stage0_8[391], stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[69],stage1_10[85],stage1_9[135],stage1_8[190]}
   );
   gpc606_5 gpc377 (
      {stage0_8[396], stage0_8[397], stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[70],stage1_10[86],stage1_9[136],stage1_8[191]}
   );
   gpc606_5 gpc378 (
      {stage0_8[402], stage0_8[403], stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[71],stage1_10[87],stage1_9[137],stage1_8[192]}
   );
   gpc606_5 gpc379 (
      {stage0_8[408], stage0_8[409], stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[72],stage1_10[88],stage1_9[138],stage1_8[193]}
   );
   gpc606_5 gpc380 (
      {stage0_8[414], stage0_8[415], stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419]},
      {stage0_10[294], stage0_10[295], stage0_10[296], stage0_10[297], stage0_10[298], stage0_10[299]},
      {stage1_12[49],stage1_11[73],stage1_10[89],stage1_9[139],stage1_8[194]}
   );
   gpc606_5 gpc381 (
      {stage0_8[420], stage0_8[421], stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425]},
      {stage0_10[300], stage0_10[301], stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305]},
      {stage1_12[50],stage1_11[74],stage1_10[90],stage1_9[140],stage1_8[195]}
   );
   gpc606_5 gpc382 (
      {stage0_8[426], stage0_8[427], stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431]},
      {stage0_10[306], stage0_10[307], stage0_10[308], stage0_10[309], stage0_10[310], stage0_10[311]},
      {stage1_12[51],stage1_11[75],stage1_10[91],stage1_9[141],stage1_8[196]}
   );
   gpc606_5 gpc383 (
      {stage0_8[432], stage0_8[433], stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437]},
      {stage0_10[312], stage0_10[313], stage0_10[314], stage0_10[315], stage0_10[316], stage0_10[317]},
      {stage1_12[52],stage1_11[76],stage1_10[92],stage1_9[142],stage1_8[197]}
   );
   gpc606_5 gpc384 (
      {stage0_8[438], stage0_8[439], stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443]},
      {stage0_10[318], stage0_10[319], stage0_10[320], stage0_10[321], stage0_10[322], stage0_10[323]},
      {stage1_12[53],stage1_11[77],stage1_10[93],stage1_9[143],stage1_8[198]}
   );
   gpc606_5 gpc385 (
      {stage0_8[444], stage0_8[445], stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449]},
      {stage0_10[324], stage0_10[325], stage0_10[326], stage0_10[327], stage0_10[328], stage0_10[329]},
      {stage1_12[54],stage1_11[78],stage1_10[94],stage1_9[144],stage1_8[199]}
   );
   gpc606_5 gpc386 (
      {stage0_8[450], stage0_8[451], stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455]},
      {stage0_10[330], stage0_10[331], stage0_10[332], stage0_10[333], stage0_10[334], stage0_10[335]},
      {stage1_12[55],stage1_11[79],stage1_10[95],stage1_9[145],stage1_8[200]}
   );
   gpc606_5 gpc387 (
      {stage0_8[456], stage0_8[457], stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461]},
      {stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339], stage0_10[340], stage0_10[341]},
      {stage1_12[56],stage1_11[80],stage1_10[96],stage1_9[146],stage1_8[201]}
   );
   gpc606_5 gpc388 (
      {stage0_8[462], stage0_8[463], stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467]},
      {stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345], stage0_10[346], stage0_10[347]},
      {stage1_12[57],stage1_11[81],stage1_10[97],stage1_9[147],stage1_8[202]}
   );
   gpc606_5 gpc389 (
      {stage0_8[468], stage0_8[469], stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473]},
      {stage0_10[348], stage0_10[349], stage0_10[350], stage0_10[351], stage0_10[352], stage0_10[353]},
      {stage1_12[58],stage1_11[82],stage1_10[98],stage1_9[148],stage1_8[203]}
   );
   gpc606_5 gpc390 (
      {stage0_8[474], stage0_8[475], stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479]},
      {stage0_10[354], stage0_10[355], stage0_10[356], stage0_10[357], stage0_10[358], stage0_10[359]},
      {stage1_12[59],stage1_11[83],stage1_10[99],stage1_9[149],stage1_8[204]}
   );
   gpc606_5 gpc391 (
      {stage0_8[480], stage0_8[481], stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485]},
      {stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363], stage0_10[364], stage0_10[365]},
      {stage1_12[60],stage1_11[84],stage1_10[100],stage1_9[150],stage1_8[205]}
   );
   gpc117_4 gpc392 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150]},
      {stage0_10[366]},
      {stage0_11[0]},
      {stage1_12[61],stage1_11[85],stage1_10[101],stage1_9[151]}
   );
   gpc117_4 gpc393 (
      {stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155], stage0_9[156], stage0_9[157]},
      {stage0_10[367]},
      {stage0_11[1]},
      {stage1_12[62],stage1_11[86],stage1_10[102],stage1_9[152]}
   );
   gpc117_4 gpc394 (
      {stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164]},
      {stage0_10[368]},
      {stage0_11[2]},
      {stage1_12[63],stage1_11[87],stage1_10[103],stage1_9[153]}
   );
   gpc117_4 gpc395 (
      {stage0_9[165], stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171]},
      {stage0_10[369]},
      {stage0_11[3]},
      {stage1_12[64],stage1_11[88],stage1_10[104],stage1_9[154]}
   );
   gpc606_5 gpc396 (
      {stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177]},
      {stage0_11[4], stage0_11[5], stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9]},
      {stage1_13[0],stage1_12[65],stage1_11[89],stage1_10[105],stage1_9[155]}
   );
   gpc606_5 gpc397 (
      {stage0_9[178], stage0_9[179], stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183]},
      {stage0_11[10], stage0_11[11], stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15]},
      {stage1_13[1],stage1_12[66],stage1_11[90],stage1_10[106],stage1_9[156]}
   );
   gpc606_5 gpc398 (
      {stage0_9[184], stage0_9[185], stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189]},
      {stage0_11[16], stage0_11[17], stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21]},
      {stage1_13[2],stage1_12[67],stage1_11[91],stage1_10[107],stage1_9[157]}
   );
   gpc606_5 gpc399 (
      {stage0_9[190], stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195]},
      {stage0_11[22], stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27]},
      {stage1_13[3],stage1_12[68],stage1_11[92],stage1_10[108],stage1_9[158]}
   );
   gpc606_5 gpc400 (
      {stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200], stage0_9[201]},
      {stage0_11[28], stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33]},
      {stage1_13[4],stage1_12[69],stage1_11[93],stage1_10[109],stage1_9[159]}
   );
   gpc606_5 gpc401 (
      {stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205], stage0_9[206], stage0_9[207]},
      {stage0_11[34], stage0_11[35], stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39]},
      {stage1_13[5],stage1_12[70],stage1_11[94],stage1_10[110],stage1_9[160]}
   );
   gpc606_5 gpc402 (
      {stage0_9[208], stage0_9[209], stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213]},
      {stage0_11[40], stage0_11[41], stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45]},
      {stage1_13[6],stage1_12[71],stage1_11[95],stage1_10[111],stage1_9[161]}
   );
   gpc606_5 gpc403 (
      {stage0_9[214], stage0_9[215], stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219]},
      {stage0_11[46], stage0_11[47], stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51]},
      {stage1_13[7],stage1_12[72],stage1_11[96],stage1_10[112],stage1_9[162]}
   );
   gpc606_5 gpc404 (
      {stage0_9[220], stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225]},
      {stage0_11[52], stage0_11[53], stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57]},
      {stage1_13[8],stage1_12[73],stage1_11[97],stage1_10[113],stage1_9[163]}
   );
   gpc606_5 gpc405 (
      {stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230], stage0_9[231]},
      {stage0_11[58], stage0_11[59], stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63]},
      {stage1_13[9],stage1_12[74],stage1_11[98],stage1_10[114],stage1_9[164]}
   );
   gpc606_5 gpc406 (
      {stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235], stage0_9[236], stage0_9[237]},
      {stage0_11[64], stage0_11[65], stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69]},
      {stage1_13[10],stage1_12[75],stage1_11[99],stage1_10[115],stage1_9[165]}
   );
   gpc606_5 gpc407 (
      {stage0_9[238], stage0_9[239], stage0_9[240], stage0_9[241], stage0_9[242], stage0_9[243]},
      {stage0_11[70], stage0_11[71], stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75]},
      {stage1_13[11],stage1_12[76],stage1_11[100],stage1_10[116],stage1_9[166]}
   );
   gpc606_5 gpc408 (
      {stage0_9[244], stage0_9[245], stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249]},
      {stage0_11[76], stage0_11[77], stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81]},
      {stage1_13[12],stage1_12[77],stage1_11[101],stage1_10[117],stage1_9[167]}
   );
   gpc606_5 gpc409 (
      {stage0_9[250], stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255]},
      {stage0_11[82], stage0_11[83], stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87]},
      {stage1_13[13],stage1_12[78],stage1_11[102],stage1_10[118],stage1_9[168]}
   );
   gpc606_5 gpc410 (
      {stage0_9[256], stage0_9[257], stage0_9[258], stage0_9[259], stage0_9[260], stage0_9[261]},
      {stage0_11[88], stage0_11[89], stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93]},
      {stage1_13[14],stage1_12[79],stage1_11[103],stage1_10[119],stage1_9[169]}
   );
   gpc606_5 gpc411 (
      {stage0_9[262], stage0_9[263], stage0_9[264], stage0_9[265], stage0_9[266], stage0_9[267]},
      {stage0_11[94], stage0_11[95], stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99]},
      {stage1_13[15],stage1_12[80],stage1_11[104],stage1_10[120],stage1_9[170]}
   );
   gpc606_5 gpc412 (
      {stage0_9[268], stage0_9[269], stage0_9[270], stage0_9[271], stage0_9[272], stage0_9[273]},
      {stage0_11[100], stage0_11[101], stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105]},
      {stage1_13[16],stage1_12[81],stage1_11[105],stage1_10[121],stage1_9[171]}
   );
   gpc606_5 gpc413 (
      {stage0_9[274], stage0_9[275], stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279]},
      {stage0_11[106], stage0_11[107], stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111]},
      {stage1_13[17],stage1_12[82],stage1_11[106],stage1_10[122],stage1_9[172]}
   );
   gpc606_5 gpc414 (
      {stage0_9[280], stage0_9[281], stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285]},
      {stage0_11[112], stage0_11[113], stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117]},
      {stage1_13[18],stage1_12[83],stage1_11[107],stage1_10[123],stage1_9[173]}
   );
   gpc606_5 gpc415 (
      {stage0_9[286], stage0_9[287], stage0_9[288], stage0_9[289], stage0_9[290], stage0_9[291]},
      {stage0_11[118], stage0_11[119], stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123]},
      {stage1_13[19],stage1_12[84],stage1_11[108],stage1_10[124],stage1_9[174]}
   );
   gpc606_5 gpc416 (
      {stage0_9[292], stage0_9[293], stage0_9[294], stage0_9[295], stage0_9[296], stage0_9[297]},
      {stage0_11[124], stage0_11[125], stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129]},
      {stage1_13[20],stage1_12[85],stage1_11[109],stage1_10[125],stage1_9[175]}
   );
   gpc606_5 gpc417 (
      {stage0_9[298], stage0_9[299], stage0_9[300], stage0_9[301], stage0_9[302], stage0_9[303]},
      {stage0_11[130], stage0_11[131], stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135]},
      {stage1_13[21],stage1_12[86],stage1_11[110],stage1_10[126],stage1_9[176]}
   );
   gpc606_5 gpc418 (
      {stage0_9[304], stage0_9[305], stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309]},
      {stage0_11[136], stage0_11[137], stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141]},
      {stage1_13[22],stage1_12[87],stage1_11[111],stage1_10[127],stage1_9[177]}
   );
   gpc606_5 gpc419 (
      {stage0_9[310], stage0_9[311], stage0_9[312], stage0_9[313], stage0_9[314], stage0_9[315]},
      {stage0_11[142], stage0_11[143], stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147]},
      {stage1_13[23],stage1_12[88],stage1_11[112],stage1_10[128],stage1_9[178]}
   );
   gpc606_5 gpc420 (
      {stage0_9[316], stage0_9[317], stage0_9[318], stage0_9[319], stage0_9[320], stage0_9[321]},
      {stage0_11[148], stage0_11[149], stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153]},
      {stage1_13[24],stage1_12[89],stage1_11[113],stage1_10[129],stage1_9[179]}
   );
   gpc606_5 gpc421 (
      {stage0_9[322], stage0_9[323], stage0_9[324], stage0_9[325], stage0_9[326], stage0_9[327]},
      {stage0_11[154], stage0_11[155], stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159]},
      {stage1_13[25],stage1_12[90],stage1_11[114],stage1_10[130],stage1_9[180]}
   );
   gpc606_5 gpc422 (
      {stage0_9[328], stage0_9[329], stage0_9[330], stage0_9[331], stage0_9[332], stage0_9[333]},
      {stage0_11[160], stage0_11[161], stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165]},
      {stage1_13[26],stage1_12[91],stage1_11[115],stage1_10[131],stage1_9[181]}
   );
   gpc606_5 gpc423 (
      {stage0_9[334], stage0_9[335], stage0_9[336], stage0_9[337], stage0_9[338], stage0_9[339]},
      {stage0_11[166], stage0_11[167], stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171]},
      {stage1_13[27],stage1_12[92],stage1_11[116],stage1_10[132],stage1_9[182]}
   );
   gpc606_5 gpc424 (
      {stage0_9[340], stage0_9[341], stage0_9[342], stage0_9[343], stage0_9[344], stage0_9[345]},
      {stage0_11[172], stage0_11[173], stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177]},
      {stage1_13[28],stage1_12[93],stage1_11[117],stage1_10[133],stage1_9[183]}
   );
   gpc606_5 gpc425 (
      {stage0_9[346], stage0_9[347], stage0_9[348], stage0_9[349], stage0_9[350], stage0_9[351]},
      {stage0_11[178], stage0_11[179], stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183]},
      {stage1_13[29],stage1_12[94],stage1_11[118],stage1_10[134],stage1_9[184]}
   );
   gpc606_5 gpc426 (
      {stage0_9[352], stage0_9[353], stage0_9[354], stage0_9[355], stage0_9[356], stage0_9[357]},
      {stage0_11[184], stage0_11[185], stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189]},
      {stage1_13[30],stage1_12[95],stage1_11[119],stage1_10[135],stage1_9[185]}
   );
   gpc606_5 gpc427 (
      {stage0_9[358], stage0_9[359], stage0_9[360], stage0_9[361], stage0_9[362], stage0_9[363]},
      {stage0_11[190], stage0_11[191], stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195]},
      {stage1_13[31],stage1_12[96],stage1_11[120],stage1_10[136],stage1_9[186]}
   );
   gpc606_5 gpc428 (
      {stage0_9[364], stage0_9[365], stage0_9[366], stage0_9[367], stage0_9[368], stage0_9[369]},
      {stage0_11[196], stage0_11[197], stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201]},
      {stage1_13[32],stage1_12[97],stage1_11[121],stage1_10[137],stage1_9[187]}
   );
   gpc606_5 gpc429 (
      {stage0_9[370], stage0_9[371], stage0_9[372], stage0_9[373], stage0_9[374], stage0_9[375]},
      {stage0_11[202], stage0_11[203], stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207]},
      {stage1_13[33],stage1_12[98],stage1_11[122],stage1_10[138],stage1_9[188]}
   );
   gpc606_5 gpc430 (
      {stage0_9[376], stage0_9[377], stage0_9[378], stage0_9[379], stage0_9[380], stage0_9[381]},
      {stage0_11[208], stage0_11[209], stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213]},
      {stage1_13[34],stage1_12[99],stage1_11[123],stage1_10[139],stage1_9[189]}
   );
   gpc606_5 gpc431 (
      {stage0_9[382], stage0_9[383], stage0_9[384], stage0_9[385], stage0_9[386], stage0_9[387]},
      {stage0_11[214], stage0_11[215], stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219]},
      {stage1_13[35],stage1_12[100],stage1_11[124],stage1_10[140],stage1_9[190]}
   );
   gpc606_5 gpc432 (
      {stage0_9[388], stage0_9[389], stage0_9[390], stage0_9[391], stage0_9[392], stage0_9[393]},
      {stage0_11[220], stage0_11[221], stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225]},
      {stage1_13[36],stage1_12[101],stage1_11[125],stage1_10[141],stage1_9[191]}
   );
   gpc606_5 gpc433 (
      {stage0_9[394], stage0_9[395], stage0_9[396], stage0_9[397], stage0_9[398], stage0_9[399]},
      {stage0_11[226], stage0_11[227], stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231]},
      {stage1_13[37],stage1_12[102],stage1_11[126],stage1_10[142],stage1_9[192]}
   );
   gpc606_5 gpc434 (
      {stage0_9[400], stage0_9[401], stage0_9[402], stage0_9[403], stage0_9[404], stage0_9[405]},
      {stage0_11[232], stage0_11[233], stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237]},
      {stage1_13[38],stage1_12[103],stage1_11[127],stage1_10[143],stage1_9[193]}
   );
   gpc606_5 gpc435 (
      {stage0_9[406], stage0_9[407], stage0_9[408], stage0_9[409], stage0_9[410], stage0_9[411]},
      {stage0_11[238], stage0_11[239], stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243]},
      {stage1_13[39],stage1_12[104],stage1_11[128],stage1_10[144],stage1_9[194]}
   );
   gpc606_5 gpc436 (
      {stage0_9[412], stage0_9[413], stage0_9[414], stage0_9[415], stage0_9[416], stage0_9[417]},
      {stage0_11[244], stage0_11[245], stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249]},
      {stage1_13[40],stage1_12[105],stage1_11[129],stage1_10[145],stage1_9[195]}
   );
   gpc606_5 gpc437 (
      {stage0_9[418], stage0_9[419], stage0_9[420], stage0_9[421], stage0_9[422], stage0_9[423]},
      {stage0_11[250], stage0_11[251], stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255]},
      {stage1_13[41],stage1_12[106],stage1_11[130],stage1_10[146],stage1_9[196]}
   );
   gpc606_5 gpc438 (
      {stage0_9[424], stage0_9[425], stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429]},
      {stage0_11[256], stage0_11[257], stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261]},
      {stage1_13[42],stage1_12[107],stage1_11[131],stage1_10[147],stage1_9[197]}
   );
   gpc606_5 gpc439 (
      {stage0_9[430], stage0_9[431], stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435]},
      {stage0_11[262], stage0_11[263], stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267]},
      {stage1_13[43],stage1_12[108],stage1_11[132],stage1_10[148],stage1_9[198]}
   );
   gpc606_5 gpc440 (
      {stage0_9[436], stage0_9[437], stage0_9[438], stage0_9[439], stage0_9[440], stage0_9[441]},
      {stage0_11[268], stage0_11[269], stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273]},
      {stage1_13[44],stage1_12[109],stage1_11[133],stage1_10[149],stage1_9[199]}
   );
   gpc606_5 gpc441 (
      {stage0_9[442], stage0_9[443], stage0_9[444], stage0_9[445], stage0_9[446], stage0_9[447]},
      {stage0_11[274], stage0_11[275], stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279]},
      {stage1_13[45],stage1_12[110],stage1_11[134],stage1_10[150],stage1_9[200]}
   );
   gpc606_5 gpc442 (
      {stage0_9[448], stage0_9[449], stage0_9[450], stage0_9[451], stage0_9[452], stage0_9[453]},
      {stage0_11[280], stage0_11[281], stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285]},
      {stage1_13[46],stage1_12[111],stage1_11[135],stage1_10[151],stage1_9[201]}
   );
   gpc606_5 gpc443 (
      {stage0_9[454], stage0_9[455], stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459]},
      {stage0_11[286], stage0_11[287], stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291]},
      {stage1_13[47],stage1_12[112],stage1_11[136],stage1_10[152],stage1_9[202]}
   );
   gpc606_5 gpc444 (
      {stage0_9[460], stage0_9[461], stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465]},
      {stage0_11[292], stage0_11[293], stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297]},
      {stage1_13[48],stage1_12[113],stage1_11[137],stage1_10[153],stage1_9[203]}
   );
   gpc606_5 gpc445 (
      {stage0_9[466], stage0_9[467], stage0_9[468], stage0_9[469], stage0_9[470], stage0_9[471]},
      {stage0_11[298], stage0_11[299], stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303]},
      {stage1_13[49],stage1_12[114],stage1_11[138],stage1_10[154],stage1_9[204]}
   );
   gpc606_5 gpc446 (
      {stage0_9[472], stage0_9[473], stage0_9[474], stage0_9[475], stage0_9[476], stage0_9[477]},
      {stage0_11[304], stage0_11[305], stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309]},
      {stage1_13[50],stage1_12[115],stage1_11[139],stage1_10[155],stage1_9[205]}
   );
   gpc615_5 gpc447 (
      {stage0_10[370], stage0_10[371], stage0_10[372], stage0_10[373], stage0_10[374]},
      {stage0_11[310]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[51],stage1_12[116],stage1_11[140],stage1_10[156]}
   );
   gpc615_5 gpc448 (
      {stage0_10[375], stage0_10[376], stage0_10[377], stage0_10[378], stage0_10[379]},
      {stage0_11[311]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[52],stage1_12[117],stage1_11[141],stage1_10[157]}
   );
   gpc615_5 gpc449 (
      {stage0_10[380], stage0_10[381], stage0_10[382], stage0_10[383], stage0_10[384]},
      {stage0_11[312]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[53],stage1_12[118],stage1_11[142],stage1_10[158]}
   );
   gpc615_5 gpc450 (
      {stage0_10[385], stage0_10[386], stage0_10[387], stage0_10[388], stage0_10[389]},
      {stage0_11[313]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[54],stage1_12[119],stage1_11[143],stage1_10[159]}
   );
   gpc615_5 gpc451 (
      {stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393], stage0_10[394]},
      {stage0_11[314]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[55],stage1_12[120],stage1_11[144],stage1_10[160]}
   );
   gpc615_5 gpc452 (
      {stage0_10[395], stage0_10[396], stage0_10[397], stage0_10[398], stage0_10[399]},
      {stage0_11[315]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[56],stage1_12[121],stage1_11[145],stage1_10[161]}
   );
   gpc615_5 gpc453 (
      {stage0_10[400], stage0_10[401], stage0_10[402], stage0_10[403], stage0_10[404]},
      {stage0_11[316]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[57],stage1_12[122],stage1_11[146],stage1_10[162]}
   );
   gpc615_5 gpc454 (
      {stage0_10[405], stage0_10[406], stage0_10[407], stage0_10[408], stage0_10[409]},
      {stage0_11[317]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[58],stage1_12[123],stage1_11[147],stage1_10[163]}
   );
   gpc615_5 gpc455 (
      {stage0_10[410], stage0_10[411], stage0_10[412], stage0_10[413], stage0_10[414]},
      {stage0_11[318]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[59],stage1_12[124],stage1_11[148],stage1_10[164]}
   );
   gpc615_5 gpc456 (
      {stage0_10[415], stage0_10[416], stage0_10[417], stage0_10[418], stage0_10[419]},
      {stage0_11[319]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[60],stage1_12[125],stage1_11[149],stage1_10[165]}
   );
   gpc615_5 gpc457 (
      {stage0_10[420], stage0_10[421], stage0_10[422], stage0_10[423], stage0_10[424]},
      {stage0_11[320]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[61],stage1_12[126],stage1_11[150],stage1_10[166]}
   );
   gpc615_5 gpc458 (
      {stage0_10[425], stage0_10[426], stage0_10[427], stage0_10[428], stage0_10[429]},
      {stage0_11[321]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[62],stage1_12[127],stage1_11[151],stage1_10[167]}
   );
   gpc615_5 gpc459 (
      {stage0_10[430], stage0_10[431], stage0_10[432], stage0_10[433], stage0_10[434]},
      {stage0_11[322]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[63],stage1_12[128],stage1_11[152],stage1_10[168]}
   );
   gpc615_5 gpc460 (
      {stage0_10[435], stage0_10[436], stage0_10[437], stage0_10[438], stage0_10[439]},
      {stage0_11[323]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[64],stage1_12[129],stage1_11[153],stage1_10[169]}
   );
   gpc615_5 gpc461 (
      {stage0_10[440], stage0_10[441], stage0_10[442], stage0_10[443], stage0_10[444]},
      {stage0_11[324]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[65],stage1_12[130],stage1_11[154],stage1_10[170]}
   );
   gpc615_5 gpc462 (
      {stage0_10[445], stage0_10[446], stage0_10[447], stage0_10[448], stage0_10[449]},
      {stage0_11[325]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[66],stage1_12[131],stage1_11[155],stage1_10[171]}
   );
   gpc615_5 gpc463 (
      {stage0_10[450], stage0_10[451], stage0_10[452], stage0_10[453], stage0_10[454]},
      {stage0_11[326]},
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage1_14[16],stage1_13[67],stage1_12[132],stage1_11[156],stage1_10[172]}
   );
   gpc615_5 gpc464 (
      {stage0_10[455], stage0_10[456], stage0_10[457], stage0_10[458], stage0_10[459]},
      {stage0_11[327]},
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage1_14[17],stage1_13[68],stage1_12[133],stage1_11[157],stage1_10[173]}
   );
   gpc615_5 gpc465 (
      {stage0_10[460], stage0_10[461], stage0_10[462], stage0_10[463], stage0_10[464]},
      {stage0_11[328]},
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage1_14[18],stage1_13[69],stage1_12[134],stage1_11[158],stage1_10[174]}
   );
   gpc615_5 gpc466 (
      {stage0_10[465], stage0_10[466], stage0_10[467], stage0_10[468], stage0_10[469]},
      {stage0_11[329]},
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage1_14[19],stage1_13[70],stage1_12[135],stage1_11[159],stage1_10[175]}
   );
   gpc615_5 gpc467 (
      {stage0_10[470], stage0_10[471], stage0_10[472], stage0_10[473], stage0_10[474]},
      {stage0_11[330]},
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage1_14[20],stage1_13[71],stage1_12[136],stage1_11[160],stage1_10[176]}
   );
   gpc615_5 gpc468 (
      {stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage0_12[126]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[21],stage1_13[72],stage1_12[137],stage1_11[161]}
   );
   gpc615_5 gpc469 (
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340]},
      {stage0_12[127]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[22],stage1_13[73],stage1_12[138],stage1_11[162]}
   );
   gpc615_5 gpc470 (
      {stage0_11[341], stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345]},
      {stage0_12[128]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[23],stage1_13[74],stage1_12[139],stage1_11[163]}
   );
   gpc615_5 gpc471 (
      {stage0_11[346], stage0_11[347], stage0_11[348], stage0_11[349], stage0_11[350]},
      {stage0_12[129]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[24],stage1_13[75],stage1_12[140],stage1_11[164]}
   );
   gpc615_5 gpc472 (
      {stage0_11[351], stage0_11[352], stage0_11[353], stage0_11[354], stage0_11[355]},
      {stage0_12[130]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[25],stage1_13[76],stage1_12[141],stage1_11[165]}
   );
   gpc615_5 gpc473 (
      {stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359], stage0_11[360]},
      {stage0_12[131]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[26],stage1_13[77],stage1_12[142],stage1_11[166]}
   );
   gpc615_5 gpc474 (
      {stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage0_12[132]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[27],stage1_13[78],stage1_12[143],stage1_11[167]}
   );
   gpc615_5 gpc475 (
      {stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369], stage0_11[370]},
      {stage0_12[133]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[28],stage1_13[79],stage1_12[144],stage1_11[168]}
   );
   gpc615_5 gpc476 (
      {stage0_11[371], stage0_11[372], stage0_11[373], stage0_11[374], stage0_11[375]},
      {stage0_12[134]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[29],stage1_13[80],stage1_12[145],stage1_11[169]}
   );
   gpc615_5 gpc477 (
      {stage0_11[376], stage0_11[377], stage0_11[378], stage0_11[379], stage0_11[380]},
      {stage0_12[135]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[30],stage1_13[81],stage1_12[146],stage1_11[170]}
   );
   gpc615_5 gpc478 (
      {stage0_11[381], stage0_11[382], stage0_11[383], stage0_11[384], stage0_11[385]},
      {stage0_12[136]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[31],stage1_13[82],stage1_12[147],stage1_11[171]}
   );
   gpc615_5 gpc479 (
      {stage0_11[386], stage0_11[387], stage0_11[388], stage0_11[389], stage0_11[390]},
      {stage0_12[137]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[32],stage1_13[83],stage1_12[148],stage1_11[172]}
   );
   gpc615_5 gpc480 (
      {stage0_11[391], stage0_11[392], stage0_11[393], stage0_11[394], stage0_11[395]},
      {stage0_12[138]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[33],stage1_13[84],stage1_12[149],stage1_11[173]}
   );
   gpc615_5 gpc481 (
      {stage0_11[396], stage0_11[397], stage0_11[398], stage0_11[399], stage0_11[400]},
      {stage0_12[139]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[34],stage1_13[85],stage1_12[150],stage1_11[174]}
   );
   gpc615_5 gpc482 (
      {stage0_11[401], stage0_11[402], stage0_11[403], stage0_11[404], stage0_11[405]},
      {stage0_12[140]},
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage1_15[14],stage1_14[35],stage1_13[86],stage1_12[151],stage1_11[175]}
   );
   gpc615_5 gpc483 (
      {stage0_11[406], stage0_11[407], stage0_11[408], stage0_11[409], stage0_11[410]},
      {stage0_12[141]},
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage1_15[15],stage1_14[36],stage1_13[87],stage1_12[152],stage1_11[176]}
   );
   gpc615_5 gpc484 (
      {stage0_11[411], stage0_11[412], stage0_11[413], stage0_11[414], stage0_11[415]},
      {stage0_12[142]},
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage1_15[16],stage1_14[37],stage1_13[88],stage1_12[153],stage1_11[177]}
   );
   gpc615_5 gpc485 (
      {stage0_11[416], stage0_11[417], stage0_11[418], stage0_11[419], stage0_11[420]},
      {stage0_12[143]},
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage1_15[17],stage1_14[38],stage1_13[89],stage1_12[154],stage1_11[178]}
   );
   gpc615_5 gpc486 (
      {stage0_11[421], stage0_11[422], stage0_11[423], stage0_11[424], stage0_11[425]},
      {stage0_12[144]},
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage1_15[18],stage1_14[39],stage1_13[90],stage1_12[155],stage1_11[179]}
   );
   gpc615_5 gpc487 (
      {stage0_11[426], stage0_11[427], stage0_11[428], stage0_11[429], stage0_11[430]},
      {stage0_12[145]},
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage1_15[19],stage1_14[40],stage1_13[91],stage1_12[156],stage1_11[180]}
   );
   gpc615_5 gpc488 (
      {stage0_11[431], stage0_11[432], stage0_11[433], stage0_11[434], stage0_11[435]},
      {stage0_12[146]},
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage1_15[20],stage1_14[41],stage1_13[92],stage1_12[157],stage1_11[181]}
   );
   gpc615_5 gpc489 (
      {stage0_11[436], stage0_11[437], stage0_11[438], stage0_11[439], stage0_11[440]},
      {stage0_12[147]},
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage1_15[21],stage1_14[42],stage1_13[93],stage1_12[158],stage1_11[182]}
   );
   gpc615_5 gpc490 (
      {stage0_11[441], stage0_11[442], stage0_11[443], stage0_11[444], stage0_11[445]},
      {stage0_12[148]},
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage1_15[22],stage1_14[43],stage1_13[94],stage1_12[159],stage1_11[183]}
   );
   gpc615_5 gpc491 (
      {stage0_11[446], stage0_11[447], stage0_11[448], stage0_11[449], stage0_11[450]},
      {stage0_12[149]},
      {stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage1_15[23],stage1_14[44],stage1_13[95],stage1_12[160],stage1_11[184]}
   );
   gpc606_5 gpc492 (
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[24],stage1_14[45],stage1_13[96],stage1_12[161]}
   );
   gpc606_5 gpc493 (
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[25],stage1_14[46],stage1_13[97],stage1_12[162]}
   );
   gpc606_5 gpc494 (
      {stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165], stage0_12[166], stage0_12[167]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[26],stage1_14[47],stage1_13[98],stage1_12[163]}
   );
   gpc606_5 gpc495 (
      {stage0_12[168], stage0_12[169], stage0_12[170], stage0_12[171], stage0_12[172], stage0_12[173]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[27],stage1_14[48],stage1_13[99],stage1_12[164]}
   );
   gpc606_5 gpc496 (
      {stage0_12[174], stage0_12[175], stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[28],stage1_14[49],stage1_13[100],stage1_12[165]}
   );
   gpc606_5 gpc497 (
      {stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183], stage0_12[184], stage0_12[185]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[29],stage1_14[50],stage1_13[101],stage1_12[166]}
   );
   gpc606_5 gpc498 (
      {stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189], stage0_12[190], stage0_12[191]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[30],stage1_14[51],stage1_13[102],stage1_12[167]}
   );
   gpc606_5 gpc499 (
      {stage0_12[192], stage0_12[193], stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[31],stage1_14[52],stage1_13[103],stage1_12[168]}
   );
   gpc606_5 gpc500 (
      {stage0_12[198], stage0_12[199], stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[32],stage1_14[53],stage1_13[104],stage1_12[169]}
   );
   gpc606_5 gpc501 (
      {stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[33],stage1_14[54],stage1_13[105],stage1_12[170]}
   );
   gpc606_5 gpc502 (
      {stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213], stage0_12[214], stage0_12[215]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[34],stage1_14[55],stage1_13[106],stage1_12[171]}
   );
   gpc606_5 gpc503 (
      {stage0_12[216], stage0_12[217], stage0_12[218], stage0_12[219], stage0_12[220], stage0_12[221]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[35],stage1_14[56],stage1_13[107],stage1_12[172]}
   );
   gpc606_5 gpc504 (
      {stage0_12[222], stage0_12[223], stage0_12[224], stage0_12[225], stage0_12[226], stage0_12[227]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[36],stage1_14[57],stage1_13[108],stage1_12[173]}
   );
   gpc606_5 gpc505 (
      {stage0_12[228], stage0_12[229], stage0_12[230], stage0_12[231], stage0_12[232], stage0_12[233]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[37],stage1_14[58],stage1_13[109],stage1_12[174]}
   );
   gpc606_5 gpc506 (
      {stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237], stage0_12[238], stage0_12[239]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[38],stage1_14[59],stage1_13[110],stage1_12[175]}
   );
   gpc606_5 gpc507 (
      {stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243], stage0_12[244], stage0_12[245]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[39],stage1_14[60],stage1_13[111],stage1_12[176]}
   );
   gpc606_5 gpc508 (
      {stage0_12[246], stage0_12[247], stage0_12[248], stage0_12[249], stage0_12[250], stage0_12[251]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[40],stage1_14[61],stage1_13[112],stage1_12[177]}
   );
   gpc606_5 gpc509 (
      {stage0_12[252], stage0_12[253], stage0_12[254], stage0_12[255], stage0_12[256], stage0_12[257]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[41],stage1_14[62],stage1_13[113],stage1_12[178]}
   );
   gpc606_5 gpc510 (
      {stage0_12[258], stage0_12[259], stage0_12[260], stage0_12[261], stage0_12[262], stage0_12[263]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[42],stage1_14[63],stage1_13[114],stage1_12[179]}
   );
   gpc606_5 gpc511 (
      {stage0_12[264], stage0_12[265], stage0_12[266], stage0_12[267], stage0_12[268], stage0_12[269]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[43],stage1_14[64],stage1_13[115],stage1_12[180]}
   );
   gpc606_5 gpc512 (
      {stage0_12[270], stage0_12[271], stage0_12[272], stage0_12[273], stage0_12[274], stage0_12[275]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[44],stage1_14[65],stage1_13[116],stage1_12[181]}
   );
   gpc606_5 gpc513 (
      {stage0_12[276], stage0_12[277], stage0_12[278], stage0_12[279], stage0_12[280], stage0_12[281]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[45],stage1_14[66],stage1_13[117],stage1_12[182]}
   );
   gpc606_5 gpc514 (
      {stage0_12[282], stage0_12[283], stage0_12[284], stage0_12[285], stage0_12[286], stage0_12[287]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[46],stage1_14[67],stage1_13[118],stage1_12[183]}
   );
   gpc606_5 gpc515 (
      {stage0_12[288], stage0_12[289], stage0_12[290], stage0_12[291], stage0_12[292], stage0_12[293]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[47],stage1_14[68],stage1_13[119],stage1_12[184]}
   );
   gpc606_5 gpc516 (
      {stage0_12[294], stage0_12[295], stage0_12[296], stage0_12[297], stage0_12[298], stage0_12[299]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[48],stage1_14[69],stage1_13[120],stage1_12[185]}
   );
   gpc606_5 gpc517 (
      {stage0_12[300], stage0_12[301], stage0_12[302], stage0_12[303], stage0_12[304], stage0_12[305]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[49],stage1_14[70],stage1_13[121],stage1_12[186]}
   );
   gpc606_5 gpc518 (
      {stage0_12[306], stage0_12[307], stage0_12[308], stage0_12[309], stage0_12[310], stage0_12[311]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[50],stage1_14[71],stage1_13[122],stage1_12[187]}
   );
   gpc606_5 gpc519 (
      {stage0_12[312], stage0_12[313], stage0_12[314], stage0_12[315], stage0_12[316], stage0_12[317]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[51],stage1_14[72],stage1_13[123],stage1_12[188]}
   );
   gpc606_5 gpc520 (
      {stage0_12[318], stage0_12[319], stage0_12[320], stage0_12[321], stage0_12[322], stage0_12[323]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[52],stage1_14[73],stage1_13[124],stage1_12[189]}
   );
   gpc606_5 gpc521 (
      {stage0_12[324], stage0_12[325], stage0_12[326], stage0_12[327], stage0_12[328], stage0_12[329]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[53],stage1_14[74],stage1_13[125],stage1_12[190]}
   );
   gpc606_5 gpc522 (
      {stage0_12[330], stage0_12[331], stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[54],stage1_14[75],stage1_13[126],stage1_12[191]}
   );
   gpc606_5 gpc523 (
      {stage0_12[336], stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340], stage0_12[341]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[55],stage1_14[76],stage1_13[127],stage1_12[192]}
   );
   gpc606_5 gpc524 (
      {stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345], stage0_12[346], stage0_12[347]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[56],stage1_14[77],stage1_13[128],stage1_12[193]}
   );
   gpc606_5 gpc525 (
      {stage0_12[348], stage0_12[349], stage0_12[350], stage0_12[351], stage0_12[352], stage0_12[353]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[57],stage1_14[78],stage1_13[129],stage1_12[194]}
   );
   gpc606_5 gpc526 (
      {stage0_12[354], stage0_12[355], stage0_12[356], stage0_12[357], stage0_12[358], stage0_12[359]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[58],stage1_14[79],stage1_13[130],stage1_12[195]}
   );
   gpc606_5 gpc527 (
      {stage0_12[360], stage0_12[361], stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[59],stage1_14[80],stage1_13[131],stage1_12[196]}
   );
   gpc606_5 gpc528 (
      {stage0_12[366], stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370], stage0_12[371]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[60],stage1_14[81],stage1_13[132],stage1_12[197]}
   );
   gpc606_5 gpc529 (
      {stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375], stage0_12[376], stage0_12[377]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[61],stage1_14[82],stage1_13[133],stage1_12[198]}
   );
   gpc606_5 gpc530 (
      {stage0_12[378], stage0_12[379], stage0_12[380], stage0_12[381], stage0_12[382], stage0_12[383]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[62],stage1_14[83],stage1_13[134],stage1_12[199]}
   );
   gpc606_5 gpc531 (
      {stage0_12[384], stage0_12[385], stage0_12[386], stage0_12[387], stage0_12[388], stage0_12[389]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[63],stage1_14[84],stage1_13[135],stage1_12[200]}
   );
   gpc606_5 gpc532 (
      {stage0_12[390], stage0_12[391], stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[64],stage1_14[85],stage1_13[136],stage1_12[201]}
   );
   gpc606_5 gpc533 (
      {stage0_12[396], stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400], stage0_12[401]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[65],stage1_14[86],stage1_13[137],stage1_12[202]}
   );
   gpc606_5 gpc534 (
      {stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405], stage0_12[406], stage0_12[407]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[66],stage1_14[87],stage1_13[138],stage1_12[203]}
   );
   gpc606_5 gpc535 (
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[43],stage1_15[67],stage1_14[88],stage1_13[139]}
   );
   gpc606_5 gpc536 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[44],stage1_15[68],stage1_14[89],stage1_13[140]}
   );
   gpc606_5 gpc537 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[45],stage1_15[69],stage1_14[90],stage1_13[141]}
   );
   gpc606_5 gpc538 (
      {stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165], stage0_13[166], stage0_13[167]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[46],stage1_15[70],stage1_14[91],stage1_13[142]}
   );
   gpc606_5 gpc539 (
      {stage0_13[168], stage0_13[169], stage0_13[170], stage0_13[171], stage0_13[172], stage0_13[173]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[47],stage1_15[71],stage1_14[92],stage1_13[143]}
   );
   gpc606_5 gpc540 (
      {stage0_13[174], stage0_13[175], stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[48],stage1_15[72],stage1_14[93],stage1_13[144]}
   );
   gpc606_5 gpc541 (
      {stage0_13[180], stage0_13[181], stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[49],stage1_15[73],stage1_14[94],stage1_13[145]}
   );
   gpc606_5 gpc542 (
      {stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189], stage0_13[190], stage0_13[191]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[50],stage1_15[74],stage1_14[95],stage1_13[146]}
   );
   gpc606_5 gpc543 (
      {stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195], stage0_13[196], stage0_13[197]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[51],stage1_15[75],stage1_14[96],stage1_13[147]}
   );
   gpc606_5 gpc544 (
      {stage0_13[198], stage0_13[199], stage0_13[200], stage0_13[201], stage0_13[202], stage0_13[203]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[52],stage1_15[76],stage1_14[97],stage1_13[148]}
   );
   gpc606_5 gpc545 (
      {stage0_13[204], stage0_13[205], stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[53],stage1_15[77],stage1_14[98],stage1_13[149]}
   );
   gpc606_5 gpc546 (
      {stage0_13[210], stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[54],stage1_15[78],stage1_14[99],stage1_13[150]}
   );
   gpc606_5 gpc547 (
      {stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220], stage0_13[221]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[55],stage1_15[79],stage1_14[100],stage1_13[151]}
   );
   gpc606_5 gpc548 (
      {stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225], stage0_13[226], stage0_13[227]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[56],stage1_15[80],stage1_14[101],stage1_13[152]}
   );
   gpc606_5 gpc549 (
      {stage0_13[228], stage0_13[229], stage0_13[230], stage0_13[231], stage0_13[232], stage0_13[233]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[57],stage1_15[81],stage1_14[102],stage1_13[153]}
   );
   gpc606_5 gpc550 (
      {stage0_13[234], stage0_13[235], stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[58],stage1_15[82],stage1_14[103],stage1_13[154]}
   );
   gpc606_5 gpc551 (
      {stage0_13[240], stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[59],stage1_15[83],stage1_14[104],stage1_13[155]}
   );
   gpc606_5 gpc552 (
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250], stage0_13[251]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[60],stage1_15[84],stage1_14[105],stage1_13[156]}
   );
   gpc606_5 gpc553 (
      {stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255], stage0_13[256], stage0_13[257]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[61],stage1_15[85],stage1_14[106],stage1_13[157]}
   );
   gpc606_5 gpc554 (
      {stage0_13[258], stage0_13[259], stage0_13[260], stage0_13[261], stage0_13[262], stage0_13[263]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[62],stage1_15[86],stage1_14[107],stage1_13[158]}
   );
   gpc606_5 gpc555 (
      {stage0_13[264], stage0_13[265], stage0_13[266], stage0_13[267], stage0_13[268], stage0_13[269]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[63],stage1_15[87],stage1_14[108],stage1_13[159]}
   );
   gpc606_5 gpc556 (
      {stage0_13[270], stage0_13[271], stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[64],stage1_15[88],stage1_14[109],stage1_13[160]}
   );
   gpc606_5 gpc557 (
      {stage0_13[276], stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280], stage0_13[281]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[65],stage1_15[89],stage1_14[110],stage1_13[161]}
   );
   gpc606_5 gpc558 (
      {stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285], stage0_13[286], stage0_13[287]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[66],stage1_15[90],stage1_14[111],stage1_13[162]}
   );
   gpc606_5 gpc559 (
      {stage0_13[288], stage0_13[289], stage0_13[290], stage0_13[291], stage0_13[292], stage0_13[293]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[67],stage1_15[91],stage1_14[112],stage1_13[163]}
   );
   gpc606_5 gpc560 (
      {stage0_13[294], stage0_13[295], stage0_13[296], stage0_13[297], stage0_13[298], stage0_13[299]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[68],stage1_15[92],stage1_14[113],stage1_13[164]}
   );
   gpc606_5 gpc561 (
      {stage0_13[300], stage0_13[301], stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[69],stage1_15[93],stage1_14[114],stage1_13[165]}
   );
   gpc606_5 gpc562 (
      {stage0_13[306], stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310], stage0_13[311]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[70],stage1_15[94],stage1_14[115],stage1_13[166]}
   );
   gpc606_5 gpc563 (
      {stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315], stage0_13[316], stage0_13[317]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[71],stage1_15[95],stage1_14[116],stage1_13[167]}
   );
   gpc606_5 gpc564 (
      {stage0_13[318], stage0_13[319], stage0_13[320], stage0_13[321], stage0_13[322], stage0_13[323]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[72],stage1_15[96],stage1_14[117],stage1_13[168]}
   );
   gpc606_5 gpc565 (
      {stage0_13[324], stage0_13[325], stage0_13[326], stage0_13[327], stage0_13[328], stage0_13[329]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[73],stage1_15[97],stage1_14[118],stage1_13[169]}
   );
   gpc606_5 gpc566 (
      {stage0_13[330], stage0_13[331], stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[74],stage1_15[98],stage1_14[119],stage1_13[170]}
   );
   gpc606_5 gpc567 (
      {stage0_13[336], stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340], stage0_13[341]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[75],stage1_15[99],stage1_14[120],stage1_13[171]}
   );
   gpc606_5 gpc568 (
      {stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345], stage0_13[346], stage0_13[347]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[76],stage1_15[100],stage1_14[121],stage1_13[172]}
   );
   gpc606_5 gpc569 (
      {stage0_13[348], stage0_13[349], stage0_13[350], stage0_13[351], stage0_13[352], stage0_13[353]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[77],stage1_15[101],stage1_14[122],stage1_13[173]}
   );
   gpc606_5 gpc570 (
      {stage0_13[354], stage0_13[355], stage0_13[356], stage0_13[357], stage0_13[358], stage0_13[359]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[78],stage1_15[102],stage1_14[123],stage1_13[174]}
   );
   gpc606_5 gpc571 (
      {stage0_13[360], stage0_13[361], stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[79],stage1_15[103],stage1_14[124],stage1_13[175]}
   );
   gpc606_5 gpc572 (
      {stage0_13[366], stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370], stage0_13[371]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[80],stage1_15[104],stage1_14[125],stage1_13[176]}
   );
   gpc606_5 gpc573 (
      {stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375], stage0_13[376], stage0_13[377]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[81],stage1_15[105],stage1_14[126],stage1_13[177]}
   );
   gpc606_5 gpc574 (
      {stage0_13[378], stage0_13[379], stage0_13[380], stage0_13[381], stage0_13[382], stage0_13[383]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[82],stage1_15[106],stage1_14[127],stage1_13[178]}
   );
   gpc606_5 gpc575 (
      {stage0_13[384], stage0_13[385], stage0_13[386], stage0_13[387], stage0_13[388], stage0_13[389]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[83],stage1_15[107],stage1_14[128],stage1_13[179]}
   );
   gpc606_5 gpc576 (
      {stage0_13[390], stage0_13[391], stage0_13[392], stage0_13[393], stage0_13[394], stage0_13[395]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[84],stage1_15[108],stage1_14[129],stage1_13[180]}
   );
   gpc606_5 gpc577 (
      {stage0_13[396], stage0_13[397], stage0_13[398], stage0_13[399], stage0_13[400], stage0_13[401]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[85],stage1_15[109],stage1_14[130],stage1_13[181]}
   );
   gpc606_5 gpc578 (
      {stage0_13[402], stage0_13[403], stage0_13[404], stage0_13[405], stage0_13[406], stage0_13[407]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[86],stage1_15[110],stage1_14[131],stage1_13[182]}
   );
   gpc606_5 gpc579 (
      {stage0_13[408], stage0_13[409], stage0_13[410], stage0_13[411], stage0_13[412], stage0_13[413]},
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268], stage0_15[269]},
      {stage1_17[44],stage1_16[87],stage1_15[111],stage1_14[132],stage1_13[183]}
   );
   gpc606_5 gpc580 (
      {stage0_13[414], stage0_13[415], stage0_13[416], stage0_13[417], stage0_13[418], stage0_13[419]},
      {stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275]},
      {stage1_17[45],stage1_16[88],stage1_15[112],stage1_14[133],stage1_13[184]}
   );
   gpc606_5 gpc581 (
      {stage0_13[420], stage0_13[421], stage0_13[422], stage0_13[423], stage0_13[424], stage0_13[425]},
      {stage0_15[276], stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage1_17[46],stage1_16[89],stage1_15[113],stage1_14[134],stage1_13[185]}
   );
   gpc606_5 gpc582 (
      {stage0_13[426], stage0_13[427], stage0_13[428], stage0_13[429], stage0_13[430], stage0_13[431]},
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287]},
      {stage1_17[47],stage1_16[90],stage1_15[114],stage1_14[135],stage1_13[186]}
   );
   gpc606_5 gpc583 (
      {stage0_13[432], stage0_13[433], stage0_13[434], stage0_13[435], stage0_13[436], stage0_13[437]},
      {stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage1_17[48],stage1_16[91],stage1_15[115],stage1_14[136],stage1_13[187]}
   );
   gpc606_5 gpc584 (
      {stage0_13[438], stage0_13[439], stage0_13[440], stage0_13[441], stage0_13[442], stage0_13[443]},
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298], stage0_15[299]},
      {stage1_17[49],stage1_16[92],stage1_15[116],stage1_14[137],stage1_13[188]}
   );
   gpc606_5 gpc585 (
      {stage0_13[444], stage0_13[445], stage0_13[446], stage0_13[447], stage0_13[448], stage0_13[449]},
      {stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305]},
      {stage1_17[50],stage1_16[93],stage1_15[117],stage1_14[138],stage1_13[189]}
   );
   gpc606_5 gpc586 (
      {stage0_13[450], stage0_13[451], stage0_13[452], stage0_13[453], stage0_13[454], stage0_13[455]},
      {stage0_15[306], stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage1_17[51],stage1_16[94],stage1_15[118],stage1_14[139],stage1_13[190]}
   );
   gpc615_5 gpc587 (
      {stage0_13[456], stage0_13[457], stage0_13[458], stage0_13[459], stage0_13[460]},
      {stage0_14[258]},
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317]},
      {stage1_17[52],stage1_16[95],stage1_15[119],stage1_14[140],stage1_13[191]}
   );
   gpc615_5 gpc588 (
      {stage0_13[461], stage0_13[462], stage0_13[463], stage0_13[464], stage0_13[465]},
      {stage0_14[259]},
      {stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage1_17[53],stage1_16[96],stage1_15[120],stage1_14[141],stage1_13[192]}
   );
   gpc615_5 gpc589 (
      {stage0_13[466], stage0_13[467], stage0_13[468], stage0_13[469], stage0_13[470]},
      {stage0_14[260]},
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328], stage0_15[329]},
      {stage1_17[54],stage1_16[97],stage1_15[121],stage1_14[142],stage1_13[193]}
   );
   gpc615_5 gpc590 (
      {stage0_13[471], stage0_13[472], stage0_13[473], stage0_13[474], stage0_13[475]},
      {stage0_14[261]},
      {stage0_15[330], stage0_15[331], stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335]},
      {stage1_17[55],stage1_16[98],stage1_15[122],stage1_14[143],stage1_13[194]}
   );
   gpc606_5 gpc591 (
      {stage0_14[262], stage0_14[263], stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[56],stage1_16[99],stage1_15[123],stage1_14[144]}
   );
   gpc606_5 gpc592 (
      {stage0_14[268], stage0_14[269], stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[57],stage1_16[100],stage1_15[124],stage1_14[145]}
   );
   gpc606_5 gpc593 (
      {stage0_14[274], stage0_14[275], stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[58],stage1_16[101],stage1_15[125],stage1_14[146]}
   );
   gpc606_5 gpc594 (
      {stage0_14[280], stage0_14[281], stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[59],stage1_16[102],stage1_15[126],stage1_14[147]}
   );
   gpc606_5 gpc595 (
      {stage0_14[286], stage0_14[287], stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[60],stage1_16[103],stage1_15[127],stage1_14[148]}
   );
   gpc606_5 gpc596 (
      {stage0_14[292], stage0_14[293], stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[61],stage1_16[104],stage1_15[128],stage1_14[149]}
   );
   gpc606_5 gpc597 (
      {stage0_14[298], stage0_14[299], stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[62],stage1_16[105],stage1_15[129],stage1_14[150]}
   );
   gpc615_5 gpc598 (
      {stage0_14[304], stage0_14[305], stage0_14[306], stage0_14[307], stage0_14[308]},
      {stage0_15[336]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[63],stage1_16[106],stage1_15[130],stage1_14[151]}
   );
   gpc615_5 gpc599 (
      {stage0_14[309], stage0_14[310], stage0_14[311], stage0_14[312], stage0_14[313]},
      {stage0_15[337]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[64],stage1_16[107],stage1_15[131],stage1_14[152]}
   );
   gpc615_5 gpc600 (
      {stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317], stage0_14[318]},
      {stage0_15[338]},
      {stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59]},
      {stage1_18[9],stage1_17[65],stage1_16[108],stage1_15[132],stage1_14[153]}
   );
   gpc615_5 gpc601 (
      {stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage0_15[339]},
      {stage0_16[60], stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65]},
      {stage1_18[10],stage1_17[66],stage1_16[109],stage1_15[133],stage1_14[154]}
   );
   gpc615_5 gpc602 (
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328]},
      {stage0_15[340]},
      {stage0_16[66], stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71]},
      {stage1_18[11],stage1_17[67],stage1_16[110],stage1_15[134],stage1_14[155]}
   );
   gpc615_5 gpc603 (
      {stage0_14[329], stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333]},
      {stage0_15[341]},
      {stage0_16[72], stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77]},
      {stage1_18[12],stage1_17[68],stage1_16[111],stage1_15[135],stage1_14[156]}
   );
   gpc615_5 gpc604 (
      {stage0_14[334], stage0_14[335], stage0_14[336], stage0_14[337], stage0_14[338]},
      {stage0_15[342]},
      {stage0_16[78], stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83]},
      {stage1_18[13],stage1_17[69],stage1_16[112],stage1_15[136],stage1_14[157]}
   );
   gpc615_5 gpc605 (
      {stage0_14[339], stage0_14[340], stage0_14[341], stage0_14[342], stage0_14[343]},
      {stage0_15[343]},
      {stage0_16[84], stage0_16[85], stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89]},
      {stage1_18[14],stage1_17[70],stage1_16[113],stage1_15[137],stage1_14[158]}
   );
   gpc615_5 gpc606 (
      {stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347], stage0_14[348]},
      {stage0_15[344]},
      {stage0_16[90], stage0_16[91], stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95]},
      {stage1_18[15],stage1_17[71],stage1_16[114],stage1_15[138],stage1_14[159]}
   );
   gpc615_5 gpc607 (
      {stage0_15[345], stage0_15[346], stage0_15[347], stage0_15[348], stage0_15[349]},
      {stage0_16[96]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[16],stage1_17[72],stage1_16[115],stage1_15[139]}
   );
   gpc615_5 gpc608 (
      {stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353], stage0_15[354]},
      {stage0_16[97]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[17],stage1_17[73],stage1_16[116],stage1_15[140]}
   );
   gpc615_5 gpc609 (
      {stage0_15[355], stage0_15[356], stage0_15[357], stage0_15[358], stage0_15[359]},
      {stage0_16[98]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[18],stage1_17[74],stage1_16[117],stage1_15[141]}
   );
   gpc615_5 gpc610 (
      {stage0_15[360], stage0_15[361], stage0_15[362], stage0_15[363], stage0_15[364]},
      {stage0_16[99]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[19],stage1_17[75],stage1_16[118],stage1_15[142]}
   );
   gpc615_5 gpc611 (
      {stage0_15[365], stage0_15[366], stage0_15[367], stage0_15[368], stage0_15[369]},
      {stage0_16[100]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[20],stage1_17[76],stage1_16[119],stage1_15[143]}
   );
   gpc615_5 gpc612 (
      {stage0_15[370], stage0_15[371], stage0_15[372], stage0_15[373], stage0_15[374]},
      {stage0_16[101]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[21],stage1_17[77],stage1_16[120],stage1_15[144]}
   );
   gpc615_5 gpc613 (
      {stage0_15[375], stage0_15[376], stage0_15[377], stage0_15[378], stage0_15[379]},
      {stage0_16[102]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[22],stage1_17[78],stage1_16[121],stage1_15[145]}
   );
   gpc615_5 gpc614 (
      {stage0_15[380], stage0_15[381], stage0_15[382], stage0_15[383], stage0_15[384]},
      {stage0_16[103]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[23],stage1_17[79],stage1_16[122],stage1_15[146]}
   );
   gpc615_5 gpc615 (
      {stage0_15[385], stage0_15[386], stage0_15[387], stage0_15[388], stage0_15[389]},
      {stage0_16[104]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[24],stage1_17[80],stage1_16[123],stage1_15[147]}
   );
   gpc615_5 gpc616 (
      {stage0_15[390], stage0_15[391], stage0_15[392], stage0_15[393], stage0_15[394]},
      {stage0_16[105]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[25],stage1_17[81],stage1_16[124],stage1_15[148]}
   );
   gpc615_5 gpc617 (
      {stage0_15[395], stage0_15[396], stage0_15[397], stage0_15[398], stage0_15[399]},
      {stage0_16[106]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[26],stage1_17[82],stage1_16[125],stage1_15[149]}
   );
   gpc615_5 gpc618 (
      {stage0_15[400], stage0_15[401], stage0_15[402], stage0_15[403], stage0_15[404]},
      {stage0_16[107]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[27],stage1_17[83],stage1_16[126],stage1_15[150]}
   );
   gpc615_5 gpc619 (
      {stage0_15[405], stage0_15[406], stage0_15[407], stage0_15[408], stage0_15[409]},
      {stage0_16[108]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[28],stage1_17[84],stage1_16[127],stage1_15[151]}
   );
   gpc615_5 gpc620 (
      {stage0_15[410], stage0_15[411], stage0_15[412], stage0_15[413], stage0_15[414]},
      {stage0_16[109]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[29],stage1_17[85],stage1_16[128],stage1_15[152]}
   );
   gpc615_5 gpc621 (
      {stage0_15[415], stage0_15[416], stage0_15[417], stage0_15[418], stage0_15[419]},
      {stage0_16[110]},
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage1_19[14],stage1_18[30],stage1_17[86],stage1_16[129],stage1_15[153]}
   );
   gpc615_5 gpc622 (
      {stage0_15[420], stage0_15[421], stage0_15[422], stage0_15[423], stage0_15[424]},
      {stage0_16[111]},
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage1_19[15],stage1_18[31],stage1_17[87],stage1_16[130],stage1_15[154]}
   );
   gpc615_5 gpc623 (
      {stage0_15[425], stage0_15[426], stage0_15[427], stage0_15[428], stage0_15[429]},
      {stage0_16[112]},
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage1_19[16],stage1_18[32],stage1_17[88],stage1_16[131],stage1_15[155]}
   );
   gpc615_5 gpc624 (
      {stage0_15[430], stage0_15[431], stage0_15[432], stage0_15[433], stage0_15[434]},
      {stage0_16[113]},
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage1_19[17],stage1_18[33],stage1_17[89],stage1_16[132],stage1_15[156]}
   );
   gpc615_5 gpc625 (
      {stage0_15[435], stage0_15[436], stage0_15[437], stage0_15[438], stage0_15[439]},
      {stage0_16[114]},
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage1_19[18],stage1_18[34],stage1_17[90],stage1_16[133],stage1_15[157]}
   );
   gpc615_5 gpc626 (
      {stage0_15[440], stage0_15[441], stage0_15[442], stage0_15[443], stage0_15[444]},
      {stage0_16[115]},
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage1_19[19],stage1_18[35],stage1_17[91],stage1_16[134],stage1_15[158]}
   );
   gpc615_5 gpc627 (
      {stage0_15[445], stage0_15[446], stage0_15[447], stage0_15[448], stage0_15[449]},
      {stage0_16[116]},
      {stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124], stage0_17[125]},
      {stage1_19[20],stage1_18[36],stage1_17[92],stage1_16[135],stage1_15[159]}
   );
   gpc615_5 gpc628 (
      {stage0_15[450], stage0_15[451], stage0_15[452], stage0_15[453], stage0_15[454]},
      {stage0_16[117]},
      {stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130], stage0_17[131]},
      {stage1_19[21],stage1_18[37],stage1_17[93],stage1_16[136],stage1_15[160]}
   );
   gpc615_5 gpc629 (
      {stage0_15[455], stage0_15[456], stage0_15[457], stage0_15[458], stage0_15[459]},
      {stage0_16[118]},
      {stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136], stage0_17[137]},
      {stage1_19[22],stage1_18[38],stage1_17[94],stage1_16[137],stage1_15[161]}
   );
   gpc615_5 gpc630 (
      {stage0_15[460], stage0_15[461], stage0_15[462], stage0_15[463], stage0_15[464]},
      {stage0_16[119]},
      {stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142], stage0_17[143]},
      {stage1_19[23],stage1_18[39],stage1_17[95],stage1_16[138],stage1_15[162]}
   );
   gpc615_5 gpc631 (
      {stage0_15[465], stage0_15[466], stage0_15[467], stage0_15[468], stage0_15[469]},
      {stage0_16[120]},
      {stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148], stage0_17[149]},
      {stage1_19[24],stage1_18[40],stage1_17[96],stage1_16[139],stage1_15[163]}
   );
   gpc615_5 gpc632 (
      {stage0_15[470], stage0_15[471], stage0_15[472], stage0_15[473], stage0_15[474]},
      {stage0_16[121]},
      {stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154], stage0_17[155]},
      {stage1_19[25],stage1_18[41],stage1_17[97],stage1_16[140],stage1_15[164]}
   );
   gpc615_5 gpc633 (
      {stage0_15[475], stage0_15[476], stage0_15[477], stage0_15[478], stage0_15[479]},
      {stage0_16[122]},
      {stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160], stage0_17[161]},
      {stage1_19[26],stage1_18[42],stage1_17[98],stage1_16[141],stage1_15[165]}
   );
   gpc606_5 gpc634 (
      {stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126], stage0_16[127], stage0_16[128]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[27],stage1_18[43],stage1_17[99],stage1_16[142]}
   );
   gpc606_5 gpc635 (
      {stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132], stage0_16[133], stage0_16[134]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[28],stage1_18[44],stage1_17[100],stage1_16[143]}
   );
   gpc606_5 gpc636 (
      {stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138], stage0_16[139], stage0_16[140]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[29],stage1_18[45],stage1_17[101],stage1_16[144]}
   );
   gpc606_5 gpc637 (
      {stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144], stage0_16[145], stage0_16[146]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[30],stage1_18[46],stage1_17[102],stage1_16[145]}
   );
   gpc606_5 gpc638 (
      {stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151], stage0_16[152]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[31],stage1_18[47],stage1_17[103],stage1_16[146]}
   );
   gpc606_5 gpc639 (
      {stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157], stage0_16[158]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[32],stage1_18[48],stage1_17[104],stage1_16[147]}
   );
   gpc606_5 gpc640 (
      {stage0_16[159], stage0_16[160], stage0_16[161], stage0_16[162], stage0_16[163], stage0_16[164]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[33],stage1_18[49],stage1_17[105],stage1_16[148]}
   );
   gpc606_5 gpc641 (
      {stage0_16[165], stage0_16[166], stage0_16[167], stage0_16[168], stage0_16[169], stage0_16[170]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[34],stage1_18[50],stage1_17[106],stage1_16[149]}
   );
   gpc606_5 gpc642 (
      {stage0_16[171], stage0_16[172], stage0_16[173], stage0_16[174], stage0_16[175], stage0_16[176]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[35],stage1_18[51],stage1_17[107],stage1_16[150]}
   );
   gpc606_5 gpc643 (
      {stage0_16[177], stage0_16[178], stage0_16[179], stage0_16[180], stage0_16[181], stage0_16[182]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[36],stage1_18[52],stage1_17[108],stage1_16[151]}
   );
   gpc606_5 gpc644 (
      {stage0_16[183], stage0_16[184], stage0_16[185], stage0_16[186], stage0_16[187], stage0_16[188]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[37],stage1_18[53],stage1_17[109],stage1_16[152]}
   );
   gpc606_5 gpc645 (
      {stage0_16[189], stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193], stage0_16[194]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[38],stage1_18[54],stage1_17[110],stage1_16[153]}
   );
   gpc606_5 gpc646 (
      {stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199], stage0_16[200]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[39],stage1_18[55],stage1_17[111],stage1_16[154]}
   );
   gpc606_5 gpc647 (
      {stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204], stage0_16[205], stage0_16[206]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[40],stage1_18[56],stage1_17[112],stage1_16[155]}
   );
   gpc606_5 gpc648 (
      {stage0_16[207], stage0_16[208], stage0_16[209], stage0_16[210], stage0_16[211], stage0_16[212]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[41],stage1_18[57],stage1_17[113],stage1_16[156]}
   );
   gpc606_5 gpc649 (
      {stage0_16[213], stage0_16[214], stage0_16[215], stage0_16[216], stage0_16[217], stage0_16[218]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[42],stage1_18[58],stage1_17[114],stage1_16[157]}
   );
   gpc606_5 gpc650 (
      {stage0_16[219], stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223], stage0_16[224]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[43],stage1_18[59],stage1_17[115],stage1_16[158]}
   );
   gpc606_5 gpc651 (
      {stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229], stage0_16[230]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[44],stage1_18[60],stage1_17[116],stage1_16[159]}
   );
   gpc606_5 gpc652 (
      {stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234], stage0_16[235], stage0_16[236]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[45],stage1_18[61],stage1_17[117],stage1_16[160]}
   );
   gpc606_5 gpc653 (
      {stage0_16[237], stage0_16[238], stage0_16[239], stage0_16[240], stage0_16[241], stage0_16[242]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[46],stage1_18[62],stage1_17[118],stage1_16[161]}
   );
   gpc606_5 gpc654 (
      {stage0_16[243], stage0_16[244], stage0_16[245], stage0_16[246], stage0_16[247], stage0_16[248]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[47],stage1_18[63],stage1_17[119],stage1_16[162]}
   );
   gpc606_5 gpc655 (
      {stage0_16[249], stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253], stage0_16[254]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[48],stage1_18[64],stage1_17[120],stage1_16[163]}
   );
   gpc606_5 gpc656 (
      {stage0_16[255], stage0_16[256], stage0_16[257], stage0_16[258], stage0_16[259], stage0_16[260]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[49],stage1_18[65],stage1_17[121],stage1_16[164]}
   );
   gpc606_5 gpc657 (
      {stage0_16[261], stage0_16[262], stage0_16[263], stage0_16[264], stage0_16[265], stage0_16[266]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[50],stage1_18[66],stage1_17[122],stage1_16[165]}
   );
   gpc606_5 gpc658 (
      {stage0_16[267], stage0_16[268], stage0_16[269], stage0_16[270], stage0_16[271], stage0_16[272]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[51],stage1_18[67],stage1_17[123],stage1_16[166]}
   );
   gpc606_5 gpc659 (
      {stage0_16[273], stage0_16[274], stage0_16[275], stage0_16[276], stage0_16[277], stage0_16[278]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[52],stage1_18[68],stage1_17[124],stage1_16[167]}
   );
   gpc606_5 gpc660 (
      {stage0_16[279], stage0_16[280], stage0_16[281], stage0_16[282], stage0_16[283], stage0_16[284]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[53],stage1_18[69],stage1_17[125],stage1_16[168]}
   );
   gpc606_5 gpc661 (
      {stage0_16[285], stage0_16[286], stage0_16[287], stage0_16[288], stage0_16[289], stage0_16[290]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[54],stage1_18[70],stage1_17[126],stage1_16[169]}
   );
   gpc606_5 gpc662 (
      {stage0_16[291], stage0_16[292], stage0_16[293], stage0_16[294], stage0_16[295], stage0_16[296]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[55],stage1_18[71],stage1_17[127],stage1_16[170]}
   );
   gpc606_5 gpc663 (
      {stage0_16[297], stage0_16[298], stage0_16[299], stage0_16[300], stage0_16[301], stage0_16[302]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[56],stage1_18[72],stage1_17[128],stage1_16[171]}
   );
   gpc606_5 gpc664 (
      {stage0_16[303], stage0_16[304], stage0_16[305], stage0_16[306], stage0_16[307], stage0_16[308]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[57],stage1_18[73],stage1_17[129],stage1_16[172]}
   );
   gpc606_5 gpc665 (
      {stage0_16[309], stage0_16[310], stage0_16[311], stage0_16[312], stage0_16[313], stage0_16[314]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[58],stage1_18[74],stage1_17[130],stage1_16[173]}
   );
   gpc606_5 gpc666 (
      {stage0_16[315], stage0_16[316], stage0_16[317], stage0_16[318], stage0_16[319], stage0_16[320]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[59],stage1_18[75],stage1_17[131],stage1_16[174]}
   );
   gpc606_5 gpc667 (
      {stage0_16[321], stage0_16[322], stage0_16[323], stage0_16[324], stage0_16[325], stage0_16[326]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[60],stage1_18[76],stage1_17[132],stage1_16[175]}
   );
   gpc606_5 gpc668 (
      {stage0_16[327], stage0_16[328], stage0_16[329], stage0_16[330], stage0_16[331], stage0_16[332]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[61],stage1_18[77],stage1_17[133],stage1_16[176]}
   );
   gpc606_5 gpc669 (
      {stage0_16[333], stage0_16[334], stage0_16[335], stage0_16[336], stage0_16[337], stage0_16[338]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[62],stage1_18[78],stage1_17[134],stage1_16[177]}
   );
   gpc606_5 gpc670 (
      {stage0_16[339], stage0_16[340], stage0_16[341], stage0_16[342], stage0_16[343], stage0_16[344]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[63],stage1_18[79],stage1_17[135],stage1_16[178]}
   );
   gpc606_5 gpc671 (
      {stage0_16[345], stage0_16[346], stage0_16[347], stage0_16[348], stage0_16[349], stage0_16[350]},
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226], stage0_18[227]},
      {stage1_20[37],stage1_19[64],stage1_18[80],stage1_17[136],stage1_16[179]}
   );
   gpc606_5 gpc672 (
      {stage0_16[351], stage0_16[352], stage0_16[353], stage0_16[354], stage0_16[355], stage0_16[356]},
      {stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231], stage0_18[232], stage0_18[233]},
      {stage1_20[38],stage1_19[65],stage1_18[81],stage1_17[137],stage1_16[180]}
   );
   gpc606_5 gpc673 (
      {stage0_16[357], stage0_16[358], stage0_16[359], stage0_16[360], stage0_16[361], stage0_16[362]},
      {stage0_18[234], stage0_18[235], stage0_18[236], stage0_18[237], stage0_18[238], stage0_18[239]},
      {stage1_20[39],stage1_19[66],stage1_18[82],stage1_17[138],stage1_16[181]}
   );
   gpc606_5 gpc674 (
      {stage0_16[363], stage0_16[364], stage0_16[365], stage0_16[366], stage0_16[367], stage0_16[368]},
      {stage0_18[240], stage0_18[241], stage0_18[242], stage0_18[243], stage0_18[244], stage0_18[245]},
      {stage1_20[40],stage1_19[67],stage1_18[83],stage1_17[139],stage1_16[182]}
   );
   gpc606_5 gpc675 (
      {stage0_16[369], stage0_16[370], stage0_16[371], stage0_16[372], stage0_16[373], stage0_16[374]},
      {stage0_18[246], stage0_18[247], stage0_18[248], stage0_18[249], stage0_18[250], stage0_18[251]},
      {stage1_20[41],stage1_19[68],stage1_18[84],stage1_17[140],stage1_16[183]}
   );
   gpc606_5 gpc676 (
      {stage0_16[375], stage0_16[376], stage0_16[377], stage0_16[378], stage0_16[379], stage0_16[380]},
      {stage0_18[252], stage0_18[253], stage0_18[254], stage0_18[255], stage0_18[256], stage0_18[257]},
      {stage1_20[42],stage1_19[69],stage1_18[85],stage1_17[141],stage1_16[184]}
   );
   gpc606_5 gpc677 (
      {stage0_16[381], stage0_16[382], stage0_16[383], stage0_16[384], stage0_16[385], stage0_16[386]},
      {stage0_18[258], stage0_18[259], stage0_18[260], stage0_18[261], stage0_18[262], stage0_18[263]},
      {stage1_20[43],stage1_19[70],stage1_18[86],stage1_17[142],stage1_16[185]}
   );
   gpc606_5 gpc678 (
      {stage0_16[387], stage0_16[388], stage0_16[389], stage0_16[390], stage0_16[391], stage0_16[392]},
      {stage0_18[264], stage0_18[265], stage0_18[266], stage0_18[267], stage0_18[268], stage0_18[269]},
      {stage1_20[44],stage1_19[71],stage1_18[87],stage1_17[143],stage1_16[186]}
   );
   gpc606_5 gpc679 (
      {stage0_16[393], stage0_16[394], stage0_16[395], stage0_16[396], stage0_16[397], stage0_16[398]},
      {stage0_18[270], stage0_18[271], stage0_18[272], stage0_18[273], stage0_18[274], stage0_18[275]},
      {stage1_20[45],stage1_19[72],stage1_18[88],stage1_17[144],stage1_16[187]}
   );
   gpc606_5 gpc680 (
      {stage0_16[399], stage0_16[400], stage0_16[401], stage0_16[402], stage0_16[403], stage0_16[404]},
      {stage0_18[276], stage0_18[277], stage0_18[278], stage0_18[279], stage0_18[280], stage0_18[281]},
      {stage1_20[46],stage1_19[73],stage1_18[89],stage1_17[145],stage1_16[188]}
   );
   gpc606_5 gpc681 (
      {stage0_16[405], stage0_16[406], stage0_16[407], stage0_16[408], stage0_16[409], stage0_16[410]},
      {stage0_18[282], stage0_18[283], stage0_18[284], stage0_18[285], stage0_18[286], stage0_18[287]},
      {stage1_20[47],stage1_19[74],stage1_18[90],stage1_17[146],stage1_16[189]}
   );
   gpc606_5 gpc682 (
      {stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166], stage0_17[167]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[48],stage1_19[75],stage1_18[91],stage1_17[147]}
   );
   gpc606_5 gpc683 (
      {stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172], stage0_17[173]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[49],stage1_19[76],stage1_18[92],stage1_17[148]}
   );
   gpc606_5 gpc684 (
      {stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178], stage0_17[179]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[50],stage1_19[77],stage1_18[93],stage1_17[149]}
   );
   gpc606_5 gpc685 (
      {stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184], stage0_17[185]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[51],stage1_19[78],stage1_18[94],stage1_17[150]}
   );
   gpc606_5 gpc686 (
      {stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190], stage0_17[191]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[52],stage1_19[79],stage1_18[95],stage1_17[151]}
   );
   gpc606_5 gpc687 (
      {stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196], stage0_17[197]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[53],stage1_19[80],stage1_18[96],stage1_17[152]}
   );
   gpc606_5 gpc688 (
      {stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202], stage0_17[203]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[54],stage1_19[81],stage1_18[97],stage1_17[153]}
   );
   gpc606_5 gpc689 (
      {stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208], stage0_17[209]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[55],stage1_19[82],stage1_18[98],stage1_17[154]}
   );
   gpc606_5 gpc690 (
      {stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214], stage0_17[215]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[56],stage1_19[83],stage1_18[99],stage1_17[155]}
   );
   gpc606_5 gpc691 (
      {stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220], stage0_17[221]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[57],stage1_19[84],stage1_18[100],stage1_17[156]}
   );
   gpc606_5 gpc692 (
      {stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226], stage0_17[227]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[58],stage1_19[85],stage1_18[101],stage1_17[157]}
   );
   gpc606_5 gpc693 (
      {stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232], stage0_17[233]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[59],stage1_19[86],stage1_18[102],stage1_17[158]}
   );
   gpc606_5 gpc694 (
      {stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238], stage0_17[239]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[60],stage1_19[87],stage1_18[103],stage1_17[159]}
   );
   gpc606_5 gpc695 (
      {stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244], stage0_17[245]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[61],stage1_19[88],stage1_18[104],stage1_17[160]}
   );
   gpc606_5 gpc696 (
      {stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250], stage0_17[251]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[62],stage1_19[89],stage1_18[105],stage1_17[161]}
   );
   gpc606_5 gpc697 (
      {stage0_17[252], stage0_17[253], stage0_17[254], stage0_17[255], stage0_17[256], stage0_17[257]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[63],stage1_19[90],stage1_18[106],stage1_17[162]}
   );
   gpc606_5 gpc698 (
      {stage0_17[258], stage0_17[259], stage0_17[260], stage0_17[261], stage0_17[262], stage0_17[263]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[64],stage1_19[91],stage1_18[107],stage1_17[163]}
   );
   gpc606_5 gpc699 (
      {stage0_17[264], stage0_17[265], stage0_17[266], stage0_17[267], stage0_17[268], stage0_17[269]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[65],stage1_19[92],stage1_18[108],stage1_17[164]}
   );
   gpc606_5 gpc700 (
      {stage0_17[270], stage0_17[271], stage0_17[272], stage0_17[273], stage0_17[274], stage0_17[275]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[66],stage1_19[93],stage1_18[109],stage1_17[165]}
   );
   gpc606_5 gpc701 (
      {stage0_17[276], stage0_17[277], stage0_17[278], stage0_17[279], stage0_17[280], stage0_17[281]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[67],stage1_19[94],stage1_18[110],stage1_17[166]}
   );
   gpc606_5 gpc702 (
      {stage0_17[282], stage0_17[283], stage0_17[284], stage0_17[285], stage0_17[286], stage0_17[287]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[68],stage1_19[95],stage1_18[111],stage1_17[167]}
   );
   gpc606_5 gpc703 (
      {stage0_17[288], stage0_17[289], stage0_17[290], stage0_17[291], stage0_17[292], stage0_17[293]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[69],stage1_19[96],stage1_18[112],stage1_17[168]}
   );
   gpc606_5 gpc704 (
      {stage0_17[294], stage0_17[295], stage0_17[296], stage0_17[297], stage0_17[298], stage0_17[299]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[70],stage1_19[97],stage1_18[113],stage1_17[169]}
   );
   gpc606_5 gpc705 (
      {stage0_17[300], stage0_17[301], stage0_17[302], stage0_17[303], stage0_17[304], stage0_17[305]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[71],stage1_19[98],stage1_18[114],stage1_17[170]}
   );
   gpc606_5 gpc706 (
      {stage0_17[306], stage0_17[307], stage0_17[308], stage0_17[309], stage0_17[310], stage0_17[311]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[72],stage1_19[99],stage1_18[115],stage1_17[171]}
   );
   gpc606_5 gpc707 (
      {stage0_17[312], stage0_17[313], stage0_17[314], stage0_17[315], stage0_17[316], stage0_17[317]},
      {stage0_19[150], stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage1_21[25],stage1_20[73],stage1_19[100],stage1_18[116],stage1_17[172]}
   );
   gpc606_5 gpc708 (
      {stage0_17[318], stage0_17[319], stage0_17[320], stage0_17[321], stage0_17[322], stage0_17[323]},
      {stage0_19[156], stage0_19[157], stage0_19[158], stage0_19[159], stage0_19[160], stage0_19[161]},
      {stage1_21[26],stage1_20[74],stage1_19[101],stage1_18[117],stage1_17[173]}
   );
   gpc606_5 gpc709 (
      {stage0_17[324], stage0_17[325], stage0_17[326], stage0_17[327], stage0_17[328], stage0_17[329]},
      {stage0_19[162], stage0_19[163], stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167]},
      {stage1_21[27],stage1_20[75],stage1_19[102],stage1_18[118],stage1_17[174]}
   );
   gpc606_5 gpc710 (
      {stage0_17[330], stage0_17[331], stage0_17[332], stage0_17[333], stage0_17[334], stage0_17[335]},
      {stage0_19[168], stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage1_21[28],stage1_20[76],stage1_19[103],stage1_18[119],stage1_17[175]}
   );
   gpc606_5 gpc711 (
      {stage0_17[336], stage0_17[337], stage0_17[338], stage0_17[339], stage0_17[340], stage0_17[341]},
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178], stage0_19[179]},
      {stage1_21[29],stage1_20[77],stage1_19[104],stage1_18[120],stage1_17[176]}
   );
   gpc606_5 gpc712 (
      {stage0_17[342], stage0_17[343], stage0_17[344], stage0_17[345], stage0_17[346], stage0_17[347]},
      {stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183], stage0_19[184], stage0_19[185]},
      {stage1_21[30],stage1_20[78],stage1_19[105],stage1_18[121],stage1_17[177]}
   );
   gpc606_5 gpc713 (
      {stage0_17[348], stage0_17[349], stage0_17[350], stage0_17[351], stage0_17[352], stage0_17[353]},
      {stage0_19[186], stage0_19[187], stage0_19[188], stage0_19[189], stage0_19[190], stage0_19[191]},
      {stage1_21[31],stage1_20[79],stage1_19[106],stage1_18[122],stage1_17[178]}
   );
   gpc606_5 gpc714 (
      {stage0_17[354], stage0_17[355], stage0_17[356], stage0_17[357], stage0_17[358], stage0_17[359]},
      {stage0_19[192], stage0_19[193], stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197]},
      {stage1_21[32],stage1_20[80],stage1_19[107],stage1_18[123],stage1_17[179]}
   );
   gpc606_5 gpc715 (
      {stage0_17[360], stage0_17[361], stage0_17[362], stage0_17[363], stage0_17[364], stage0_17[365]},
      {stage0_19[198], stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage1_21[33],stage1_20[81],stage1_19[108],stage1_18[124],stage1_17[180]}
   );
   gpc606_5 gpc716 (
      {stage0_17[366], stage0_17[367], stage0_17[368], stage0_17[369], stage0_17[370], stage0_17[371]},
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208], stage0_19[209]},
      {stage1_21[34],stage1_20[82],stage1_19[109],stage1_18[125],stage1_17[181]}
   );
   gpc606_5 gpc717 (
      {stage0_17[372], stage0_17[373], stage0_17[374], stage0_17[375], stage0_17[376], stage0_17[377]},
      {stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213], stage0_19[214], stage0_19[215]},
      {stage1_21[35],stage1_20[83],stage1_19[110],stage1_18[126],stage1_17[182]}
   );
   gpc606_5 gpc718 (
      {stage0_17[378], stage0_17[379], stage0_17[380], stage0_17[381], stage0_17[382], stage0_17[383]},
      {stage0_19[216], stage0_19[217], stage0_19[218], stage0_19[219], stage0_19[220], stage0_19[221]},
      {stage1_21[36],stage1_20[84],stage1_19[111],stage1_18[127],stage1_17[183]}
   );
   gpc606_5 gpc719 (
      {stage0_17[384], stage0_17[385], stage0_17[386], stage0_17[387], stage0_17[388], stage0_17[389]},
      {stage0_19[222], stage0_19[223], stage0_19[224], stage0_19[225], stage0_19[226], stage0_19[227]},
      {stage1_21[37],stage1_20[85],stage1_19[112],stage1_18[128],stage1_17[184]}
   );
   gpc606_5 gpc720 (
      {stage0_17[390], stage0_17[391], stage0_17[392], stage0_17[393], stage0_17[394], stage0_17[395]},
      {stage0_19[228], stage0_19[229], stage0_19[230], stage0_19[231], stage0_19[232], stage0_19[233]},
      {stage1_21[38],stage1_20[86],stage1_19[113],stage1_18[129],stage1_17[185]}
   );
   gpc606_5 gpc721 (
      {stage0_17[396], stage0_17[397], stage0_17[398], stage0_17[399], stage0_17[400], stage0_17[401]},
      {stage0_19[234], stage0_19[235], stage0_19[236], stage0_19[237], stage0_19[238], stage0_19[239]},
      {stage1_21[39],stage1_20[87],stage1_19[114],stage1_18[130],stage1_17[186]}
   );
   gpc606_5 gpc722 (
      {stage0_18[288], stage0_18[289], stage0_18[290], stage0_18[291], stage0_18[292], stage0_18[293]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[40],stage1_20[88],stage1_19[115],stage1_18[131]}
   );
   gpc606_5 gpc723 (
      {stage0_18[294], stage0_18[295], stage0_18[296], stage0_18[297], stage0_18[298], stage0_18[299]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[41],stage1_20[89],stage1_19[116],stage1_18[132]}
   );
   gpc606_5 gpc724 (
      {stage0_18[300], stage0_18[301], stage0_18[302], stage0_18[303], stage0_18[304], stage0_18[305]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[42],stage1_20[90],stage1_19[117],stage1_18[133]}
   );
   gpc606_5 gpc725 (
      {stage0_18[306], stage0_18[307], stage0_18[308], stage0_18[309], stage0_18[310], stage0_18[311]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[43],stage1_20[91],stage1_19[118],stage1_18[134]}
   );
   gpc615_5 gpc726 (
      {stage0_18[312], stage0_18[313], stage0_18[314], stage0_18[315], stage0_18[316]},
      {stage0_19[240]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[44],stage1_20[92],stage1_19[119],stage1_18[135]}
   );
   gpc615_5 gpc727 (
      {stage0_18[317], stage0_18[318], stage0_18[319], stage0_18[320], stage0_18[321]},
      {stage0_19[241]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[45],stage1_20[93],stage1_19[120],stage1_18[136]}
   );
   gpc615_5 gpc728 (
      {stage0_18[322], stage0_18[323], stage0_18[324], stage0_18[325], stage0_18[326]},
      {stage0_19[242]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[46],stage1_20[94],stage1_19[121],stage1_18[137]}
   );
   gpc615_5 gpc729 (
      {stage0_18[327], stage0_18[328], stage0_18[329], stage0_18[330], stage0_18[331]},
      {stage0_19[243]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[47],stage1_20[95],stage1_19[122],stage1_18[138]}
   );
   gpc615_5 gpc730 (
      {stage0_18[332], stage0_18[333], stage0_18[334], stage0_18[335], stage0_18[336]},
      {stage0_19[244]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[48],stage1_20[96],stage1_19[123],stage1_18[139]}
   );
   gpc615_5 gpc731 (
      {stage0_18[337], stage0_18[338], stage0_18[339], stage0_18[340], stage0_18[341]},
      {stage0_19[245]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[49],stage1_20[97],stage1_19[124],stage1_18[140]}
   );
   gpc615_5 gpc732 (
      {stage0_18[342], stage0_18[343], stage0_18[344], stage0_18[345], stage0_18[346]},
      {stage0_19[246]},
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65]},
      {stage1_22[10],stage1_21[50],stage1_20[98],stage1_19[125],stage1_18[141]}
   );
   gpc615_5 gpc733 (
      {stage0_18[347], stage0_18[348], stage0_18[349], stage0_18[350], stage0_18[351]},
      {stage0_19[247]},
      {stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69], stage0_20[70], stage0_20[71]},
      {stage1_22[11],stage1_21[51],stage1_20[99],stage1_19[126],stage1_18[142]}
   );
   gpc615_5 gpc734 (
      {stage0_18[352], stage0_18[353], stage0_18[354], stage0_18[355], stage0_18[356]},
      {stage0_19[248]},
      {stage0_20[72], stage0_20[73], stage0_20[74], stage0_20[75], stage0_20[76], stage0_20[77]},
      {stage1_22[12],stage1_21[52],stage1_20[100],stage1_19[127],stage1_18[143]}
   );
   gpc615_5 gpc735 (
      {stage0_18[357], stage0_18[358], stage0_18[359], stage0_18[360], stage0_18[361]},
      {stage0_19[249]},
      {stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81], stage0_20[82], stage0_20[83]},
      {stage1_22[13],stage1_21[53],stage1_20[101],stage1_19[128],stage1_18[144]}
   );
   gpc615_5 gpc736 (
      {stage0_18[362], stage0_18[363], stage0_18[364], stage0_18[365], stage0_18[366]},
      {stage0_19[250]},
      {stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88], stage0_20[89]},
      {stage1_22[14],stage1_21[54],stage1_20[102],stage1_19[129],stage1_18[145]}
   );
   gpc615_5 gpc737 (
      {stage0_18[367], stage0_18[368], stage0_18[369], stage0_18[370], stage0_18[371]},
      {stage0_19[251]},
      {stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94], stage0_20[95]},
      {stage1_22[15],stage1_21[55],stage1_20[103],stage1_19[130],stage1_18[146]}
   );
   gpc615_5 gpc738 (
      {stage0_18[372], stage0_18[373], stage0_18[374], stage0_18[375], stage0_18[376]},
      {stage0_19[252]},
      {stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99], stage0_20[100], stage0_20[101]},
      {stage1_22[16],stage1_21[56],stage1_20[104],stage1_19[131],stage1_18[147]}
   );
   gpc615_5 gpc739 (
      {stage0_18[377], stage0_18[378], stage0_18[379], stage0_18[380], stage0_18[381]},
      {stage0_19[253]},
      {stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105], stage0_20[106], stage0_20[107]},
      {stage1_22[17],stage1_21[57],stage1_20[105],stage1_19[132],stage1_18[148]}
   );
   gpc615_5 gpc740 (
      {stage0_18[382], stage0_18[383], stage0_18[384], stage0_18[385], stage0_18[386]},
      {stage0_19[254]},
      {stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111], stage0_20[112], stage0_20[113]},
      {stage1_22[18],stage1_21[58],stage1_20[106],stage1_19[133],stage1_18[149]}
   );
   gpc615_5 gpc741 (
      {stage0_18[387], stage0_18[388], stage0_18[389], stage0_18[390], stage0_18[391]},
      {stage0_19[255]},
      {stage0_20[114], stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118], stage0_20[119]},
      {stage1_22[19],stage1_21[59],stage1_20[107],stage1_19[134],stage1_18[150]}
   );
   gpc615_5 gpc742 (
      {stage0_18[392], stage0_18[393], stage0_18[394], stage0_18[395], stage0_18[396]},
      {stage0_19[256]},
      {stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124], stage0_20[125]},
      {stage1_22[20],stage1_21[60],stage1_20[108],stage1_19[135],stage1_18[151]}
   );
   gpc615_5 gpc743 (
      {stage0_18[397], stage0_18[398], stage0_18[399], stage0_18[400], stage0_18[401]},
      {stage0_19[257]},
      {stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130], stage0_20[131]},
      {stage1_22[21],stage1_21[61],stage1_20[109],stage1_19[136],stage1_18[152]}
   );
   gpc615_5 gpc744 (
      {stage0_18[402], stage0_18[403], stage0_18[404], stage0_18[405], stage0_18[406]},
      {stage0_19[258]},
      {stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136], stage0_20[137]},
      {stage1_22[22],stage1_21[62],stage1_20[110],stage1_19[137],stage1_18[153]}
   );
   gpc615_5 gpc745 (
      {stage0_18[407], stage0_18[408], stage0_18[409], stage0_18[410], stage0_18[411]},
      {stage0_19[259]},
      {stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141], stage0_20[142], stage0_20[143]},
      {stage1_22[23],stage1_21[63],stage1_20[111],stage1_19[138],stage1_18[154]}
   );
   gpc615_5 gpc746 (
      {stage0_18[412], stage0_18[413], stage0_18[414], stage0_18[415], stage0_18[416]},
      {stage0_19[260]},
      {stage0_20[144], stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148], stage0_20[149]},
      {stage1_22[24],stage1_21[64],stage1_20[112],stage1_19[139],stage1_18[155]}
   );
   gpc615_5 gpc747 (
      {stage0_18[417], stage0_18[418], stage0_18[419], stage0_18[420], stage0_18[421]},
      {stage0_19[261]},
      {stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154], stage0_20[155]},
      {stage1_22[25],stage1_21[65],stage1_20[113],stage1_19[140],stage1_18[156]}
   );
   gpc615_5 gpc748 (
      {stage0_18[422], stage0_18[423], stage0_18[424], stage0_18[425], stage0_18[426]},
      {stage0_19[262]},
      {stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160], stage0_20[161]},
      {stage1_22[26],stage1_21[66],stage1_20[114],stage1_19[141],stage1_18[157]}
   );
   gpc615_5 gpc749 (
      {stage0_18[427], stage0_18[428], stage0_18[429], stage0_18[430], stage0_18[431]},
      {stage0_19[263]},
      {stage0_20[162], stage0_20[163], stage0_20[164], stage0_20[165], stage0_20[166], stage0_20[167]},
      {stage1_22[27],stage1_21[67],stage1_20[115],stage1_19[142],stage1_18[158]}
   );
   gpc615_5 gpc750 (
      {stage0_18[432], stage0_18[433], stage0_18[434], stage0_18[435], stage0_18[436]},
      {stage0_19[264]},
      {stage0_20[168], stage0_20[169], stage0_20[170], stage0_20[171], stage0_20[172], stage0_20[173]},
      {stage1_22[28],stage1_21[68],stage1_20[116],stage1_19[143],stage1_18[159]}
   );
   gpc615_5 gpc751 (
      {stage0_18[437], stage0_18[438], stage0_18[439], stage0_18[440], stage0_18[441]},
      {stage0_19[265]},
      {stage0_20[174], stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178], stage0_20[179]},
      {stage1_22[29],stage1_21[69],stage1_20[117],stage1_19[144],stage1_18[160]}
   );
   gpc615_5 gpc752 (
      {stage0_18[442], stage0_18[443], stage0_18[444], stage0_18[445], stage0_18[446]},
      {stage0_19[266]},
      {stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184], stage0_20[185]},
      {stage1_22[30],stage1_21[70],stage1_20[118],stage1_19[145],stage1_18[161]}
   );
   gpc606_5 gpc753 (
      {stage0_19[267], stage0_19[268], stage0_19[269], stage0_19[270], stage0_19[271], stage0_19[272]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[31],stage1_21[71],stage1_20[119],stage1_19[146]}
   );
   gpc606_5 gpc754 (
      {stage0_19[273], stage0_19[274], stage0_19[275], stage0_19[276], stage0_19[277], stage0_19[278]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[32],stage1_21[72],stage1_20[120],stage1_19[147]}
   );
   gpc606_5 gpc755 (
      {stage0_19[279], stage0_19[280], stage0_19[281], stage0_19[282], stage0_19[283], stage0_19[284]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[33],stage1_21[73],stage1_20[121],stage1_19[148]}
   );
   gpc606_5 gpc756 (
      {stage0_19[285], stage0_19[286], stage0_19[287], stage0_19[288], stage0_19[289], stage0_19[290]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[34],stage1_21[74],stage1_20[122],stage1_19[149]}
   );
   gpc606_5 gpc757 (
      {stage0_19[291], stage0_19[292], stage0_19[293], stage0_19[294], stage0_19[295], stage0_19[296]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[35],stage1_21[75],stage1_20[123],stage1_19[150]}
   );
   gpc615_5 gpc758 (
      {stage0_19[297], stage0_19[298], stage0_19[299], stage0_19[300], stage0_19[301]},
      {stage0_20[186]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[36],stage1_21[76],stage1_20[124],stage1_19[151]}
   );
   gpc615_5 gpc759 (
      {stage0_19[302], stage0_19[303], stage0_19[304], stage0_19[305], stage0_19[306]},
      {stage0_20[187]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[37],stage1_21[77],stage1_20[125],stage1_19[152]}
   );
   gpc615_5 gpc760 (
      {stage0_19[307], stage0_19[308], stage0_19[309], stage0_19[310], stage0_19[311]},
      {stage0_20[188]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[38],stage1_21[78],stage1_20[126],stage1_19[153]}
   );
   gpc615_5 gpc761 (
      {stage0_19[312], stage0_19[313], stage0_19[314], stage0_19[315], stage0_19[316]},
      {stage0_20[189]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[39],stage1_21[79],stage1_20[127],stage1_19[154]}
   );
   gpc615_5 gpc762 (
      {stage0_19[317], stage0_19[318], stage0_19[319], stage0_19[320], stage0_19[321]},
      {stage0_20[190]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[40],stage1_21[80],stage1_20[128],stage1_19[155]}
   );
   gpc615_5 gpc763 (
      {stage0_19[322], stage0_19[323], stage0_19[324], stage0_19[325], stage0_19[326]},
      {stage0_20[191]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[41],stage1_21[81],stage1_20[129],stage1_19[156]}
   );
   gpc615_5 gpc764 (
      {stage0_19[327], stage0_19[328], stage0_19[329], stage0_19[330], stage0_19[331]},
      {stage0_20[192]},
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage1_23[11],stage1_22[42],stage1_21[82],stage1_20[130],stage1_19[157]}
   );
   gpc615_5 gpc765 (
      {stage0_19[332], stage0_19[333], stage0_19[334], stage0_19[335], stage0_19[336]},
      {stage0_20[193]},
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage1_23[12],stage1_22[43],stage1_21[83],stage1_20[131],stage1_19[158]}
   );
   gpc615_5 gpc766 (
      {stage0_19[337], stage0_19[338], stage0_19[339], stage0_19[340], stage0_19[341]},
      {stage0_20[194]},
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage1_23[13],stage1_22[44],stage1_21[84],stage1_20[132],stage1_19[159]}
   );
   gpc615_5 gpc767 (
      {stage0_19[342], stage0_19[343], stage0_19[344], stage0_19[345], stage0_19[346]},
      {stage0_20[195]},
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage1_23[14],stage1_22[45],stage1_21[85],stage1_20[133],stage1_19[160]}
   );
   gpc606_5 gpc768 (
      {stage0_20[196], stage0_20[197], stage0_20[198], stage0_20[199], stage0_20[200], stage0_20[201]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[15],stage1_22[46],stage1_21[86],stage1_20[134]}
   );
   gpc606_5 gpc769 (
      {stage0_20[202], stage0_20[203], stage0_20[204], stage0_20[205], stage0_20[206], stage0_20[207]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[16],stage1_22[47],stage1_21[87],stage1_20[135]}
   );
   gpc606_5 gpc770 (
      {stage0_20[208], stage0_20[209], stage0_20[210], stage0_20[211], stage0_20[212], stage0_20[213]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[17],stage1_22[48],stage1_21[88],stage1_20[136]}
   );
   gpc606_5 gpc771 (
      {stage0_20[214], stage0_20[215], stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[18],stage1_22[49],stage1_21[89],stage1_20[137]}
   );
   gpc606_5 gpc772 (
      {stage0_20[220], stage0_20[221], stage0_20[222], stage0_20[223], stage0_20[224], stage0_20[225]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[19],stage1_22[50],stage1_21[90],stage1_20[138]}
   );
   gpc606_5 gpc773 (
      {stage0_20[226], stage0_20[227], stage0_20[228], stage0_20[229], stage0_20[230], stage0_20[231]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[20],stage1_22[51],stage1_21[91],stage1_20[139]}
   );
   gpc606_5 gpc774 (
      {stage0_20[232], stage0_20[233], stage0_20[234], stage0_20[235], stage0_20[236], stage0_20[237]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[21],stage1_22[52],stage1_21[92],stage1_20[140]}
   );
   gpc606_5 gpc775 (
      {stage0_20[238], stage0_20[239], stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[22],stage1_22[53],stage1_21[93],stage1_20[141]}
   );
   gpc606_5 gpc776 (
      {stage0_20[244], stage0_20[245], stage0_20[246], stage0_20[247], stage0_20[248], stage0_20[249]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[23],stage1_22[54],stage1_21[94],stage1_20[142]}
   );
   gpc606_5 gpc777 (
      {stage0_20[250], stage0_20[251], stage0_20[252], stage0_20[253], stage0_20[254], stage0_20[255]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[24],stage1_22[55],stage1_21[95],stage1_20[143]}
   );
   gpc606_5 gpc778 (
      {stage0_20[256], stage0_20[257], stage0_20[258], stage0_20[259], stage0_20[260], stage0_20[261]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[25],stage1_22[56],stage1_21[96],stage1_20[144]}
   );
   gpc606_5 gpc779 (
      {stage0_20[262], stage0_20[263], stage0_20[264], stage0_20[265], stage0_20[266], stage0_20[267]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[26],stage1_22[57],stage1_21[97],stage1_20[145]}
   );
   gpc606_5 gpc780 (
      {stage0_20[268], stage0_20[269], stage0_20[270], stage0_20[271], stage0_20[272], stage0_20[273]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[27],stage1_22[58],stage1_21[98],stage1_20[146]}
   );
   gpc606_5 gpc781 (
      {stage0_20[274], stage0_20[275], stage0_20[276], stage0_20[277], stage0_20[278], stage0_20[279]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[28],stage1_22[59],stage1_21[99],stage1_20[147]}
   );
   gpc606_5 gpc782 (
      {stage0_20[280], stage0_20[281], stage0_20[282], stage0_20[283], stage0_20[284], stage0_20[285]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[29],stage1_22[60],stage1_21[100],stage1_20[148]}
   );
   gpc606_5 gpc783 (
      {stage0_20[286], stage0_20[287], stage0_20[288], stage0_20[289], stage0_20[290], stage0_20[291]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[30],stage1_22[61],stage1_21[101],stage1_20[149]}
   );
   gpc606_5 gpc784 (
      {stage0_20[292], stage0_20[293], stage0_20[294], stage0_20[295], stage0_20[296], stage0_20[297]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[31],stage1_22[62],stage1_21[102],stage1_20[150]}
   );
   gpc606_5 gpc785 (
      {stage0_20[298], stage0_20[299], stage0_20[300], stage0_20[301], stage0_20[302], stage0_20[303]},
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106], stage0_22[107]},
      {stage1_24[17],stage1_23[32],stage1_22[63],stage1_21[103],stage1_20[151]}
   );
   gpc606_5 gpc786 (
      {stage0_20[304], stage0_20[305], stage0_20[306], stage0_20[307], stage0_20[308], stage0_20[309]},
      {stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112], stage0_22[113]},
      {stage1_24[18],stage1_23[33],stage1_22[64],stage1_21[104],stage1_20[152]}
   );
   gpc606_5 gpc787 (
      {stage0_20[310], stage0_20[311], stage0_20[312], stage0_20[313], stage0_20[314], stage0_20[315]},
      {stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118], stage0_22[119]},
      {stage1_24[19],stage1_23[34],stage1_22[65],stage1_21[105],stage1_20[153]}
   );
   gpc606_5 gpc788 (
      {stage0_20[316], stage0_20[317], stage0_20[318], stage0_20[319], stage0_20[320], stage0_20[321]},
      {stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124], stage0_22[125]},
      {stage1_24[20],stage1_23[35],stage1_22[66],stage1_21[106],stage1_20[154]}
   );
   gpc606_5 gpc789 (
      {stage0_20[322], stage0_20[323], stage0_20[324], stage0_20[325], stage0_20[326], stage0_20[327]},
      {stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130], stage0_22[131]},
      {stage1_24[21],stage1_23[36],stage1_22[67],stage1_21[107],stage1_20[155]}
   );
   gpc606_5 gpc790 (
      {stage0_20[328], stage0_20[329], stage0_20[330], stage0_20[331], stage0_20[332], stage0_20[333]},
      {stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136], stage0_22[137]},
      {stage1_24[22],stage1_23[37],stage1_22[68],stage1_21[108],stage1_20[156]}
   );
   gpc606_5 gpc791 (
      {stage0_20[334], stage0_20[335], stage0_20[336], stage0_20[337], stage0_20[338], stage0_20[339]},
      {stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141], stage0_22[142], stage0_22[143]},
      {stage1_24[23],stage1_23[38],stage1_22[69],stage1_21[109],stage1_20[157]}
   );
   gpc606_5 gpc792 (
      {stage0_20[340], stage0_20[341], stage0_20[342], stage0_20[343], stage0_20[344], stage0_20[345]},
      {stage0_22[144], stage0_22[145], stage0_22[146], stage0_22[147], stage0_22[148], stage0_22[149]},
      {stage1_24[24],stage1_23[39],stage1_22[70],stage1_21[110],stage1_20[158]}
   );
   gpc606_5 gpc793 (
      {stage0_20[346], stage0_20[347], stage0_20[348], stage0_20[349], stage0_20[350], stage0_20[351]},
      {stage0_22[150], stage0_22[151], stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155]},
      {stage1_24[25],stage1_23[40],stage1_22[71],stage1_21[111],stage1_20[159]}
   );
   gpc606_5 gpc794 (
      {stage0_20[352], stage0_20[353], stage0_20[354], stage0_20[355], stage0_20[356], stage0_20[357]},
      {stage0_22[156], stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage1_24[26],stage1_23[41],stage1_22[72],stage1_21[112],stage1_20[160]}
   );
   gpc606_5 gpc795 (
      {stage0_20[358], stage0_20[359], stage0_20[360], stage0_20[361], stage0_20[362], stage0_20[363]},
      {stage0_22[162], stage0_22[163], stage0_22[164], stage0_22[165], stage0_22[166], stage0_22[167]},
      {stage1_24[27],stage1_23[42],stage1_22[73],stage1_21[113],stage1_20[161]}
   );
   gpc606_5 gpc796 (
      {stage0_20[364], stage0_20[365], stage0_20[366], stage0_20[367], stage0_20[368], stage0_20[369]},
      {stage0_22[168], stage0_22[169], stage0_22[170], stage0_22[171], stage0_22[172], stage0_22[173]},
      {stage1_24[28],stage1_23[43],stage1_22[74],stage1_21[114],stage1_20[162]}
   );
   gpc606_5 gpc797 (
      {stage0_20[370], stage0_20[371], stage0_20[372], stage0_20[373], stage0_20[374], stage0_20[375]},
      {stage0_22[174], stage0_22[175], stage0_22[176], stage0_22[177], stage0_22[178], stage0_22[179]},
      {stage1_24[29],stage1_23[44],stage1_22[75],stage1_21[115],stage1_20[163]}
   );
   gpc606_5 gpc798 (
      {stage0_20[376], stage0_20[377], stage0_20[378], stage0_20[379], stage0_20[380], stage0_20[381]},
      {stage0_22[180], stage0_22[181], stage0_22[182], stage0_22[183], stage0_22[184], stage0_22[185]},
      {stage1_24[30],stage1_23[45],stage1_22[76],stage1_21[116],stage1_20[164]}
   );
   gpc606_5 gpc799 (
      {stage0_20[382], stage0_20[383], stage0_20[384], stage0_20[385], stage0_20[386], stage0_20[387]},
      {stage0_22[186], stage0_22[187], stage0_22[188], stage0_22[189], stage0_22[190], stage0_22[191]},
      {stage1_24[31],stage1_23[46],stage1_22[77],stage1_21[117],stage1_20[165]}
   );
   gpc606_5 gpc800 (
      {stage0_20[388], stage0_20[389], stage0_20[390], stage0_20[391], stage0_20[392], stage0_20[393]},
      {stage0_22[192], stage0_22[193], stage0_22[194], stage0_22[195], stage0_22[196], stage0_22[197]},
      {stage1_24[32],stage1_23[47],stage1_22[78],stage1_21[118],stage1_20[166]}
   );
   gpc606_5 gpc801 (
      {stage0_20[394], stage0_20[395], stage0_20[396], stage0_20[397], stage0_20[398], stage0_20[399]},
      {stage0_22[198], stage0_22[199], stage0_22[200], stage0_22[201], stage0_22[202], stage0_22[203]},
      {stage1_24[33],stage1_23[48],stage1_22[79],stage1_21[119],stage1_20[167]}
   );
   gpc606_5 gpc802 (
      {stage0_20[400], stage0_20[401], stage0_20[402], stage0_20[403], stage0_20[404], stage0_20[405]},
      {stage0_22[204], stage0_22[205], stage0_22[206], stage0_22[207], stage0_22[208], stage0_22[209]},
      {stage1_24[34],stage1_23[49],stage1_22[80],stage1_21[120],stage1_20[168]}
   );
   gpc606_5 gpc803 (
      {stage0_20[406], stage0_20[407], stage0_20[408], stage0_20[409], stage0_20[410], stage0_20[411]},
      {stage0_22[210], stage0_22[211], stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215]},
      {stage1_24[35],stage1_23[50],stage1_22[81],stage1_21[121],stage1_20[169]}
   );
   gpc606_5 gpc804 (
      {stage0_20[412], stage0_20[413], stage0_20[414], stage0_20[415], stage0_20[416], stage0_20[417]},
      {stage0_22[216], stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage1_24[36],stage1_23[51],stage1_22[82],stage1_21[122],stage1_20[170]}
   );
   gpc606_5 gpc805 (
      {stage0_20[418], stage0_20[419], stage0_20[420], stage0_20[421], stage0_20[422], stage0_20[423]},
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226], stage0_22[227]},
      {stage1_24[37],stage1_23[52],stage1_22[83],stage1_21[123],stage1_20[171]}
   );
   gpc606_5 gpc806 (
      {stage0_20[424], stage0_20[425], stage0_20[426], stage0_20[427], stage0_20[428], stage0_20[429]},
      {stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231], stage0_22[232], stage0_22[233]},
      {stage1_24[38],stage1_23[53],stage1_22[84],stage1_21[124],stage1_20[172]}
   );
   gpc606_5 gpc807 (
      {stage0_20[430], stage0_20[431], stage0_20[432], stage0_20[433], stage0_20[434], stage0_20[435]},
      {stage0_22[234], stage0_22[235], stage0_22[236], stage0_22[237], stage0_22[238], stage0_22[239]},
      {stage1_24[39],stage1_23[54],stage1_22[85],stage1_21[125],stage1_20[173]}
   );
   gpc606_5 gpc808 (
      {stage0_20[436], stage0_20[437], stage0_20[438], stage0_20[439], stage0_20[440], stage0_20[441]},
      {stage0_22[240], stage0_22[241], stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245]},
      {stage1_24[40],stage1_23[55],stage1_22[86],stage1_21[126],stage1_20[174]}
   );
   gpc606_5 gpc809 (
      {stage0_20[442], stage0_20[443], stage0_20[444], stage0_20[445], stage0_20[446], stage0_20[447]},
      {stage0_22[246], stage0_22[247], stage0_22[248], stage0_22[249], stage0_22[250], stage0_22[251]},
      {stage1_24[41],stage1_23[56],stage1_22[87],stage1_21[127],stage1_20[175]}
   );
   gpc606_5 gpc810 (
      {stage0_20[448], stage0_20[449], stage0_20[450], stage0_20[451], stage0_20[452], stage0_20[453]},
      {stage0_22[252], stage0_22[253], stage0_22[254], stage0_22[255], stage0_22[256], stage0_22[257]},
      {stage1_24[42],stage1_23[57],stage1_22[88],stage1_21[128],stage1_20[176]}
   );
   gpc606_5 gpc811 (
      {stage0_20[454], stage0_20[455], stage0_20[456], stage0_20[457], stage0_20[458], stage0_20[459]},
      {stage0_22[258], stage0_22[259], stage0_22[260], stage0_22[261], stage0_22[262], stage0_22[263]},
      {stage1_24[43],stage1_23[58],stage1_22[89],stage1_21[129],stage1_20[177]}
   );
   gpc606_5 gpc812 (
      {stage0_20[460], stage0_20[461], stage0_20[462], stage0_20[463], stage0_20[464], stage0_20[465]},
      {stage0_22[264], stage0_22[265], stage0_22[266], stage0_22[267], stage0_22[268], stage0_22[269]},
      {stage1_24[44],stage1_23[59],stage1_22[90],stage1_21[130],stage1_20[178]}
   );
   gpc606_5 gpc813 (
      {stage0_20[466], stage0_20[467], stage0_20[468], stage0_20[469], stage0_20[470], stage0_20[471]},
      {stage0_22[270], stage0_22[271], stage0_22[272], stage0_22[273], stage0_22[274], stage0_22[275]},
      {stage1_24[45],stage1_23[60],stage1_22[91],stage1_21[131],stage1_20[179]}
   );
   gpc606_5 gpc814 (
      {stage0_20[472], stage0_20[473], stage0_20[474], stage0_20[475], stage0_20[476], stage0_20[477]},
      {stage0_22[276], stage0_22[277], stage0_22[278], stage0_22[279], stage0_22[280], stage0_22[281]},
      {stage1_24[46],stage1_23[61],stage1_22[92],stage1_21[132],stage1_20[180]}
   );
   gpc606_5 gpc815 (
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[47],stage1_23[62],stage1_22[93],stage1_21[133]}
   );
   gpc606_5 gpc816 (
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[48],stage1_23[63],stage1_22[94],stage1_21[134]}
   );
   gpc606_5 gpc817 (
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[49],stage1_23[64],stage1_22[95],stage1_21[135]}
   );
   gpc606_5 gpc818 (
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[50],stage1_23[65],stage1_22[96],stage1_21[136]}
   );
   gpc606_5 gpc819 (
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[51],stage1_23[66],stage1_22[97],stage1_21[137]}
   );
   gpc606_5 gpc820 (
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[52],stage1_23[67],stage1_22[98],stage1_21[138]}
   );
   gpc606_5 gpc821 (
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[53],stage1_23[68],stage1_22[99],stage1_21[139]}
   );
   gpc606_5 gpc822 (
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[54],stage1_23[69],stage1_22[100],stage1_21[140]}
   );
   gpc606_5 gpc823 (
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[55],stage1_23[70],stage1_22[101],stage1_21[141]}
   );
   gpc606_5 gpc824 (
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[56],stage1_23[71],stage1_22[102],stage1_21[142]}
   );
   gpc606_5 gpc825 (
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[57],stage1_23[72],stage1_22[103],stage1_21[143]}
   );
   gpc606_5 gpc826 (
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[58],stage1_23[73],stage1_22[104],stage1_21[144]}
   );
   gpc606_5 gpc827 (
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[59],stage1_23[74],stage1_22[105],stage1_21[145]}
   );
   gpc606_5 gpc828 (
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[60],stage1_23[75],stage1_22[106],stage1_21[146]}
   );
   gpc606_5 gpc829 (
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[61],stage1_23[76],stage1_22[107],stage1_21[147]}
   );
   gpc606_5 gpc830 (
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[62],stage1_23[77],stage1_22[108],stage1_21[148]}
   );
   gpc606_5 gpc831 (
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[63],stage1_23[78],stage1_22[109],stage1_21[149]}
   );
   gpc606_5 gpc832 (
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage0_23[102], stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107]},
      {stage1_25[17],stage1_24[64],stage1_23[79],stage1_22[110],stage1_21[150]}
   );
   gpc606_5 gpc833 (
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage0_23[108], stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113]},
      {stage1_25[18],stage1_24[65],stage1_23[80],stage1_22[111],stage1_21[151]}
   );
   gpc606_5 gpc834 (
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage0_23[114], stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119]},
      {stage1_25[19],stage1_24[66],stage1_23[81],stage1_22[112],stage1_21[152]}
   );
   gpc606_5 gpc835 (
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage0_23[120], stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage1_25[20],stage1_24[67],stage1_23[82],stage1_22[113],stage1_21[153]}
   );
   gpc606_5 gpc836 (
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage0_23[126], stage0_23[127], stage0_23[128], stage0_23[129], stage0_23[130], stage0_23[131]},
      {stage1_25[21],stage1_24[68],stage1_23[83],stage1_22[114],stage1_21[154]}
   );
   gpc606_5 gpc837 (
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage0_23[132], stage0_23[133], stage0_23[134], stage0_23[135], stage0_23[136], stage0_23[137]},
      {stage1_25[22],stage1_24[69],stage1_23[84],stage1_22[115],stage1_21[155]}
   );
   gpc606_5 gpc838 (
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage0_23[138], stage0_23[139], stage0_23[140], stage0_23[141], stage0_23[142], stage0_23[143]},
      {stage1_25[23],stage1_24[70],stage1_23[85],stage1_22[116],stage1_21[156]}
   );
   gpc606_5 gpc839 (
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage0_23[144], stage0_23[145], stage0_23[146], stage0_23[147], stage0_23[148], stage0_23[149]},
      {stage1_25[24],stage1_24[71],stage1_23[86],stage1_22[117],stage1_21[157]}
   );
   gpc606_5 gpc840 (
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage1_25[25],stage1_24[72],stage1_23[87],stage1_22[118],stage1_21[158]}
   );
   gpc606_5 gpc841 (
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249], stage0_21[250], stage0_21[251]},
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160], stage0_23[161]},
      {stage1_25[26],stage1_24[73],stage1_23[88],stage1_22[119],stage1_21[159]}
   );
   gpc606_5 gpc842 (
      {stage0_21[252], stage0_21[253], stage0_21[254], stage0_21[255], stage0_21[256], stage0_21[257]},
      {stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165], stage0_23[166], stage0_23[167]},
      {stage1_25[27],stage1_24[74],stage1_23[89],stage1_22[120],stage1_21[160]}
   );
   gpc606_5 gpc843 (
      {stage0_21[258], stage0_21[259], stage0_21[260], stage0_21[261], stage0_21[262], stage0_21[263]},
      {stage0_23[168], stage0_23[169], stage0_23[170], stage0_23[171], stage0_23[172], stage0_23[173]},
      {stage1_25[28],stage1_24[75],stage1_23[90],stage1_22[121],stage1_21[161]}
   );
   gpc606_5 gpc844 (
      {stage0_21[264], stage0_21[265], stage0_21[266], stage0_21[267], stage0_21[268], stage0_21[269]},
      {stage0_23[174], stage0_23[175], stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179]},
      {stage1_25[29],stage1_24[76],stage1_23[91],stage1_22[122],stage1_21[162]}
   );
   gpc606_5 gpc845 (
      {stage0_21[270], stage0_21[271], stage0_21[272], stage0_21[273], stage0_21[274], stage0_21[275]},
      {stage0_23[180], stage0_23[181], stage0_23[182], stage0_23[183], stage0_23[184], stage0_23[185]},
      {stage1_25[30],stage1_24[77],stage1_23[92],stage1_22[123],stage1_21[163]}
   );
   gpc606_5 gpc846 (
      {stage0_21[276], stage0_21[277], stage0_21[278], stage0_21[279], stage0_21[280], stage0_21[281]},
      {stage0_23[186], stage0_23[187], stage0_23[188], stage0_23[189], stage0_23[190], stage0_23[191]},
      {stage1_25[31],stage1_24[78],stage1_23[93],stage1_22[124],stage1_21[164]}
   );
   gpc606_5 gpc847 (
      {stage0_21[282], stage0_21[283], stage0_21[284], stage0_21[285], stage0_21[286], stage0_21[287]},
      {stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195], stage0_23[196], stage0_23[197]},
      {stage1_25[32],stage1_24[79],stage1_23[94],stage1_22[125],stage1_21[165]}
   );
   gpc606_5 gpc848 (
      {stage0_21[288], stage0_21[289], stage0_21[290], stage0_21[291], stage0_21[292], stage0_21[293]},
      {stage0_23[198], stage0_23[199], stage0_23[200], stage0_23[201], stage0_23[202], stage0_23[203]},
      {stage1_25[33],stage1_24[80],stage1_23[95],stage1_22[126],stage1_21[166]}
   );
   gpc606_5 gpc849 (
      {stage0_21[294], stage0_21[295], stage0_21[296], stage0_21[297], stage0_21[298], stage0_21[299]},
      {stage0_23[204], stage0_23[205], stage0_23[206], stage0_23[207], stage0_23[208], stage0_23[209]},
      {stage1_25[34],stage1_24[81],stage1_23[96],stage1_22[127],stage1_21[167]}
   );
   gpc606_5 gpc850 (
      {stage0_21[300], stage0_21[301], stage0_21[302], stage0_21[303], stage0_21[304], stage0_21[305]},
      {stage0_23[210], stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214], stage0_23[215]},
      {stage1_25[35],stage1_24[82],stage1_23[97],stage1_22[128],stage1_21[168]}
   );
   gpc606_5 gpc851 (
      {stage0_21[306], stage0_21[307], stage0_21[308], stage0_21[309], stage0_21[310], stage0_21[311]},
      {stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220], stage0_23[221]},
      {stage1_25[36],stage1_24[83],stage1_23[98],stage1_22[129],stage1_21[169]}
   );
   gpc606_5 gpc852 (
      {stage0_21[312], stage0_21[313], stage0_21[314], stage0_21[315], stage0_21[316], stage0_21[317]},
      {stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225], stage0_23[226], stage0_23[227]},
      {stage1_25[37],stage1_24[84],stage1_23[99],stage1_22[130],stage1_21[170]}
   );
   gpc606_5 gpc853 (
      {stage0_21[318], stage0_21[319], stage0_21[320], stage0_21[321], stage0_21[322], stage0_21[323]},
      {stage0_23[228], stage0_23[229], stage0_23[230], stage0_23[231], stage0_23[232], stage0_23[233]},
      {stage1_25[38],stage1_24[85],stage1_23[100],stage1_22[131],stage1_21[171]}
   );
   gpc606_5 gpc854 (
      {stage0_21[324], stage0_21[325], stage0_21[326], stage0_21[327], stage0_21[328], stage0_21[329]},
      {stage0_23[234], stage0_23[235], stage0_23[236], stage0_23[237], stage0_23[238], stage0_23[239]},
      {stage1_25[39],stage1_24[86],stage1_23[101],stage1_22[132],stage1_21[172]}
   );
   gpc606_5 gpc855 (
      {stage0_21[330], stage0_21[331], stage0_21[332], stage0_21[333], stage0_21[334], stage0_21[335]},
      {stage0_23[240], stage0_23[241], stage0_23[242], stage0_23[243], stage0_23[244], stage0_23[245]},
      {stage1_25[40],stage1_24[87],stage1_23[102],stage1_22[133],stage1_21[173]}
   );
   gpc606_5 gpc856 (
      {stage0_21[336], stage0_21[337], stage0_21[338], stage0_21[339], stage0_21[340], stage0_21[341]},
      {stage0_23[246], stage0_23[247], stage0_23[248], stage0_23[249], stage0_23[250], stage0_23[251]},
      {stage1_25[41],stage1_24[88],stage1_23[103],stage1_22[134],stage1_21[174]}
   );
   gpc606_5 gpc857 (
      {stage0_21[342], stage0_21[343], stage0_21[344], stage0_21[345], stage0_21[346], stage0_21[347]},
      {stage0_23[252], stage0_23[253], stage0_23[254], stage0_23[255], stage0_23[256], stage0_23[257]},
      {stage1_25[42],stage1_24[89],stage1_23[104],stage1_22[135],stage1_21[175]}
   );
   gpc606_5 gpc858 (
      {stage0_21[348], stage0_21[349], stage0_21[350], stage0_21[351], stage0_21[352], stage0_21[353]},
      {stage0_23[258], stage0_23[259], stage0_23[260], stage0_23[261], stage0_23[262], stage0_23[263]},
      {stage1_25[43],stage1_24[90],stage1_23[105],stage1_22[136],stage1_21[176]}
   );
   gpc606_5 gpc859 (
      {stage0_21[354], stage0_21[355], stage0_21[356], stage0_21[357], stage0_21[358], stage0_21[359]},
      {stage0_23[264], stage0_23[265], stage0_23[266], stage0_23[267], stage0_23[268], stage0_23[269]},
      {stage1_25[44],stage1_24[91],stage1_23[106],stage1_22[137],stage1_21[177]}
   );
   gpc606_5 gpc860 (
      {stage0_21[360], stage0_21[361], stage0_21[362], stage0_21[363], stage0_21[364], stage0_21[365]},
      {stage0_23[270], stage0_23[271], stage0_23[272], stage0_23[273], stage0_23[274], stage0_23[275]},
      {stage1_25[45],stage1_24[92],stage1_23[107],stage1_22[138],stage1_21[178]}
   );
   gpc606_5 gpc861 (
      {stage0_21[366], stage0_21[367], stage0_21[368], stage0_21[369], stage0_21[370], stage0_21[371]},
      {stage0_23[276], stage0_23[277], stage0_23[278], stage0_23[279], stage0_23[280], stage0_23[281]},
      {stage1_25[46],stage1_24[93],stage1_23[108],stage1_22[139],stage1_21[179]}
   );
   gpc606_5 gpc862 (
      {stage0_21[372], stage0_21[373], stage0_21[374], stage0_21[375], stage0_21[376], stage0_21[377]},
      {stage0_23[282], stage0_23[283], stage0_23[284], stage0_23[285], stage0_23[286], stage0_23[287]},
      {stage1_25[47],stage1_24[94],stage1_23[109],stage1_22[140],stage1_21[180]}
   );
   gpc606_5 gpc863 (
      {stage0_21[378], stage0_21[379], stage0_21[380], stage0_21[381], stage0_21[382], stage0_21[383]},
      {stage0_23[288], stage0_23[289], stage0_23[290], stage0_23[291], stage0_23[292], stage0_23[293]},
      {stage1_25[48],stage1_24[95],stage1_23[110],stage1_22[141],stage1_21[181]}
   );
   gpc606_5 gpc864 (
      {stage0_21[384], stage0_21[385], stage0_21[386], stage0_21[387], stage0_21[388], stage0_21[389]},
      {stage0_23[294], stage0_23[295], stage0_23[296], stage0_23[297], stage0_23[298], stage0_23[299]},
      {stage1_25[49],stage1_24[96],stage1_23[111],stage1_22[142],stage1_21[182]}
   );
   gpc606_5 gpc865 (
      {stage0_21[390], stage0_21[391], stage0_21[392], stage0_21[393], stage0_21[394], stage0_21[395]},
      {stage0_23[300], stage0_23[301], stage0_23[302], stage0_23[303], stage0_23[304], stage0_23[305]},
      {stage1_25[50],stage1_24[97],stage1_23[112],stage1_22[143],stage1_21[183]}
   );
   gpc606_5 gpc866 (
      {stage0_21[396], stage0_21[397], stage0_21[398], stage0_21[399], stage0_21[400], stage0_21[401]},
      {stage0_23[306], stage0_23[307], stage0_23[308], stage0_23[309], stage0_23[310], stage0_23[311]},
      {stage1_25[51],stage1_24[98],stage1_23[113],stage1_22[144],stage1_21[184]}
   );
   gpc606_5 gpc867 (
      {stage0_21[402], stage0_21[403], stage0_21[404], stage0_21[405], stage0_21[406], stage0_21[407]},
      {stage0_23[312], stage0_23[313], stage0_23[314], stage0_23[315], stage0_23[316], stage0_23[317]},
      {stage1_25[52],stage1_24[99],stage1_23[114],stage1_22[145],stage1_21[185]}
   );
   gpc606_5 gpc868 (
      {stage0_21[408], stage0_21[409], stage0_21[410], stage0_21[411], stage0_21[412], stage0_21[413]},
      {stage0_23[318], stage0_23[319], stage0_23[320], stage0_23[321], stage0_23[322], stage0_23[323]},
      {stage1_25[53],stage1_24[100],stage1_23[115],stage1_22[146],stage1_21[186]}
   );
   gpc606_5 gpc869 (
      {stage0_21[414], stage0_21[415], stage0_21[416], stage0_21[417], stage0_21[418], stage0_21[419]},
      {stage0_23[324], stage0_23[325], stage0_23[326], stage0_23[327], stage0_23[328], stage0_23[329]},
      {stage1_25[54],stage1_24[101],stage1_23[116],stage1_22[147],stage1_21[187]}
   );
   gpc606_5 gpc870 (
      {stage0_21[420], stage0_21[421], stage0_21[422], stage0_21[423], stage0_21[424], stage0_21[425]},
      {stage0_23[330], stage0_23[331], stage0_23[332], stage0_23[333], stage0_23[334], stage0_23[335]},
      {stage1_25[55],stage1_24[102],stage1_23[117],stage1_22[148],stage1_21[188]}
   );
   gpc606_5 gpc871 (
      {stage0_21[426], stage0_21[427], stage0_21[428], stage0_21[429], stage0_21[430], stage0_21[431]},
      {stage0_23[336], stage0_23[337], stage0_23[338], stage0_23[339], stage0_23[340], stage0_23[341]},
      {stage1_25[56],stage1_24[103],stage1_23[118],stage1_22[149],stage1_21[189]}
   );
   gpc606_5 gpc872 (
      {stage0_21[432], stage0_21[433], stage0_21[434], stage0_21[435], stage0_21[436], stage0_21[437]},
      {stage0_23[342], stage0_23[343], stage0_23[344], stage0_23[345], stage0_23[346], stage0_23[347]},
      {stage1_25[57],stage1_24[104],stage1_23[119],stage1_22[150],stage1_21[190]}
   );
   gpc606_5 gpc873 (
      {stage0_21[438], stage0_21[439], stage0_21[440], stage0_21[441], stage0_21[442], stage0_21[443]},
      {stage0_23[348], stage0_23[349], stage0_23[350], stage0_23[351], stage0_23[352], stage0_23[353]},
      {stage1_25[58],stage1_24[105],stage1_23[120],stage1_22[151],stage1_21[191]}
   );
   gpc606_5 gpc874 (
      {stage0_21[444], stage0_21[445], stage0_21[446], stage0_21[447], stage0_21[448], stage0_21[449]},
      {stage0_23[354], stage0_23[355], stage0_23[356], stage0_23[357], stage0_23[358], stage0_23[359]},
      {stage1_25[59],stage1_24[106],stage1_23[121],stage1_22[152],stage1_21[192]}
   );
   gpc606_5 gpc875 (
      {stage0_21[450], stage0_21[451], stage0_21[452], stage0_21[453], stage0_21[454], stage0_21[455]},
      {stage0_23[360], stage0_23[361], stage0_23[362], stage0_23[363], stage0_23[364], stage0_23[365]},
      {stage1_25[60],stage1_24[107],stage1_23[122],stage1_22[153],stage1_21[193]}
   );
   gpc606_5 gpc876 (
      {stage0_21[456], stage0_21[457], stage0_21[458], stage0_21[459], stage0_21[460], stage0_21[461]},
      {stage0_23[366], stage0_23[367], stage0_23[368], stage0_23[369], stage0_23[370], stage0_23[371]},
      {stage1_25[61],stage1_24[108],stage1_23[123],stage1_22[154],stage1_21[194]}
   );
   gpc606_5 gpc877 (
      {stage0_21[462], stage0_21[463], stage0_21[464], stage0_21[465], stage0_21[466], stage0_21[467]},
      {stage0_23[372], stage0_23[373], stage0_23[374], stage0_23[375], stage0_23[376], stage0_23[377]},
      {stage1_25[62],stage1_24[109],stage1_23[124],stage1_22[155],stage1_21[195]}
   );
   gpc606_5 gpc878 (
      {stage0_21[468], stage0_21[469], stage0_21[470], stage0_21[471], stage0_21[472], stage0_21[473]},
      {stage0_23[378], stage0_23[379], stage0_23[380], stage0_23[381], stage0_23[382], stage0_23[383]},
      {stage1_25[63],stage1_24[110],stage1_23[125],stage1_22[156],stage1_21[196]}
   );
   gpc606_5 gpc879 (
      {stage0_21[474], stage0_21[475], stage0_21[476], stage0_21[477], stage0_21[478], stage0_21[479]},
      {stage0_23[384], stage0_23[385], stage0_23[386], stage0_23[387], stage0_23[388], stage0_23[389]},
      {stage1_25[64],stage1_24[111],stage1_23[126],stage1_22[157],stage1_21[197]}
   );
   gpc606_5 gpc880 (
      {stage0_21[480], stage0_21[481], stage0_21[482], stage0_21[483], stage0_21[484], stage0_21[485]},
      {stage0_23[390], stage0_23[391], stage0_23[392], stage0_23[393], stage0_23[394], stage0_23[395]},
      {stage1_25[65],stage1_24[112],stage1_23[127],stage1_22[158],stage1_21[198]}
   );
   gpc615_5 gpc881 (
      {stage0_22[282], stage0_22[283], stage0_22[284], stage0_22[285], stage0_22[286]},
      {stage0_23[396]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[66],stage1_24[113],stage1_23[128],stage1_22[159]}
   );
   gpc615_5 gpc882 (
      {stage0_22[287], stage0_22[288], stage0_22[289], stage0_22[290], stage0_22[291]},
      {stage0_23[397]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[67],stage1_24[114],stage1_23[129],stage1_22[160]}
   );
   gpc615_5 gpc883 (
      {stage0_22[292], stage0_22[293], stage0_22[294], stage0_22[295], stage0_22[296]},
      {stage0_23[398]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[68],stage1_24[115],stage1_23[130],stage1_22[161]}
   );
   gpc615_5 gpc884 (
      {stage0_22[297], stage0_22[298], stage0_22[299], stage0_22[300], stage0_22[301]},
      {stage0_23[399]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[69],stage1_24[116],stage1_23[131],stage1_22[162]}
   );
   gpc615_5 gpc885 (
      {stage0_22[302], stage0_22[303], stage0_22[304], stage0_22[305], stage0_22[306]},
      {stage0_23[400]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[70],stage1_24[117],stage1_23[132],stage1_22[163]}
   );
   gpc615_5 gpc886 (
      {stage0_22[307], stage0_22[308], stage0_22[309], stage0_22[310], stage0_22[311]},
      {stage0_23[401]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[71],stage1_24[118],stage1_23[133],stage1_22[164]}
   );
   gpc615_5 gpc887 (
      {stage0_22[312], stage0_22[313], stage0_22[314], stage0_22[315], stage0_22[316]},
      {stage0_23[402]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[72],stage1_24[119],stage1_23[134],stage1_22[165]}
   );
   gpc615_5 gpc888 (
      {stage0_22[317], stage0_22[318], stage0_22[319], stage0_22[320], stage0_22[321]},
      {stage0_23[403]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[73],stage1_24[120],stage1_23[135],stage1_22[166]}
   );
   gpc615_5 gpc889 (
      {stage0_22[322], stage0_22[323], stage0_22[324], stage0_22[325], stage0_22[326]},
      {stage0_23[404]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[74],stage1_24[121],stage1_23[136],stage1_22[167]}
   );
   gpc615_5 gpc890 (
      {stage0_22[327], stage0_22[328], stage0_22[329], stage0_22[330], stage0_22[331]},
      {stage0_23[405]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[75],stage1_24[122],stage1_23[137],stage1_22[168]}
   );
   gpc615_5 gpc891 (
      {stage0_22[332], stage0_22[333], stage0_22[334], stage0_22[335], stage0_22[336]},
      {stage0_23[406]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[76],stage1_24[123],stage1_23[138],stage1_22[169]}
   );
   gpc615_5 gpc892 (
      {stage0_22[337], stage0_22[338], stage0_22[339], stage0_22[340], stage0_22[341]},
      {stage0_23[407]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[77],stage1_24[124],stage1_23[139],stage1_22[170]}
   );
   gpc615_5 gpc893 (
      {stage0_22[342], stage0_22[343], stage0_22[344], stage0_22[345], stage0_22[346]},
      {stage0_23[408]},
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage1_26[12],stage1_25[78],stage1_24[125],stage1_23[140],stage1_22[171]}
   );
   gpc615_5 gpc894 (
      {stage0_22[347], stage0_22[348], stage0_22[349], stage0_22[350], stage0_22[351]},
      {stage0_23[409]},
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage1_26[13],stage1_25[79],stage1_24[126],stage1_23[141],stage1_22[172]}
   );
   gpc615_5 gpc895 (
      {stage0_22[352], stage0_22[353], stage0_22[354], stage0_22[355], stage0_22[356]},
      {stage0_23[410]},
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage1_26[14],stage1_25[80],stage1_24[127],stage1_23[142],stage1_22[173]}
   );
   gpc615_5 gpc896 (
      {stage0_22[357], stage0_22[358], stage0_22[359], stage0_22[360], stage0_22[361]},
      {stage0_23[411]},
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage1_26[15],stage1_25[81],stage1_24[128],stage1_23[143],stage1_22[174]}
   );
   gpc615_5 gpc897 (
      {stage0_22[362], stage0_22[363], stage0_22[364], stage0_22[365], stage0_22[366]},
      {stage0_23[412]},
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage1_26[16],stage1_25[82],stage1_24[129],stage1_23[144],stage1_22[175]}
   );
   gpc615_5 gpc898 (
      {stage0_22[367], stage0_22[368], stage0_22[369], stage0_22[370], stage0_22[371]},
      {stage0_23[413]},
      {stage0_24[102], stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107]},
      {stage1_26[17],stage1_25[83],stage1_24[130],stage1_23[145],stage1_22[176]}
   );
   gpc615_5 gpc899 (
      {stage0_22[372], stage0_22[373], stage0_22[374], stage0_22[375], stage0_22[376]},
      {stage0_23[414]},
      {stage0_24[108], stage0_24[109], stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113]},
      {stage1_26[18],stage1_25[84],stage1_24[131],stage1_23[146],stage1_22[177]}
   );
   gpc615_5 gpc900 (
      {stage0_22[377], stage0_22[378], stage0_22[379], stage0_22[380], stage0_22[381]},
      {stage0_23[415]},
      {stage0_24[114], stage0_24[115], stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119]},
      {stage1_26[19],stage1_25[85],stage1_24[132],stage1_23[147],stage1_22[178]}
   );
   gpc615_5 gpc901 (
      {stage0_22[382], stage0_22[383], stage0_22[384], stage0_22[385], stage0_22[386]},
      {stage0_23[416]},
      {stage0_24[120], stage0_24[121], stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125]},
      {stage1_26[20],stage1_25[86],stage1_24[133],stage1_23[148],stage1_22[179]}
   );
   gpc615_5 gpc902 (
      {stage0_22[387], stage0_22[388], stage0_22[389], stage0_22[390], stage0_22[391]},
      {stage0_23[417]},
      {stage0_24[126], stage0_24[127], stage0_24[128], stage0_24[129], stage0_24[130], stage0_24[131]},
      {stage1_26[21],stage1_25[87],stage1_24[134],stage1_23[149],stage1_22[180]}
   );
   gpc615_5 gpc903 (
      {stage0_22[392], stage0_22[393], stage0_22[394], stage0_22[395], stage0_22[396]},
      {stage0_23[418]},
      {stage0_24[132], stage0_24[133], stage0_24[134], stage0_24[135], stage0_24[136], stage0_24[137]},
      {stage1_26[22],stage1_25[88],stage1_24[135],stage1_23[150],stage1_22[181]}
   );
   gpc615_5 gpc904 (
      {stage0_22[397], stage0_22[398], stage0_22[399], stage0_22[400], stage0_22[401]},
      {stage0_23[419]},
      {stage0_24[138], stage0_24[139], stage0_24[140], stage0_24[141], stage0_24[142], stage0_24[143]},
      {stage1_26[23],stage1_25[89],stage1_24[136],stage1_23[151],stage1_22[182]}
   );
   gpc615_5 gpc905 (
      {stage0_22[402], stage0_22[403], stage0_22[404], stage0_22[405], stage0_22[406]},
      {stage0_23[420]},
      {stage0_24[144], stage0_24[145], stage0_24[146], stage0_24[147], stage0_24[148], stage0_24[149]},
      {stage1_26[24],stage1_25[90],stage1_24[137],stage1_23[152],stage1_22[183]}
   );
   gpc615_5 gpc906 (
      {stage0_22[407], stage0_22[408], stage0_22[409], stage0_22[410], stage0_22[411]},
      {stage0_23[421]},
      {stage0_24[150], stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154], stage0_24[155]},
      {stage1_26[25],stage1_25[91],stage1_24[138],stage1_23[153],stage1_22[184]}
   );
   gpc615_5 gpc907 (
      {stage0_22[412], stage0_22[413], stage0_22[414], stage0_22[415], stage0_22[416]},
      {stage0_23[422]},
      {stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160], stage0_24[161]},
      {stage1_26[26],stage1_25[92],stage1_24[139],stage1_23[154],stage1_22[185]}
   );
   gpc615_5 gpc908 (
      {stage0_22[417], stage0_22[418], stage0_22[419], stage0_22[420], stage0_22[421]},
      {stage0_23[423]},
      {stage0_24[162], stage0_24[163], stage0_24[164], stage0_24[165], stage0_24[166], stage0_24[167]},
      {stage1_26[27],stage1_25[93],stage1_24[140],stage1_23[155],stage1_22[186]}
   );
   gpc615_5 gpc909 (
      {stage0_23[424], stage0_23[425], stage0_23[426], stage0_23[427], stage0_23[428]},
      {stage0_24[168]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[28],stage1_25[94],stage1_24[141],stage1_23[156]}
   );
   gpc615_5 gpc910 (
      {stage0_23[429], stage0_23[430], stage0_23[431], stage0_23[432], stage0_23[433]},
      {stage0_24[169]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[29],stage1_25[95],stage1_24[142],stage1_23[157]}
   );
   gpc615_5 gpc911 (
      {stage0_23[434], stage0_23[435], stage0_23[436], stage0_23[437], stage0_23[438]},
      {stage0_24[170]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[30],stage1_25[96],stage1_24[143],stage1_23[158]}
   );
   gpc615_5 gpc912 (
      {stage0_23[439], stage0_23[440], stage0_23[441], stage0_23[442], stage0_23[443]},
      {stage0_24[171]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[31],stage1_25[97],stage1_24[144],stage1_23[159]}
   );
   gpc615_5 gpc913 (
      {stage0_23[444], stage0_23[445], stage0_23[446], stage0_23[447], stage0_23[448]},
      {stage0_24[172]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[32],stage1_25[98],stage1_24[145],stage1_23[160]}
   );
   gpc615_5 gpc914 (
      {stage0_23[449], stage0_23[450], stage0_23[451], stage0_23[452], stage0_23[453]},
      {stage0_24[173]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[33],stage1_25[99],stage1_24[146],stage1_23[161]}
   );
   gpc615_5 gpc915 (
      {stage0_23[454], stage0_23[455], stage0_23[456], stage0_23[457], stage0_23[458]},
      {stage0_24[174]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[34],stage1_25[100],stage1_24[147],stage1_23[162]}
   );
   gpc615_5 gpc916 (
      {stage0_23[459], stage0_23[460], stage0_23[461], stage0_23[462], stage0_23[463]},
      {stage0_24[175]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[35],stage1_25[101],stage1_24[148],stage1_23[163]}
   );
   gpc615_5 gpc917 (
      {stage0_23[464], stage0_23[465], stage0_23[466], stage0_23[467], stage0_23[468]},
      {stage0_24[176]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[36],stage1_25[102],stage1_24[149],stage1_23[164]}
   );
   gpc615_5 gpc918 (
      {stage0_23[469], stage0_23[470], stage0_23[471], stage0_23[472], stage0_23[473]},
      {stage0_24[177]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[37],stage1_25[103],stage1_24[150],stage1_23[165]}
   );
   gpc606_5 gpc919 (
      {stage0_24[178], stage0_24[179], stage0_24[180], stage0_24[181], stage0_24[182], stage0_24[183]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[10],stage1_26[38],stage1_25[104],stage1_24[151]}
   );
   gpc606_5 gpc920 (
      {stage0_24[184], stage0_24[185], stage0_24[186], stage0_24[187], stage0_24[188], stage0_24[189]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[11],stage1_26[39],stage1_25[105],stage1_24[152]}
   );
   gpc606_5 gpc921 (
      {stage0_24[190], stage0_24[191], stage0_24[192], stage0_24[193], stage0_24[194], stage0_24[195]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[12],stage1_26[40],stage1_25[106],stage1_24[153]}
   );
   gpc615_5 gpc922 (
      {stage0_24[196], stage0_24[197], stage0_24[198], stage0_24[199], stage0_24[200]},
      {stage0_25[60]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[13],stage1_26[41],stage1_25[107],stage1_24[154]}
   );
   gpc615_5 gpc923 (
      {stage0_24[201], stage0_24[202], stage0_24[203], stage0_24[204], stage0_24[205]},
      {stage0_25[61]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[14],stage1_26[42],stage1_25[108],stage1_24[155]}
   );
   gpc615_5 gpc924 (
      {stage0_24[206], stage0_24[207], stage0_24[208], stage0_24[209], stage0_24[210]},
      {stage0_25[62]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[15],stage1_26[43],stage1_25[109],stage1_24[156]}
   );
   gpc615_5 gpc925 (
      {stage0_24[211], stage0_24[212], stage0_24[213], stage0_24[214], stage0_24[215]},
      {stage0_25[63]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[16],stage1_26[44],stage1_25[110],stage1_24[157]}
   );
   gpc615_5 gpc926 (
      {stage0_24[216], stage0_24[217], stage0_24[218], stage0_24[219], stage0_24[220]},
      {stage0_25[64]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[17],stage1_26[45],stage1_25[111],stage1_24[158]}
   );
   gpc615_5 gpc927 (
      {stage0_24[221], stage0_24[222], stage0_24[223], stage0_24[224], stage0_24[225]},
      {stage0_25[65]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[18],stage1_26[46],stage1_25[112],stage1_24[159]}
   );
   gpc615_5 gpc928 (
      {stage0_24[226], stage0_24[227], stage0_24[228], stage0_24[229], stage0_24[230]},
      {stage0_25[66]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[19],stage1_26[47],stage1_25[113],stage1_24[160]}
   );
   gpc615_5 gpc929 (
      {stage0_24[231], stage0_24[232], stage0_24[233], stage0_24[234], stage0_24[235]},
      {stage0_25[67]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[20],stage1_26[48],stage1_25[114],stage1_24[161]}
   );
   gpc615_5 gpc930 (
      {stage0_24[236], stage0_24[237], stage0_24[238], stage0_24[239], stage0_24[240]},
      {stage0_25[68]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[21],stage1_26[49],stage1_25[115],stage1_24[162]}
   );
   gpc615_5 gpc931 (
      {stage0_24[241], stage0_24[242], stage0_24[243], stage0_24[244], stage0_24[245]},
      {stage0_25[69]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[22],stage1_26[50],stage1_25[116],stage1_24[163]}
   );
   gpc615_5 gpc932 (
      {stage0_24[246], stage0_24[247], stage0_24[248], stage0_24[249], stage0_24[250]},
      {stage0_25[70]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[23],stage1_26[51],stage1_25[117],stage1_24[164]}
   );
   gpc615_5 gpc933 (
      {stage0_24[251], stage0_24[252], stage0_24[253], stage0_24[254], stage0_24[255]},
      {stage0_25[71]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[24],stage1_26[52],stage1_25[118],stage1_24[165]}
   );
   gpc615_5 gpc934 (
      {stage0_24[256], stage0_24[257], stage0_24[258], stage0_24[259], stage0_24[260]},
      {stage0_25[72]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[25],stage1_26[53],stage1_25[119],stage1_24[166]}
   );
   gpc615_5 gpc935 (
      {stage0_24[261], stage0_24[262], stage0_24[263], stage0_24[264], stage0_24[265]},
      {stage0_25[73]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[26],stage1_26[54],stage1_25[120],stage1_24[167]}
   );
   gpc615_5 gpc936 (
      {stage0_24[266], stage0_24[267], stage0_24[268], stage0_24[269], stage0_24[270]},
      {stage0_25[74]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[27],stage1_26[55],stage1_25[121],stage1_24[168]}
   );
   gpc615_5 gpc937 (
      {stage0_24[271], stage0_24[272], stage0_24[273], stage0_24[274], stage0_24[275]},
      {stage0_25[75]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[28],stage1_26[56],stage1_25[122],stage1_24[169]}
   );
   gpc615_5 gpc938 (
      {stage0_24[276], stage0_24[277], stage0_24[278], stage0_24[279], stage0_24[280]},
      {stage0_25[76]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[29],stage1_26[57],stage1_25[123],stage1_24[170]}
   );
   gpc615_5 gpc939 (
      {stage0_24[281], stage0_24[282], stage0_24[283], stage0_24[284], stage0_24[285]},
      {stage0_25[77]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[30],stage1_26[58],stage1_25[124],stage1_24[171]}
   );
   gpc615_5 gpc940 (
      {stage0_24[286], stage0_24[287], stage0_24[288], stage0_24[289], stage0_24[290]},
      {stage0_25[78]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[31],stage1_26[59],stage1_25[125],stage1_24[172]}
   );
   gpc615_5 gpc941 (
      {stage0_24[291], stage0_24[292], stage0_24[293], stage0_24[294], stage0_24[295]},
      {stage0_25[79]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[32],stage1_26[60],stage1_25[126],stage1_24[173]}
   );
   gpc615_5 gpc942 (
      {stage0_24[296], stage0_24[297], stage0_24[298], stage0_24[299], stage0_24[300]},
      {stage0_25[80]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[33],stage1_26[61],stage1_25[127],stage1_24[174]}
   );
   gpc615_5 gpc943 (
      {stage0_24[301], stage0_24[302], stage0_24[303], stage0_24[304], stage0_24[305]},
      {stage0_25[81]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[34],stage1_26[62],stage1_25[128],stage1_24[175]}
   );
   gpc615_5 gpc944 (
      {stage0_24[306], stage0_24[307], stage0_24[308], stage0_24[309], stage0_24[310]},
      {stage0_25[82]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[35],stage1_26[63],stage1_25[129],stage1_24[176]}
   );
   gpc615_5 gpc945 (
      {stage0_24[311], stage0_24[312], stage0_24[313], stage0_24[314], stage0_24[315]},
      {stage0_25[83]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[36],stage1_26[64],stage1_25[130],stage1_24[177]}
   );
   gpc615_5 gpc946 (
      {stage0_24[316], stage0_24[317], stage0_24[318], stage0_24[319], stage0_24[320]},
      {stage0_25[84]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[37],stage1_26[65],stage1_25[131],stage1_24[178]}
   );
   gpc615_5 gpc947 (
      {stage0_24[321], stage0_24[322], stage0_24[323], stage0_24[324], stage0_24[325]},
      {stage0_25[85]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[38],stage1_26[66],stage1_25[132],stage1_24[179]}
   );
   gpc615_5 gpc948 (
      {stage0_24[326], stage0_24[327], stage0_24[328], stage0_24[329], stage0_24[330]},
      {stage0_25[86]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[39],stage1_26[67],stage1_25[133],stage1_24[180]}
   );
   gpc615_5 gpc949 (
      {stage0_24[331], stage0_24[332], stage0_24[333], stage0_24[334], stage0_24[335]},
      {stage0_25[87]},
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184], stage0_26[185]},
      {stage1_28[30],stage1_27[40],stage1_26[68],stage1_25[134],stage1_24[181]}
   );
   gpc615_5 gpc950 (
      {stage0_24[336], stage0_24[337], stage0_24[338], stage0_24[339], stage0_24[340]},
      {stage0_25[88]},
      {stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189], stage0_26[190], stage0_26[191]},
      {stage1_28[31],stage1_27[41],stage1_26[69],stage1_25[135],stage1_24[182]}
   );
   gpc615_5 gpc951 (
      {stage0_24[341], stage0_24[342], stage0_24[343], stage0_24[344], stage0_24[345]},
      {stage0_25[89]},
      {stage0_26[192], stage0_26[193], stage0_26[194], stage0_26[195], stage0_26[196], stage0_26[197]},
      {stage1_28[32],stage1_27[42],stage1_26[70],stage1_25[136],stage1_24[183]}
   );
   gpc615_5 gpc952 (
      {stage0_24[346], stage0_24[347], stage0_24[348], stage0_24[349], stage0_24[350]},
      {stage0_25[90]},
      {stage0_26[198], stage0_26[199], stage0_26[200], stage0_26[201], stage0_26[202], stage0_26[203]},
      {stage1_28[33],stage1_27[43],stage1_26[71],stage1_25[137],stage1_24[184]}
   );
   gpc615_5 gpc953 (
      {stage0_24[351], stage0_24[352], stage0_24[353], stage0_24[354], stage0_24[355]},
      {stage0_25[91]},
      {stage0_26[204], stage0_26[205], stage0_26[206], stage0_26[207], stage0_26[208], stage0_26[209]},
      {stage1_28[34],stage1_27[44],stage1_26[72],stage1_25[138],stage1_24[185]}
   );
   gpc615_5 gpc954 (
      {stage0_24[356], stage0_24[357], stage0_24[358], stage0_24[359], stage0_24[360]},
      {stage0_25[92]},
      {stage0_26[210], stage0_26[211], stage0_26[212], stage0_26[213], stage0_26[214], stage0_26[215]},
      {stage1_28[35],stage1_27[45],stage1_26[73],stage1_25[139],stage1_24[186]}
   );
   gpc615_5 gpc955 (
      {stage0_24[361], stage0_24[362], stage0_24[363], stage0_24[364], stage0_24[365]},
      {stage0_25[93]},
      {stage0_26[216], stage0_26[217], stage0_26[218], stage0_26[219], stage0_26[220], stage0_26[221]},
      {stage1_28[36],stage1_27[46],stage1_26[74],stage1_25[140],stage1_24[187]}
   );
   gpc615_5 gpc956 (
      {stage0_24[366], stage0_24[367], stage0_24[368], stage0_24[369], stage0_24[370]},
      {stage0_25[94]},
      {stage0_26[222], stage0_26[223], stage0_26[224], stage0_26[225], stage0_26[226], stage0_26[227]},
      {stage1_28[37],stage1_27[47],stage1_26[75],stage1_25[141],stage1_24[188]}
   );
   gpc615_5 gpc957 (
      {stage0_24[371], stage0_24[372], stage0_24[373], stage0_24[374], stage0_24[375]},
      {stage0_25[95]},
      {stage0_26[228], stage0_26[229], stage0_26[230], stage0_26[231], stage0_26[232], stage0_26[233]},
      {stage1_28[38],stage1_27[48],stage1_26[76],stage1_25[142],stage1_24[189]}
   );
   gpc615_5 gpc958 (
      {stage0_24[376], stage0_24[377], stage0_24[378], stage0_24[379], stage0_24[380]},
      {stage0_25[96]},
      {stage0_26[234], stage0_26[235], stage0_26[236], stage0_26[237], stage0_26[238], stage0_26[239]},
      {stage1_28[39],stage1_27[49],stage1_26[77],stage1_25[143],stage1_24[190]}
   );
   gpc615_5 gpc959 (
      {stage0_24[381], stage0_24[382], stage0_24[383], stage0_24[384], stage0_24[385]},
      {stage0_25[97]},
      {stage0_26[240], stage0_26[241], stage0_26[242], stage0_26[243], stage0_26[244], stage0_26[245]},
      {stage1_28[40],stage1_27[50],stage1_26[78],stage1_25[144],stage1_24[191]}
   );
   gpc615_5 gpc960 (
      {stage0_24[386], stage0_24[387], stage0_24[388], stage0_24[389], stage0_24[390]},
      {stage0_25[98]},
      {stage0_26[246], stage0_26[247], stage0_26[248], stage0_26[249], stage0_26[250], stage0_26[251]},
      {stage1_28[41],stage1_27[51],stage1_26[79],stage1_25[145],stage1_24[192]}
   );
   gpc615_5 gpc961 (
      {stage0_24[391], stage0_24[392], stage0_24[393], stage0_24[394], stage0_24[395]},
      {stage0_25[99]},
      {stage0_26[252], stage0_26[253], stage0_26[254], stage0_26[255], stage0_26[256], stage0_26[257]},
      {stage1_28[42],stage1_27[52],stage1_26[80],stage1_25[146],stage1_24[193]}
   );
   gpc615_5 gpc962 (
      {stage0_24[396], stage0_24[397], stage0_24[398], stage0_24[399], stage0_24[400]},
      {stage0_25[100]},
      {stage0_26[258], stage0_26[259], stage0_26[260], stage0_26[261], stage0_26[262], stage0_26[263]},
      {stage1_28[43],stage1_27[53],stage1_26[81],stage1_25[147],stage1_24[194]}
   );
   gpc615_5 gpc963 (
      {stage0_24[401], stage0_24[402], stage0_24[403], stage0_24[404], stage0_24[405]},
      {stage0_25[101]},
      {stage0_26[264], stage0_26[265], stage0_26[266], stage0_26[267], stage0_26[268], stage0_26[269]},
      {stage1_28[44],stage1_27[54],stage1_26[82],stage1_25[148],stage1_24[195]}
   );
   gpc615_5 gpc964 (
      {stage0_24[406], stage0_24[407], stage0_24[408], stage0_24[409], stage0_24[410]},
      {stage0_25[102]},
      {stage0_26[270], stage0_26[271], stage0_26[272], stage0_26[273], stage0_26[274], stage0_26[275]},
      {stage1_28[45],stage1_27[55],stage1_26[83],stage1_25[149],stage1_24[196]}
   );
   gpc615_5 gpc965 (
      {stage0_24[411], stage0_24[412], stage0_24[413], stage0_24[414], stage0_24[415]},
      {stage0_25[103]},
      {stage0_26[276], stage0_26[277], stage0_26[278], stage0_26[279], stage0_26[280], stage0_26[281]},
      {stage1_28[46],stage1_27[56],stage1_26[84],stage1_25[150],stage1_24[197]}
   );
   gpc615_5 gpc966 (
      {stage0_24[416], stage0_24[417], stage0_24[418], stage0_24[419], stage0_24[420]},
      {stage0_25[104]},
      {stage0_26[282], stage0_26[283], stage0_26[284], stage0_26[285], stage0_26[286], stage0_26[287]},
      {stage1_28[47],stage1_27[57],stage1_26[85],stage1_25[151],stage1_24[198]}
   );
   gpc615_5 gpc967 (
      {stage0_24[421], stage0_24[422], stage0_24[423], stage0_24[424], stage0_24[425]},
      {stage0_25[105]},
      {stage0_26[288], stage0_26[289], stage0_26[290], stage0_26[291], stage0_26[292], stage0_26[293]},
      {stage1_28[48],stage1_27[58],stage1_26[86],stage1_25[152],stage1_24[199]}
   );
   gpc615_5 gpc968 (
      {stage0_24[426], stage0_24[427], stage0_24[428], stage0_24[429], stage0_24[430]},
      {stage0_25[106]},
      {stage0_26[294], stage0_26[295], stage0_26[296], stage0_26[297], stage0_26[298], stage0_26[299]},
      {stage1_28[49],stage1_27[59],stage1_26[87],stage1_25[153],stage1_24[200]}
   );
   gpc615_5 gpc969 (
      {stage0_24[431], stage0_24[432], stage0_24[433], stage0_24[434], stage0_24[435]},
      {stage0_25[107]},
      {stage0_26[300], stage0_26[301], stage0_26[302], stage0_26[303], stage0_26[304], stage0_26[305]},
      {stage1_28[50],stage1_27[60],stage1_26[88],stage1_25[154],stage1_24[201]}
   );
   gpc615_5 gpc970 (
      {stage0_24[436], stage0_24[437], stage0_24[438], stage0_24[439], stage0_24[440]},
      {stage0_25[108]},
      {stage0_26[306], stage0_26[307], stage0_26[308], stage0_26[309], stage0_26[310], stage0_26[311]},
      {stage1_28[51],stage1_27[61],stage1_26[89],stage1_25[155],stage1_24[202]}
   );
   gpc615_5 gpc971 (
      {stage0_24[441], stage0_24[442], stage0_24[443], stage0_24[444], stage0_24[445]},
      {stage0_25[109]},
      {stage0_26[312], stage0_26[313], stage0_26[314], stage0_26[315], stage0_26[316], stage0_26[317]},
      {stage1_28[52],stage1_27[62],stage1_26[90],stage1_25[156],stage1_24[203]}
   );
   gpc615_5 gpc972 (
      {stage0_24[446], stage0_24[447], stage0_24[448], stage0_24[449], stage0_24[450]},
      {stage0_25[110]},
      {stage0_26[318], stage0_26[319], stage0_26[320], stage0_26[321], stage0_26[322], stage0_26[323]},
      {stage1_28[53],stage1_27[63],stage1_26[91],stage1_25[157],stage1_24[204]}
   );
   gpc615_5 gpc973 (
      {stage0_24[451], stage0_24[452], stage0_24[453], stage0_24[454], stage0_24[455]},
      {stage0_25[111]},
      {stage0_26[324], stage0_26[325], stage0_26[326], stage0_26[327], stage0_26[328], stage0_26[329]},
      {stage1_28[54],stage1_27[64],stage1_26[92],stage1_25[158],stage1_24[205]}
   );
   gpc615_5 gpc974 (
      {stage0_24[456], stage0_24[457], stage0_24[458], stage0_24[459], stage0_24[460]},
      {stage0_25[112]},
      {stage0_26[330], stage0_26[331], stage0_26[332], stage0_26[333], stage0_26[334], stage0_26[335]},
      {stage1_28[55],stage1_27[65],stage1_26[93],stage1_25[159],stage1_24[206]}
   );
   gpc615_5 gpc975 (
      {stage0_24[461], stage0_24[462], stage0_24[463], stage0_24[464], stage0_24[465]},
      {stage0_25[113]},
      {stage0_26[336], stage0_26[337], stage0_26[338], stage0_26[339], stage0_26[340], stage0_26[341]},
      {stage1_28[56],stage1_27[66],stage1_26[94],stage1_25[160],stage1_24[207]}
   );
   gpc615_5 gpc976 (
      {stage0_24[466], stage0_24[467], stage0_24[468], stage0_24[469], stage0_24[470]},
      {stage0_25[114]},
      {stage0_26[342], stage0_26[343], stage0_26[344], stage0_26[345], stage0_26[346], stage0_26[347]},
      {stage1_28[57],stage1_27[67],stage1_26[95],stage1_25[161],stage1_24[208]}
   );
   gpc615_5 gpc977 (
      {stage0_24[471], stage0_24[472], stage0_24[473], stage0_24[474], stage0_24[475]},
      {stage0_25[115]},
      {stage0_26[348], stage0_26[349], stage0_26[350], stage0_26[351], stage0_26[352], stage0_26[353]},
      {stage1_28[58],stage1_27[68],stage1_26[96],stage1_25[162],stage1_24[209]}
   );
   gpc615_5 gpc978 (
      {stage0_24[476], stage0_24[477], stage0_24[478], stage0_24[479], stage0_24[480]},
      {stage0_25[116]},
      {stage0_26[354], stage0_26[355], stage0_26[356], stage0_26[357], stage0_26[358], stage0_26[359]},
      {stage1_28[59],stage1_27[69],stage1_26[97],stage1_25[163],stage1_24[210]}
   );
   gpc615_5 gpc979 (
      {stage0_24[481], stage0_24[482], stage0_24[483], stage0_24[484], stage0_24[485]},
      {stage0_25[117]},
      {stage0_26[360], stage0_26[361], stage0_26[362], stage0_26[363], stage0_26[364], stage0_26[365]},
      {stage1_28[60],stage1_27[70],stage1_26[98],stage1_25[164],stage1_24[211]}
   );
   gpc606_5 gpc980 (
      {stage0_25[118], stage0_25[119], stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[61],stage1_27[71],stage1_26[99],stage1_25[165]}
   );
   gpc606_5 gpc981 (
      {stage0_25[124], stage0_25[125], stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[62],stage1_27[72],stage1_26[100],stage1_25[166]}
   );
   gpc606_5 gpc982 (
      {stage0_25[130], stage0_25[131], stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[63],stage1_27[73],stage1_26[101],stage1_25[167]}
   );
   gpc606_5 gpc983 (
      {stage0_25[136], stage0_25[137], stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[64],stage1_27[74],stage1_26[102],stage1_25[168]}
   );
   gpc606_5 gpc984 (
      {stage0_25[142], stage0_25[143], stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[65],stage1_27[75],stage1_26[103],stage1_25[169]}
   );
   gpc606_5 gpc985 (
      {stage0_25[148], stage0_25[149], stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[66],stage1_27[76],stage1_26[104],stage1_25[170]}
   );
   gpc606_5 gpc986 (
      {stage0_25[154], stage0_25[155], stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[67],stage1_27[77],stage1_26[105],stage1_25[171]}
   );
   gpc606_5 gpc987 (
      {stage0_25[160], stage0_25[161], stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[68],stage1_27[78],stage1_26[106],stage1_25[172]}
   );
   gpc606_5 gpc988 (
      {stage0_25[166], stage0_25[167], stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[69],stage1_27[79],stage1_26[107],stage1_25[173]}
   );
   gpc606_5 gpc989 (
      {stage0_25[172], stage0_25[173], stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[70],stage1_27[80],stage1_26[108],stage1_25[174]}
   );
   gpc606_5 gpc990 (
      {stage0_25[178], stage0_25[179], stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[71],stage1_27[81],stage1_26[109],stage1_25[175]}
   );
   gpc606_5 gpc991 (
      {stage0_25[184], stage0_25[185], stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[72],stage1_27[82],stage1_26[110],stage1_25[176]}
   );
   gpc606_5 gpc992 (
      {stage0_25[190], stage0_25[191], stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[73],stage1_27[83],stage1_26[111],stage1_25[177]}
   );
   gpc606_5 gpc993 (
      {stage0_25[196], stage0_25[197], stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[74],stage1_27[84],stage1_26[112],stage1_25[178]}
   );
   gpc606_5 gpc994 (
      {stage0_25[202], stage0_25[203], stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[75],stage1_27[85],stage1_26[113],stage1_25[179]}
   );
   gpc606_5 gpc995 (
      {stage0_25[208], stage0_25[209], stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[76],stage1_27[86],stage1_26[114],stage1_25[180]}
   );
   gpc606_5 gpc996 (
      {stage0_25[214], stage0_25[215], stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[77],stage1_27[87],stage1_26[115],stage1_25[181]}
   );
   gpc606_5 gpc997 (
      {stage0_25[220], stage0_25[221], stage0_25[222], stage0_25[223], stage0_25[224], stage0_25[225]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[78],stage1_27[88],stage1_26[116],stage1_25[182]}
   );
   gpc615_5 gpc998 (
      {stage0_25[226], stage0_25[227], stage0_25[228], stage0_25[229], stage0_25[230]},
      {stage0_26[366]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[79],stage1_27[89],stage1_26[117],stage1_25[183]}
   );
   gpc615_5 gpc999 (
      {stage0_25[231], stage0_25[232], stage0_25[233], stage0_25[234], stage0_25[235]},
      {stage0_26[367]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[80],stage1_27[90],stage1_26[118],stage1_25[184]}
   );
   gpc615_5 gpc1000 (
      {stage0_25[236], stage0_25[237], stage0_25[238], stage0_25[239], stage0_25[240]},
      {stage0_26[368]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[81],stage1_27[91],stage1_26[119],stage1_25[185]}
   );
   gpc615_5 gpc1001 (
      {stage0_25[241], stage0_25[242], stage0_25[243], stage0_25[244], stage0_25[245]},
      {stage0_26[369]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[82],stage1_27[92],stage1_26[120],stage1_25[186]}
   );
   gpc615_5 gpc1002 (
      {stage0_25[246], stage0_25[247], stage0_25[248], stage0_25[249], stage0_25[250]},
      {stage0_26[370]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[83],stage1_27[93],stage1_26[121],stage1_25[187]}
   );
   gpc615_5 gpc1003 (
      {stage0_25[251], stage0_25[252], stage0_25[253], stage0_25[254], stage0_25[255]},
      {stage0_26[371]},
      {stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141], stage0_27[142], stage0_27[143]},
      {stage1_29[23],stage1_28[84],stage1_27[94],stage1_26[122],stage1_25[188]}
   );
   gpc615_5 gpc1004 (
      {stage0_25[256], stage0_25[257], stage0_25[258], stage0_25[259], stage0_25[260]},
      {stage0_26[372]},
      {stage0_27[144], stage0_27[145], stage0_27[146], stage0_27[147], stage0_27[148], stage0_27[149]},
      {stage1_29[24],stage1_28[85],stage1_27[95],stage1_26[123],stage1_25[189]}
   );
   gpc615_5 gpc1005 (
      {stage0_25[261], stage0_25[262], stage0_25[263], stage0_25[264], stage0_25[265]},
      {stage0_26[373]},
      {stage0_27[150], stage0_27[151], stage0_27[152], stage0_27[153], stage0_27[154], stage0_27[155]},
      {stage1_29[25],stage1_28[86],stage1_27[96],stage1_26[124],stage1_25[190]}
   );
   gpc615_5 gpc1006 (
      {stage0_25[266], stage0_25[267], stage0_25[268], stage0_25[269], stage0_25[270]},
      {stage0_26[374]},
      {stage0_27[156], stage0_27[157], stage0_27[158], stage0_27[159], stage0_27[160], stage0_27[161]},
      {stage1_29[26],stage1_28[87],stage1_27[97],stage1_26[125],stage1_25[191]}
   );
   gpc615_5 gpc1007 (
      {stage0_25[271], stage0_25[272], stage0_25[273], stage0_25[274], stage0_25[275]},
      {stage0_26[375]},
      {stage0_27[162], stage0_27[163], stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167]},
      {stage1_29[27],stage1_28[88],stage1_27[98],stage1_26[126],stage1_25[192]}
   );
   gpc615_5 gpc1008 (
      {stage0_25[276], stage0_25[277], stage0_25[278], stage0_25[279], stage0_25[280]},
      {stage0_26[376]},
      {stage0_27[168], stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage1_29[28],stage1_28[89],stage1_27[99],stage1_26[127],stage1_25[193]}
   );
   gpc615_5 gpc1009 (
      {stage0_25[281], stage0_25[282], stage0_25[283], stage0_25[284], stage0_25[285]},
      {stage0_26[377]},
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178], stage0_27[179]},
      {stage1_29[29],stage1_28[90],stage1_27[100],stage1_26[128],stage1_25[194]}
   );
   gpc615_5 gpc1010 (
      {stage0_25[286], stage0_25[287], stage0_25[288], stage0_25[289], stage0_25[290]},
      {stage0_26[378]},
      {stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183], stage0_27[184], stage0_27[185]},
      {stage1_29[30],stage1_28[91],stage1_27[101],stage1_26[129],stage1_25[195]}
   );
   gpc615_5 gpc1011 (
      {stage0_25[291], stage0_25[292], stage0_25[293], stage0_25[294], stage0_25[295]},
      {stage0_26[379]},
      {stage0_27[186], stage0_27[187], stage0_27[188], stage0_27[189], stage0_27[190], stage0_27[191]},
      {stage1_29[31],stage1_28[92],stage1_27[102],stage1_26[130],stage1_25[196]}
   );
   gpc615_5 gpc1012 (
      {stage0_25[296], stage0_25[297], stage0_25[298], stage0_25[299], stage0_25[300]},
      {stage0_26[380]},
      {stage0_27[192], stage0_27[193], stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197]},
      {stage1_29[32],stage1_28[93],stage1_27[103],stage1_26[131],stage1_25[197]}
   );
   gpc615_5 gpc1013 (
      {stage0_25[301], stage0_25[302], stage0_25[303], stage0_25[304], stage0_25[305]},
      {stage0_26[381]},
      {stage0_27[198], stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage1_29[33],stage1_28[94],stage1_27[104],stage1_26[132],stage1_25[198]}
   );
   gpc615_5 gpc1014 (
      {stage0_25[306], stage0_25[307], stage0_25[308], stage0_25[309], stage0_25[310]},
      {stage0_26[382]},
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208], stage0_27[209]},
      {stage1_29[34],stage1_28[95],stage1_27[105],stage1_26[133],stage1_25[199]}
   );
   gpc615_5 gpc1015 (
      {stage0_25[311], stage0_25[312], stage0_25[313], stage0_25[314], stage0_25[315]},
      {stage0_26[383]},
      {stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213], stage0_27[214], stage0_27[215]},
      {stage1_29[35],stage1_28[96],stage1_27[106],stage1_26[134],stage1_25[200]}
   );
   gpc615_5 gpc1016 (
      {stage0_25[316], stage0_25[317], stage0_25[318], stage0_25[319], stage0_25[320]},
      {stage0_26[384]},
      {stage0_27[216], stage0_27[217], stage0_27[218], stage0_27[219], stage0_27[220], stage0_27[221]},
      {stage1_29[36],stage1_28[97],stage1_27[107],stage1_26[135],stage1_25[201]}
   );
   gpc615_5 gpc1017 (
      {stage0_25[321], stage0_25[322], stage0_25[323], stage0_25[324], stage0_25[325]},
      {stage0_26[385]},
      {stage0_27[222], stage0_27[223], stage0_27[224], stage0_27[225], stage0_27[226], stage0_27[227]},
      {stage1_29[37],stage1_28[98],stage1_27[108],stage1_26[136],stage1_25[202]}
   );
   gpc615_5 gpc1018 (
      {stage0_25[326], stage0_25[327], stage0_25[328], stage0_25[329], stage0_25[330]},
      {stage0_26[386]},
      {stage0_27[228], stage0_27[229], stage0_27[230], stage0_27[231], stage0_27[232], stage0_27[233]},
      {stage1_29[38],stage1_28[99],stage1_27[109],stage1_26[137],stage1_25[203]}
   );
   gpc615_5 gpc1019 (
      {stage0_25[331], stage0_25[332], stage0_25[333], stage0_25[334], stage0_25[335]},
      {stage0_26[387]},
      {stage0_27[234], stage0_27[235], stage0_27[236], stage0_27[237], stage0_27[238], stage0_27[239]},
      {stage1_29[39],stage1_28[100],stage1_27[110],stage1_26[138],stage1_25[204]}
   );
   gpc615_5 gpc1020 (
      {stage0_25[336], stage0_25[337], stage0_25[338], stage0_25[339], stage0_25[340]},
      {stage0_26[388]},
      {stage0_27[240], stage0_27[241], stage0_27[242], stage0_27[243], stage0_27[244], stage0_27[245]},
      {stage1_29[40],stage1_28[101],stage1_27[111],stage1_26[139],stage1_25[205]}
   );
   gpc615_5 gpc1021 (
      {stage0_25[341], stage0_25[342], stage0_25[343], stage0_25[344], stage0_25[345]},
      {stage0_26[389]},
      {stage0_27[246], stage0_27[247], stage0_27[248], stage0_27[249], stage0_27[250], stage0_27[251]},
      {stage1_29[41],stage1_28[102],stage1_27[112],stage1_26[140],stage1_25[206]}
   );
   gpc615_5 gpc1022 (
      {stage0_25[346], stage0_25[347], stage0_25[348], stage0_25[349], stage0_25[350]},
      {stage0_26[390]},
      {stage0_27[252], stage0_27[253], stage0_27[254], stage0_27[255], stage0_27[256], stage0_27[257]},
      {stage1_29[42],stage1_28[103],stage1_27[113],stage1_26[141],stage1_25[207]}
   );
   gpc615_5 gpc1023 (
      {stage0_25[351], stage0_25[352], stage0_25[353], stage0_25[354], stage0_25[355]},
      {stage0_26[391]},
      {stage0_27[258], stage0_27[259], stage0_27[260], stage0_27[261], stage0_27[262], stage0_27[263]},
      {stage1_29[43],stage1_28[104],stage1_27[114],stage1_26[142],stage1_25[208]}
   );
   gpc615_5 gpc1024 (
      {stage0_25[356], stage0_25[357], stage0_25[358], stage0_25[359], stage0_25[360]},
      {stage0_26[392]},
      {stage0_27[264], stage0_27[265], stage0_27[266], stage0_27[267], stage0_27[268], stage0_27[269]},
      {stage1_29[44],stage1_28[105],stage1_27[115],stage1_26[143],stage1_25[209]}
   );
   gpc615_5 gpc1025 (
      {stage0_25[361], stage0_25[362], stage0_25[363], stage0_25[364], stage0_25[365]},
      {stage0_26[393]},
      {stage0_27[270], stage0_27[271], stage0_27[272], stage0_27[273], stage0_27[274], stage0_27[275]},
      {stage1_29[45],stage1_28[106],stage1_27[116],stage1_26[144],stage1_25[210]}
   );
   gpc615_5 gpc1026 (
      {stage0_25[366], stage0_25[367], stage0_25[368], stage0_25[369], stage0_25[370]},
      {stage0_26[394]},
      {stage0_27[276], stage0_27[277], stage0_27[278], stage0_27[279], stage0_27[280], stage0_27[281]},
      {stage1_29[46],stage1_28[107],stage1_27[117],stage1_26[145],stage1_25[211]}
   );
   gpc615_5 gpc1027 (
      {stage0_25[371], stage0_25[372], stage0_25[373], stage0_25[374], stage0_25[375]},
      {stage0_26[395]},
      {stage0_27[282], stage0_27[283], stage0_27[284], stage0_27[285], stage0_27[286], stage0_27[287]},
      {stage1_29[47],stage1_28[108],stage1_27[118],stage1_26[146],stage1_25[212]}
   );
   gpc615_5 gpc1028 (
      {stage0_25[376], stage0_25[377], stage0_25[378], stage0_25[379], stage0_25[380]},
      {stage0_26[396]},
      {stage0_27[288], stage0_27[289], stage0_27[290], stage0_27[291], stage0_27[292], stage0_27[293]},
      {stage1_29[48],stage1_28[109],stage1_27[119],stage1_26[147],stage1_25[213]}
   );
   gpc615_5 gpc1029 (
      {stage0_25[381], stage0_25[382], stage0_25[383], stage0_25[384], stage0_25[385]},
      {stage0_26[397]},
      {stage0_27[294], stage0_27[295], stage0_27[296], stage0_27[297], stage0_27[298], stage0_27[299]},
      {stage1_29[49],stage1_28[110],stage1_27[120],stage1_26[148],stage1_25[214]}
   );
   gpc615_5 gpc1030 (
      {stage0_25[386], stage0_25[387], stage0_25[388], stage0_25[389], stage0_25[390]},
      {stage0_26[398]},
      {stage0_27[300], stage0_27[301], stage0_27[302], stage0_27[303], stage0_27[304], stage0_27[305]},
      {stage1_29[50],stage1_28[111],stage1_27[121],stage1_26[149],stage1_25[215]}
   );
   gpc615_5 gpc1031 (
      {stage0_25[391], stage0_25[392], stage0_25[393], stage0_25[394], stage0_25[395]},
      {stage0_26[399]},
      {stage0_27[306], stage0_27[307], stage0_27[308], stage0_27[309], stage0_27[310], stage0_27[311]},
      {stage1_29[51],stage1_28[112],stage1_27[122],stage1_26[150],stage1_25[216]}
   );
   gpc615_5 gpc1032 (
      {stage0_25[396], stage0_25[397], stage0_25[398], stage0_25[399], stage0_25[400]},
      {stage0_26[400]},
      {stage0_27[312], stage0_27[313], stage0_27[314], stage0_27[315], stage0_27[316], stage0_27[317]},
      {stage1_29[52],stage1_28[113],stage1_27[123],stage1_26[151],stage1_25[217]}
   );
   gpc615_5 gpc1033 (
      {stage0_25[401], stage0_25[402], stage0_25[403], stage0_25[404], stage0_25[405]},
      {stage0_26[401]},
      {stage0_27[318], stage0_27[319], stage0_27[320], stage0_27[321], stage0_27[322], stage0_27[323]},
      {stage1_29[53],stage1_28[114],stage1_27[124],stage1_26[152],stage1_25[218]}
   );
   gpc615_5 gpc1034 (
      {stage0_25[406], stage0_25[407], stage0_25[408], stage0_25[409], stage0_25[410]},
      {stage0_26[402]},
      {stage0_27[324], stage0_27[325], stage0_27[326], stage0_27[327], stage0_27[328], stage0_27[329]},
      {stage1_29[54],stage1_28[115],stage1_27[125],stage1_26[153],stage1_25[219]}
   );
   gpc615_5 gpc1035 (
      {stage0_25[411], stage0_25[412], stage0_25[413], stage0_25[414], stage0_25[415]},
      {stage0_26[403]},
      {stage0_27[330], stage0_27[331], stage0_27[332], stage0_27[333], stage0_27[334], stage0_27[335]},
      {stage1_29[55],stage1_28[116],stage1_27[126],stage1_26[154],stage1_25[220]}
   );
   gpc615_5 gpc1036 (
      {stage0_25[416], stage0_25[417], stage0_25[418], stage0_25[419], stage0_25[420]},
      {stage0_26[404]},
      {stage0_27[336], stage0_27[337], stage0_27[338], stage0_27[339], stage0_27[340], stage0_27[341]},
      {stage1_29[56],stage1_28[117],stage1_27[127],stage1_26[155],stage1_25[221]}
   );
   gpc615_5 gpc1037 (
      {stage0_25[421], stage0_25[422], stage0_25[423], stage0_25[424], stage0_25[425]},
      {stage0_26[405]},
      {stage0_27[342], stage0_27[343], stage0_27[344], stage0_27[345], stage0_27[346], stage0_27[347]},
      {stage1_29[57],stage1_28[118],stage1_27[128],stage1_26[156],stage1_25[222]}
   );
   gpc615_5 gpc1038 (
      {stage0_25[426], stage0_25[427], stage0_25[428], stage0_25[429], stage0_25[430]},
      {stage0_26[406]},
      {stage0_27[348], stage0_27[349], stage0_27[350], stage0_27[351], stage0_27[352], stage0_27[353]},
      {stage1_29[58],stage1_28[119],stage1_27[129],stage1_26[157],stage1_25[223]}
   );
   gpc615_5 gpc1039 (
      {stage0_25[431], stage0_25[432], stage0_25[433], stage0_25[434], stage0_25[435]},
      {stage0_26[407]},
      {stage0_27[354], stage0_27[355], stage0_27[356], stage0_27[357], stage0_27[358], stage0_27[359]},
      {stage1_29[59],stage1_28[120],stage1_27[130],stage1_26[158],stage1_25[224]}
   );
   gpc615_5 gpc1040 (
      {stage0_25[436], stage0_25[437], stage0_25[438], stage0_25[439], stage0_25[440]},
      {stage0_26[408]},
      {stage0_27[360], stage0_27[361], stage0_27[362], stage0_27[363], stage0_27[364], stage0_27[365]},
      {stage1_29[60],stage1_28[121],stage1_27[131],stage1_26[159],stage1_25[225]}
   );
   gpc615_5 gpc1041 (
      {stage0_25[441], stage0_25[442], stage0_25[443], stage0_25[444], stage0_25[445]},
      {stage0_26[409]},
      {stage0_27[366], stage0_27[367], stage0_27[368], stage0_27[369], stage0_27[370], stage0_27[371]},
      {stage1_29[61],stage1_28[122],stage1_27[132],stage1_26[160],stage1_25[226]}
   );
   gpc615_5 gpc1042 (
      {stage0_25[446], stage0_25[447], stage0_25[448], stage0_25[449], stage0_25[450]},
      {stage0_26[410]},
      {stage0_27[372], stage0_27[373], stage0_27[374], stage0_27[375], stage0_27[376], stage0_27[377]},
      {stage1_29[62],stage1_28[123],stage1_27[133],stage1_26[161],stage1_25[227]}
   );
   gpc615_5 gpc1043 (
      {stage0_25[451], stage0_25[452], stage0_25[453], stage0_25[454], stage0_25[455]},
      {stage0_26[411]},
      {stage0_27[378], stage0_27[379], stage0_27[380], stage0_27[381], stage0_27[382], stage0_27[383]},
      {stage1_29[63],stage1_28[124],stage1_27[134],stage1_26[162],stage1_25[228]}
   );
   gpc615_5 gpc1044 (
      {stage0_25[456], stage0_25[457], stage0_25[458], stage0_25[459], stage0_25[460]},
      {stage0_26[412]},
      {stage0_27[384], stage0_27[385], stage0_27[386], stage0_27[387], stage0_27[388], stage0_27[389]},
      {stage1_29[64],stage1_28[125],stage1_27[135],stage1_26[163],stage1_25[229]}
   );
   gpc615_5 gpc1045 (
      {stage0_25[461], stage0_25[462], stage0_25[463], stage0_25[464], stage0_25[465]},
      {stage0_26[413]},
      {stage0_27[390], stage0_27[391], stage0_27[392], stage0_27[393], stage0_27[394], stage0_27[395]},
      {stage1_29[65],stage1_28[126],stage1_27[136],stage1_26[164],stage1_25[230]}
   );
   gpc615_5 gpc1046 (
      {stage0_25[466], stage0_25[467], stage0_25[468], stage0_25[469], stage0_25[470]},
      {stage0_26[414]},
      {stage0_27[396], stage0_27[397], stage0_27[398], stage0_27[399], stage0_27[400], stage0_27[401]},
      {stage1_29[66],stage1_28[127],stage1_27[137],stage1_26[165],stage1_25[231]}
   );
   gpc615_5 gpc1047 (
      {stage0_25[471], stage0_25[472], stage0_25[473], stage0_25[474], stage0_25[475]},
      {stage0_26[415]},
      {stage0_27[402], stage0_27[403], stage0_27[404], stage0_27[405], stage0_27[406], stage0_27[407]},
      {stage1_29[67],stage1_28[128],stage1_27[138],stage1_26[166],stage1_25[232]}
   );
   gpc615_5 gpc1048 (
      {stage0_25[476], stage0_25[477], stage0_25[478], stage0_25[479], stage0_25[480]},
      {stage0_26[416]},
      {stage0_27[408], stage0_27[409], stage0_27[410], stage0_27[411], stage0_27[412], stage0_27[413]},
      {stage1_29[68],stage1_28[129],stage1_27[139],stage1_26[167],stage1_25[233]}
   );
   gpc615_5 gpc1049 (
      {stage0_25[481], stage0_25[482], stage0_25[483], stage0_25[484], stage0_25[485]},
      {stage0_26[417]},
      {stage0_27[414], stage0_27[415], stage0_27[416], stage0_27[417], stage0_27[418], stage0_27[419]},
      {stage1_29[69],stage1_28[130],stage1_27[140],stage1_26[168],stage1_25[234]}
   );
   gpc606_5 gpc1050 (
      {stage0_26[418], stage0_26[419], stage0_26[420], stage0_26[421], stage0_26[422], stage0_26[423]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[70],stage1_28[131],stage1_27[141],stage1_26[169]}
   );
   gpc606_5 gpc1051 (
      {stage0_26[424], stage0_26[425], stage0_26[426], stage0_26[427], stage0_26[428], stage0_26[429]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[71],stage1_28[132],stage1_27[142],stage1_26[170]}
   );
   gpc615_5 gpc1052 (
      {stage0_26[430], stage0_26[431], stage0_26[432], stage0_26[433], stage0_26[434]},
      {stage0_27[420]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[72],stage1_28[133],stage1_27[143],stage1_26[171]}
   );
   gpc615_5 gpc1053 (
      {stage0_26[435], stage0_26[436], stage0_26[437], stage0_26[438], stage0_26[439]},
      {stage0_27[421]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[73],stage1_28[134],stage1_27[144],stage1_26[172]}
   );
   gpc615_5 gpc1054 (
      {stage0_26[440], stage0_26[441], stage0_26[442], stage0_26[443], stage0_26[444]},
      {stage0_27[422]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[74],stage1_28[135],stage1_27[145],stage1_26[173]}
   );
   gpc606_5 gpc1055 (
      {stage0_27[423], stage0_27[424], stage0_27[425], stage0_27[426], stage0_27[427], stage0_27[428]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[5],stage1_29[75],stage1_28[136],stage1_27[146]}
   );
   gpc606_5 gpc1056 (
      {stage0_27[429], stage0_27[430], stage0_27[431], stage0_27[432], stage0_27[433], stage0_27[434]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[6],stage1_29[76],stage1_28[137],stage1_27[147]}
   );
   gpc606_5 gpc1057 (
      {stage0_27[435], stage0_27[436], stage0_27[437], stage0_27[438], stage0_27[439], stage0_27[440]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[7],stage1_29[77],stage1_28[138],stage1_27[148]}
   );
   gpc606_5 gpc1058 (
      {stage0_27[441], stage0_27[442], stage0_27[443], stage0_27[444], stage0_27[445], stage0_27[446]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[8],stage1_29[78],stage1_28[139],stage1_27[149]}
   );
   gpc606_5 gpc1059 (
      {stage0_27[447], stage0_27[448], stage0_27[449], stage0_27[450], stage0_27[451], stage0_27[452]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[9],stage1_29[79],stage1_28[140],stage1_27[150]}
   );
   gpc606_5 gpc1060 (
      {stage0_27[453], stage0_27[454], stage0_27[455], stage0_27[456], stage0_27[457], stage0_27[458]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[10],stage1_29[80],stage1_28[141],stage1_27[151]}
   );
   gpc606_5 gpc1061 (
      {stage0_27[459], stage0_27[460], stage0_27[461], stage0_27[462], stage0_27[463], stage0_27[464]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[11],stage1_29[81],stage1_28[142],stage1_27[152]}
   );
   gpc606_5 gpc1062 (
      {stage0_27[465], stage0_27[466], stage0_27[467], stage0_27[468], stage0_27[469], stage0_27[470]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[12],stage1_29[82],stage1_28[143],stage1_27[153]}
   );
   gpc606_5 gpc1063 (
      {stage0_27[471], stage0_27[472], stage0_27[473], stage0_27[474], stage0_27[475], stage0_27[476]},
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage1_31[8],stage1_30[13],stage1_29[83],stage1_28[144],stage1_27[154]}
   );
   gpc606_5 gpc1064 (
      {stage0_27[477], stage0_27[478], stage0_27[479], stage0_27[480], stage0_27[481], stage0_27[482]},
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage1_31[9],stage1_30[14],stage1_29[84],stage1_28[145],stage1_27[155]}
   );
   gpc606_5 gpc1065 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[10],stage1_30[15],stage1_29[85],stage1_28[146]}
   );
   gpc606_5 gpc1066 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[11],stage1_30[16],stage1_29[86],stage1_28[147]}
   );
   gpc606_5 gpc1067 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[12],stage1_30[17],stage1_29[87],stage1_28[148]}
   );
   gpc606_5 gpc1068 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[13],stage1_30[18],stage1_29[88],stage1_28[149]}
   );
   gpc606_5 gpc1069 (
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[14],stage1_30[19],stage1_29[89],stage1_28[150]}
   );
   gpc606_5 gpc1070 (
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[15],stage1_30[20],stage1_29[90],stage1_28[151]}
   );
   gpc606_5 gpc1071 (
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[16],stage1_30[21],stage1_29[91],stage1_28[152]}
   );
   gpc606_5 gpc1072 (
      {stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[17],stage1_30[22],stage1_29[92],stage1_28[153]}
   );
   gpc606_5 gpc1073 (
      {stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[18],stage1_30[23],stage1_29[93],stage1_28[154]}
   );
   gpc606_5 gpc1074 (
      {stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[19],stage1_30[24],stage1_29[94],stage1_28[155]}
   );
   gpc606_5 gpc1075 (
      {stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[20],stage1_30[25],stage1_29[95],stage1_28[156]}
   );
   gpc606_5 gpc1076 (
      {stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[21],stage1_30[26],stage1_29[96],stage1_28[157]}
   );
   gpc606_5 gpc1077 (
      {stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[22],stage1_30[27],stage1_29[97],stage1_28[158]}
   );
   gpc606_5 gpc1078 (
      {stage0_28[108], stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[23],stage1_30[28],stage1_29[98],stage1_28[159]}
   );
   gpc606_5 gpc1079 (
      {stage0_28[114], stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[24],stage1_30[29],stage1_29[99],stage1_28[160]}
   );
   gpc606_5 gpc1080 (
      {stage0_28[120], stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[25],stage1_30[30],stage1_29[100],stage1_28[161]}
   );
   gpc606_5 gpc1081 (
      {stage0_28[126], stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[26],stage1_30[31],stage1_29[101],stage1_28[162]}
   );
   gpc606_5 gpc1082 (
      {stage0_28[132], stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[27],stage1_30[32],stage1_29[102],stage1_28[163]}
   );
   gpc606_5 gpc1083 (
      {stage0_28[138], stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143]},
      {stage0_30[108], stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113]},
      {stage1_32[18],stage1_31[28],stage1_30[33],stage1_29[103],stage1_28[164]}
   );
   gpc606_5 gpc1084 (
      {stage0_28[144], stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149]},
      {stage0_30[114], stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119]},
      {stage1_32[19],stage1_31[29],stage1_30[34],stage1_29[104],stage1_28[165]}
   );
   gpc606_5 gpc1085 (
      {stage0_28[150], stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155]},
      {stage0_30[120], stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125]},
      {stage1_32[20],stage1_31[30],stage1_30[35],stage1_29[105],stage1_28[166]}
   );
   gpc606_5 gpc1086 (
      {stage0_28[156], stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161]},
      {stage0_30[126], stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131]},
      {stage1_32[21],stage1_31[31],stage1_30[36],stage1_29[106],stage1_28[167]}
   );
   gpc606_5 gpc1087 (
      {stage0_28[162], stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167]},
      {stage0_30[132], stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137]},
      {stage1_32[22],stage1_31[32],stage1_30[37],stage1_29[107],stage1_28[168]}
   );
   gpc606_5 gpc1088 (
      {stage0_28[168], stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173]},
      {stage0_30[138], stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143]},
      {stage1_32[23],stage1_31[33],stage1_30[38],stage1_29[108],stage1_28[169]}
   );
   gpc606_5 gpc1089 (
      {stage0_28[174], stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179]},
      {stage0_30[144], stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149]},
      {stage1_32[24],stage1_31[34],stage1_30[39],stage1_29[109],stage1_28[170]}
   );
   gpc606_5 gpc1090 (
      {stage0_28[180], stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185]},
      {stage0_30[150], stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155]},
      {stage1_32[25],stage1_31[35],stage1_30[40],stage1_29[110],stage1_28[171]}
   );
   gpc606_5 gpc1091 (
      {stage0_28[186], stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191]},
      {stage0_30[156], stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161]},
      {stage1_32[26],stage1_31[36],stage1_30[41],stage1_29[111],stage1_28[172]}
   );
   gpc606_5 gpc1092 (
      {stage0_28[192], stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197]},
      {stage0_30[162], stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167]},
      {stage1_32[27],stage1_31[37],stage1_30[42],stage1_29[112],stage1_28[173]}
   );
   gpc606_5 gpc1093 (
      {stage0_28[198], stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203]},
      {stage0_30[168], stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173]},
      {stage1_32[28],stage1_31[38],stage1_30[43],stage1_29[113],stage1_28[174]}
   );
   gpc606_5 gpc1094 (
      {stage0_28[204], stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209]},
      {stage0_30[174], stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179]},
      {stage1_32[29],stage1_31[39],stage1_30[44],stage1_29[114],stage1_28[175]}
   );
   gpc606_5 gpc1095 (
      {stage0_28[210], stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215]},
      {stage0_30[180], stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185]},
      {stage1_32[30],stage1_31[40],stage1_30[45],stage1_29[115],stage1_28[176]}
   );
   gpc606_5 gpc1096 (
      {stage0_28[216], stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221]},
      {stage0_30[186], stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191]},
      {stage1_32[31],stage1_31[41],stage1_30[46],stage1_29[116],stage1_28[177]}
   );
   gpc606_5 gpc1097 (
      {stage0_28[222], stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227]},
      {stage0_30[192], stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197]},
      {stage1_32[32],stage1_31[42],stage1_30[47],stage1_29[117],stage1_28[178]}
   );
   gpc606_5 gpc1098 (
      {stage0_28[228], stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233]},
      {stage0_30[198], stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage1_32[33],stage1_31[43],stage1_30[48],stage1_29[118],stage1_28[179]}
   );
   gpc606_5 gpc1099 (
      {stage0_28[234], stage0_28[235], stage0_28[236], stage0_28[237], stage0_28[238], stage0_28[239]},
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208], stage0_30[209]},
      {stage1_32[34],stage1_31[44],stage1_30[49],stage1_29[119],stage1_28[180]}
   );
   gpc606_5 gpc1100 (
      {stage0_28[240], stage0_28[241], stage0_28[242], stage0_28[243], stage0_28[244], stage0_28[245]},
      {stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213], stage0_30[214], stage0_30[215]},
      {stage1_32[35],stage1_31[45],stage1_30[50],stage1_29[120],stage1_28[181]}
   );
   gpc606_5 gpc1101 (
      {stage0_28[246], stage0_28[247], stage0_28[248], stage0_28[249], stage0_28[250], stage0_28[251]},
      {stage0_30[216], stage0_30[217], stage0_30[218], stage0_30[219], stage0_30[220], stage0_30[221]},
      {stage1_32[36],stage1_31[46],stage1_30[51],stage1_29[121],stage1_28[182]}
   );
   gpc606_5 gpc1102 (
      {stage0_28[252], stage0_28[253], stage0_28[254], stage0_28[255], stage0_28[256], stage0_28[257]},
      {stage0_30[222], stage0_30[223], stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227]},
      {stage1_32[37],stage1_31[47],stage1_30[52],stage1_29[122],stage1_28[183]}
   );
   gpc606_5 gpc1103 (
      {stage0_28[258], stage0_28[259], stage0_28[260], stage0_28[261], stage0_28[262], stage0_28[263]},
      {stage0_30[228], stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage1_32[38],stage1_31[48],stage1_30[53],stage1_29[123],stage1_28[184]}
   );
   gpc606_5 gpc1104 (
      {stage0_28[264], stage0_28[265], stage0_28[266], stage0_28[267], stage0_28[268], stage0_28[269]},
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238], stage0_30[239]},
      {stage1_32[39],stage1_31[49],stage1_30[54],stage1_29[124],stage1_28[185]}
   );
   gpc606_5 gpc1105 (
      {stage0_28[270], stage0_28[271], stage0_28[272], stage0_28[273], stage0_28[274], stage0_28[275]},
      {stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243], stage0_30[244], stage0_30[245]},
      {stage1_32[40],stage1_31[50],stage1_30[55],stage1_29[125],stage1_28[186]}
   );
   gpc606_5 gpc1106 (
      {stage0_28[276], stage0_28[277], stage0_28[278], stage0_28[279], stage0_28[280], stage0_28[281]},
      {stage0_30[246], stage0_30[247], stage0_30[248], stage0_30[249], stage0_30[250], stage0_30[251]},
      {stage1_32[41],stage1_31[51],stage1_30[56],stage1_29[126],stage1_28[187]}
   );
   gpc606_5 gpc1107 (
      {stage0_28[282], stage0_28[283], stage0_28[284], stage0_28[285], stage0_28[286], stage0_28[287]},
      {stage0_30[252], stage0_30[253], stage0_30[254], stage0_30[255], stage0_30[256], stage0_30[257]},
      {stage1_32[42],stage1_31[52],stage1_30[57],stage1_29[127],stage1_28[188]}
   );
   gpc606_5 gpc1108 (
      {stage0_28[288], stage0_28[289], stage0_28[290], stage0_28[291], stage0_28[292], stage0_28[293]},
      {stage0_30[258], stage0_30[259], stage0_30[260], stage0_30[261], stage0_30[262], stage0_30[263]},
      {stage1_32[43],stage1_31[53],stage1_30[58],stage1_29[128],stage1_28[189]}
   );
   gpc606_5 gpc1109 (
      {stage0_28[294], stage0_28[295], stage0_28[296], stage0_28[297], stage0_28[298], stage0_28[299]},
      {stage0_30[264], stage0_30[265], stage0_30[266], stage0_30[267], stage0_30[268], stage0_30[269]},
      {stage1_32[44],stage1_31[54],stage1_30[59],stage1_29[129],stage1_28[190]}
   );
   gpc606_5 gpc1110 (
      {stage0_28[300], stage0_28[301], stage0_28[302], stage0_28[303], stage0_28[304], stage0_28[305]},
      {stage0_30[270], stage0_30[271], stage0_30[272], stage0_30[273], stage0_30[274], stage0_30[275]},
      {stage1_32[45],stage1_31[55],stage1_30[60],stage1_29[130],stage1_28[191]}
   );
   gpc606_5 gpc1111 (
      {stage0_28[306], stage0_28[307], stage0_28[308], stage0_28[309], stage0_28[310], stage0_28[311]},
      {stage0_30[276], stage0_30[277], stage0_30[278], stage0_30[279], stage0_30[280], stage0_30[281]},
      {stage1_32[46],stage1_31[56],stage1_30[61],stage1_29[131],stage1_28[192]}
   );
   gpc606_5 gpc1112 (
      {stage0_28[312], stage0_28[313], stage0_28[314], stage0_28[315], stage0_28[316], stage0_28[317]},
      {stage0_30[282], stage0_30[283], stage0_30[284], stage0_30[285], stage0_30[286], stage0_30[287]},
      {stage1_32[47],stage1_31[57],stage1_30[62],stage1_29[132],stage1_28[193]}
   );
   gpc606_5 gpc1113 (
      {stage0_28[318], stage0_28[319], stage0_28[320], stage0_28[321], stage0_28[322], stage0_28[323]},
      {stage0_30[288], stage0_30[289], stage0_30[290], stage0_30[291], stage0_30[292], stage0_30[293]},
      {stage1_32[48],stage1_31[58],stage1_30[63],stage1_29[133],stage1_28[194]}
   );
   gpc606_5 gpc1114 (
      {stage0_28[324], stage0_28[325], stage0_28[326], stage0_28[327], stage0_28[328], stage0_28[329]},
      {stage0_30[294], stage0_30[295], stage0_30[296], stage0_30[297], stage0_30[298], stage0_30[299]},
      {stage1_32[49],stage1_31[59],stage1_30[64],stage1_29[134],stage1_28[195]}
   );
   gpc606_5 gpc1115 (
      {stage0_28[330], stage0_28[331], stage0_28[332], stage0_28[333], stage0_28[334], stage0_28[335]},
      {stage0_30[300], stage0_30[301], stage0_30[302], stage0_30[303], stage0_30[304], stage0_30[305]},
      {stage1_32[50],stage1_31[60],stage1_30[65],stage1_29[135],stage1_28[196]}
   );
   gpc606_5 gpc1116 (
      {stage0_28[336], stage0_28[337], stage0_28[338], stage0_28[339], stage0_28[340], stage0_28[341]},
      {stage0_30[306], stage0_30[307], stage0_30[308], stage0_30[309], stage0_30[310], stage0_30[311]},
      {stage1_32[51],stage1_31[61],stage1_30[66],stage1_29[136],stage1_28[197]}
   );
   gpc606_5 gpc1117 (
      {stage0_28[342], stage0_28[343], stage0_28[344], stage0_28[345], stage0_28[346], stage0_28[347]},
      {stage0_30[312], stage0_30[313], stage0_30[314], stage0_30[315], stage0_30[316], stage0_30[317]},
      {stage1_32[52],stage1_31[62],stage1_30[67],stage1_29[137],stage1_28[198]}
   );
   gpc606_5 gpc1118 (
      {stage0_28[348], stage0_28[349], stage0_28[350], stage0_28[351], stage0_28[352], stage0_28[353]},
      {stage0_30[318], stage0_30[319], stage0_30[320], stage0_30[321], stage0_30[322], stage0_30[323]},
      {stage1_32[53],stage1_31[63],stage1_30[68],stage1_29[138],stage1_28[199]}
   );
   gpc606_5 gpc1119 (
      {stage0_28[354], stage0_28[355], stage0_28[356], stage0_28[357], stage0_28[358], stage0_28[359]},
      {stage0_30[324], stage0_30[325], stage0_30[326], stage0_30[327], stage0_30[328], stage0_30[329]},
      {stage1_32[54],stage1_31[64],stage1_30[69],stage1_29[139],stage1_28[200]}
   );
   gpc606_5 gpc1120 (
      {stage0_28[360], stage0_28[361], stage0_28[362], stage0_28[363], stage0_28[364], stage0_28[365]},
      {stage0_30[330], stage0_30[331], stage0_30[332], stage0_30[333], stage0_30[334], stage0_30[335]},
      {stage1_32[55],stage1_31[65],stage1_30[70],stage1_29[140],stage1_28[201]}
   );
   gpc606_5 gpc1121 (
      {stage0_28[366], stage0_28[367], stage0_28[368], stage0_28[369], stage0_28[370], stage0_28[371]},
      {stage0_30[336], stage0_30[337], stage0_30[338], stage0_30[339], stage0_30[340], stage0_30[341]},
      {stage1_32[56],stage1_31[66],stage1_30[71],stage1_29[141],stage1_28[202]}
   );
   gpc606_5 gpc1122 (
      {stage0_28[372], stage0_28[373], stage0_28[374], stage0_28[375], stage0_28[376], stage0_28[377]},
      {stage0_30[342], stage0_30[343], stage0_30[344], stage0_30[345], stage0_30[346], stage0_30[347]},
      {stage1_32[57],stage1_31[67],stage1_30[72],stage1_29[142],stage1_28[203]}
   );
   gpc606_5 gpc1123 (
      {stage0_28[378], stage0_28[379], stage0_28[380], stage0_28[381], stage0_28[382], stage0_28[383]},
      {stage0_30[348], stage0_30[349], stage0_30[350], stage0_30[351], stage0_30[352], stage0_30[353]},
      {stage1_32[58],stage1_31[68],stage1_30[73],stage1_29[143],stage1_28[204]}
   );
   gpc606_5 gpc1124 (
      {stage0_28[384], stage0_28[385], stage0_28[386], stage0_28[387], stage0_28[388], stage0_28[389]},
      {stage0_30[354], stage0_30[355], stage0_30[356], stage0_30[357], stage0_30[358], stage0_30[359]},
      {stage1_32[59],stage1_31[69],stage1_30[74],stage1_29[144],stage1_28[205]}
   );
   gpc606_5 gpc1125 (
      {stage0_28[390], stage0_28[391], stage0_28[392], stage0_28[393], stage0_28[394], stage0_28[395]},
      {stage0_30[360], stage0_30[361], stage0_30[362], stage0_30[363], stage0_30[364], stage0_30[365]},
      {stage1_32[60],stage1_31[70],stage1_30[75],stage1_29[145],stage1_28[206]}
   );
   gpc606_5 gpc1126 (
      {stage0_28[396], stage0_28[397], stage0_28[398], stage0_28[399], stage0_28[400], stage0_28[401]},
      {stage0_30[366], stage0_30[367], stage0_30[368], stage0_30[369], stage0_30[370], stage0_30[371]},
      {stage1_32[61],stage1_31[71],stage1_30[76],stage1_29[146],stage1_28[207]}
   );
   gpc606_5 gpc1127 (
      {stage0_28[402], stage0_28[403], stage0_28[404], stage0_28[405], stage0_28[406], stage0_28[407]},
      {stage0_30[372], stage0_30[373], stage0_30[374], stage0_30[375], stage0_30[376], stage0_30[377]},
      {stage1_32[62],stage1_31[72],stage1_30[77],stage1_29[147],stage1_28[208]}
   );
   gpc606_5 gpc1128 (
      {stage0_28[408], stage0_28[409], stage0_28[410], stage0_28[411], stage0_28[412], stage0_28[413]},
      {stage0_30[378], stage0_30[379], stage0_30[380], stage0_30[381], stage0_30[382], stage0_30[383]},
      {stage1_32[63],stage1_31[73],stage1_30[78],stage1_29[148],stage1_28[209]}
   );
   gpc606_5 gpc1129 (
      {stage0_28[414], stage0_28[415], stage0_28[416], stage0_28[417], stage0_28[418], stage0_28[419]},
      {stage0_30[384], stage0_30[385], stage0_30[386], stage0_30[387], stage0_30[388], stage0_30[389]},
      {stage1_32[64],stage1_31[74],stage1_30[79],stage1_29[149],stage1_28[210]}
   );
   gpc606_5 gpc1130 (
      {stage0_28[420], stage0_28[421], stage0_28[422], stage0_28[423], stage0_28[424], stage0_28[425]},
      {stage0_30[390], stage0_30[391], stage0_30[392], stage0_30[393], stage0_30[394], stage0_30[395]},
      {stage1_32[65],stage1_31[75],stage1_30[80],stage1_29[150],stage1_28[211]}
   );
   gpc606_5 gpc1131 (
      {stage0_28[426], stage0_28[427], stage0_28[428], stage0_28[429], stage0_28[430], stage0_28[431]},
      {stage0_30[396], stage0_30[397], stage0_30[398], stage0_30[399], stage0_30[400], stage0_30[401]},
      {stage1_32[66],stage1_31[76],stage1_30[81],stage1_29[151],stage1_28[212]}
   );
   gpc606_5 gpc1132 (
      {stage0_28[432], stage0_28[433], stage0_28[434], stage0_28[435], stage0_28[436], stage0_28[437]},
      {stage0_30[402], stage0_30[403], stage0_30[404], stage0_30[405], stage0_30[406], stage0_30[407]},
      {stage1_32[67],stage1_31[77],stage1_30[82],stage1_29[152],stage1_28[213]}
   );
   gpc606_5 gpc1133 (
      {stage0_28[438], stage0_28[439], stage0_28[440], stage0_28[441], stage0_28[442], stage0_28[443]},
      {stage0_30[408], stage0_30[409], stage0_30[410], stage0_30[411], stage0_30[412], stage0_30[413]},
      {stage1_32[68],stage1_31[78],stage1_30[83],stage1_29[153],stage1_28[214]}
   );
   gpc606_5 gpc1134 (
      {stage0_28[444], stage0_28[445], stage0_28[446], stage0_28[447], stage0_28[448], stage0_28[449]},
      {stage0_30[414], stage0_30[415], stage0_30[416], stage0_30[417], stage0_30[418], stage0_30[419]},
      {stage1_32[69],stage1_31[79],stage1_30[84],stage1_29[154],stage1_28[215]}
   );
   gpc606_5 gpc1135 (
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[70],stage1_31[80],stage1_30[85],stage1_29[155]}
   );
   gpc606_5 gpc1136 (
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[71],stage1_31[81],stage1_30[86],stage1_29[156]}
   );
   gpc606_5 gpc1137 (
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[72],stage1_31[82],stage1_30[87],stage1_29[157]}
   );
   gpc606_5 gpc1138 (
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[73],stage1_31[83],stage1_30[88],stage1_29[158]}
   );
   gpc606_5 gpc1139 (
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[74],stage1_31[84],stage1_30[89],stage1_29[159]}
   );
   gpc606_5 gpc1140 (
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[75],stage1_31[85],stage1_30[90],stage1_29[160]}
   );
   gpc606_5 gpc1141 (
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[76],stage1_31[86],stage1_30[91],stage1_29[161]}
   );
   gpc606_5 gpc1142 (
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[77],stage1_31[87],stage1_30[92],stage1_29[162]}
   );
   gpc606_5 gpc1143 (
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[78],stage1_31[88],stage1_30[93],stage1_29[163]}
   );
   gpc606_5 gpc1144 (
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[79],stage1_31[89],stage1_30[94],stage1_29[164]}
   );
   gpc606_5 gpc1145 (
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[80],stage1_31[90],stage1_30[95],stage1_29[165]}
   );
   gpc606_5 gpc1146 (
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[81],stage1_31[91],stage1_30[96],stage1_29[166]}
   );
   gpc606_5 gpc1147 (
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[82],stage1_31[92],stage1_30[97],stage1_29[167]}
   );
   gpc606_5 gpc1148 (
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[83],stage1_31[93],stage1_30[98],stage1_29[168]}
   );
   gpc606_5 gpc1149 (
      {stage0_29[144], stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[84],stage1_31[94],stage1_30[99],stage1_29[169]}
   );
   gpc606_5 gpc1150 (
      {stage0_29[150], stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[85],stage1_31[95],stage1_30[100],stage1_29[170]}
   );
   gpc606_5 gpc1151 (
      {stage0_29[156], stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161]},
      {stage0_31[96], stage0_31[97], stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101]},
      {stage1_33[16],stage1_32[86],stage1_31[96],stage1_30[101],stage1_29[171]}
   );
   gpc606_5 gpc1152 (
      {stage0_29[162], stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167]},
      {stage0_31[102], stage0_31[103], stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107]},
      {stage1_33[17],stage1_32[87],stage1_31[97],stage1_30[102],stage1_29[172]}
   );
   gpc606_5 gpc1153 (
      {stage0_29[168], stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173]},
      {stage0_31[108], stage0_31[109], stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113]},
      {stage1_33[18],stage1_32[88],stage1_31[98],stage1_30[103],stage1_29[173]}
   );
   gpc606_5 gpc1154 (
      {stage0_29[174], stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179]},
      {stage0_31[114], stage0_31[115], stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119]},
      {stage1_33[19],stage1_32[89],stage1_31[99],stage1_30[104],stage1_29[174]}
   );
   gpc606_5 gpc1155 (
      {stage0_29[180], stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185]},
      {stage0_31[120], stage0_31[121], stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125]},
      {stage1_33[20],stage1_32[90],stage1_31[100],stage1_30[105],stage1_29[175]}
   );
   gpc615_5 gpc1156 (
      {stage0_29[186], stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190]},
      {stage0_30[420]},
      {stage0_31[126], stage0_31[127], stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131]},
      {stage1_33[21],stage1_32[91],stage1_31[101],stage1_30[106],stage1_29[176]}
   );
   gpc615_5 gpc1157 (
      {stage0_29[191], stage0_29[192], stage0_29[193], stage0_29[194], stage0_29[195]},
      {stage0_30[421]},
      {stage0_31[132], stage0_31[133], stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137]},
      {stage1_33[22],stage1_32[92],stage1_31[102],stage1_30[107],stage1_29[177]}
   );
   gpc615_5 gpc1158 (
      {stage0_29[196], stage0_29[197], stage0_29[198], stage0_29[199], stage0_29[200]},
      {stage0_30[422]},
      {stage0_31[138], stage0_31[139], stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143]},
      {stage1_33[23],stage1_32[93],stage1_31[103],stage1_30[108],stage1_29[178]}
   );
   gpc615_5 gpc1159 (
      {stage0_29[201], stage0_29[202], stage0_29[203], stage0_29[204], stage0_29[205]},
      {stage0_30[423]},
      {stage0_31[144], stage0_31[145], stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149]},
      {stage1_33[24],stage1_32[94],stage1_31[104],stage1_30[109],stage1_29[179]}
   );
   gpc615_5 gpc1160 (
      {stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209], stage0_29[210]},
      {stage0_30[424]},
      {stage0_31[150], stage0_31[151], stage0_31[152], stage0_31[153], stage0_31[154], stage0_31[155]},
      {stage1_33[25],stage1_32[95],stage1_31[105],stage1_30[110],stage1_29[180]}
   );
   gpc615_5 gpc1161 (
      {stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215]},
      {stage0_30[425]},
      {stage0_31[156], stage0_31[157], stage0_31[158], stage0_31[159], stage0_31[160], stage0_31[161]},
      {stage1_33[26],stage1_32[96],stage1_31[106],stage1_30[111],stage1_29[181]}
   );
   gpc615_5 gpc1162 (
      {stage0_29[216], stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220]},
      {stage0_30[426]},
      {stage0_31[162], stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage1_33[27],stage1_32[97],stage1_31[107],stage1_30[112],stage1_29[182]}
   );
   gpc615_5 gpc1163 (
      {stage0_29[221], stage0_29[222], stage0_29[223], stage0_29[224], stage0_29[225]},
      {stage0_30[427]},
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172], stage0_31[173]},
      {stage1_33[28],stage1_32[98],stage1_31[108],stage1_30[113],stage1_29[183]}
   );
   gpc615_5 gpc1164 (
      {stage0_29[226], stage0_29[227], stage0_29[228], stage0_29[229], stage0_29[230]},
      {stage0_30[428]},
      {stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177], stage0_31[178], stage0_31[179]},
      {stage1_33[29],stage1_32[99],stage1_31[109],stage1_30[114],stage1_29[184]}
   );
   gpc615_5 gpc1165 (
      {stage0_29[231], stage0_29[232], stage0_29[233], stage0_29[234], stage0_29[235]},
      {stage0_30[429]},
      {stage0_31[180], stage0_31[181], stage0_31[182], stage0_31[183], stage0_31[184], stage0_31[185]},
      {stage1_33[30],stage1_32[100],stage1_31[110],stage1_30[115],stage1_29[185]}
   );
   gpc615_5 gpc1166 (
      {stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239], stage0_29[240]},
      {stage0_30[430]},
      {stage0_31[186], stage0_31[187], stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191]},
      {stage1_33[31],stage1_32[101],stage1_31[111],stage1_30[116],stage1_29[186]}
   );
   gpc615_5 gpc1167 (
      {stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245]},
      {stage0_30[431]},
      {stage0_31[192], stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage1_33[32],stage1_32[102],stage1_31[112],stage1_30[117],stage1_29[187]}
   );
   gpc615_5 gpc1168 (
      {stage0_29[246], stage0_29[247], stage0_29[248], stage0_29[249], stage0_29[250]},
      {stage0_30[432]},
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202], stage0_31[203]},
      {stage1_33[33],stage1_32[103],stage1_31[113],stage1_30[118],stage1_29[188]}
   );
   gpc615_5 gpc1169 (
      {stage0_29[251], stage0_29[252], stage0_29[253], stage0_29[254], stage0_29[255]},
      {stage0_30[433]},
      {stage0_31[204], stage0_31[205], stage0_31[206], stage0_31[207], stage0_31[208], stage0_31[209]},
      {stage1_33[34],stage1_32[104],stage1_31[114],stage1_30[119],stage1_29[189]}
   );
   gpc615_5 gpc1170 (
      {stage0_29[256], stage0_29[257], stage0_29[258], stage0_29[259], stage0_29[260]},
      {stage0_30[434]},
      {stage0_31[210], stage0_31[211], stage0_31[212], stage0_31[213], stage0_31[214], stage0_31[215]},
      {stage1_33[35],stage1_32[105],stage1_31[115],stage1_30[120],stage1_29[190]}
   );
   gpc615_5 gpc1171 (
      {stage0_29[261], stage0_29[262], stage0_29[263], stage0_29[264], stage0_29[265]},
      {stage0_30[435]},
      {stage0_31[216], stage0_31[217], stage0_31[218], stage0_31[219], stage0_31[220], stage0_31[221]},
      {stage1_33[36],stage1_32[106],stage1_31[116],stage1_30[121],stage1_29[191]}
   );
   gpc615_5 gpc1172 (
      {stage0_29[266], stage0_29[267], stage0_29[268], stage0_29[269], stage0_29[270]},
      {stage0_30[436]},
      {stage0_31[222], stage0_31[223], stage0_31[224], stage0_31[225], stage0_31[226], stage0_31[227]},
      {stage1_33[37],stage1_32[107],stage1_31[117],stage1_30[122],stage1_29[192]}
   );
   gpc615_5 gpc1173 (
      {stage0_29[271], stage0_29[272], stage0_29[273], stage0_29[274], stage0_29[275]},
      {stage0_30[437]},
      {stage0_31[228], stage0_31[229], stage0_31[230], stage0_31[231], stage0_31[232], stage0_31[233]},
      {stage1_33[38],stage1_32[108],stage1_31[118],stage1_30[123],stage1_29[193]}
   );
   gpc615_5 gpc1174 (
      {stage0_29[276], stage0_29[277], stage0_29[278], stage0_29[279], stage0_29[280]},
      {stage0_30[438]},
      {stage0_31[234], stage0_31[235], stage0_31[236], stage0_31[237], stage0_31[238], stage0_31[239]},
      {stage1_33[39],stage1_32[109],stage1_31[119],stage1_30[124],stage1_29[194]}
   );
   gpc615_5 gpc1175 (
      {stage0_29[281], stage0_29[282], stage0_29[283], stage0_29[284], stage0_29[285]},
      {stage0_30[439]},
      {stage0_31[240], stage0_31[241], stage0_31[242], stage0_31[243], stage0_31[244], stage0_31[245]},
      {stage1_33[40],stage1_32[110],stage1_31[120],stage1_30[125],stage1_29[195]}
   );
   gpc615_5 gpc1176 (
      {stage0_29[286], stage0_29[287], stage0_29[288], stage0_29[289], stage0_29[290]},
      {stage0_30[440]},
      {stage0_31[246], stage0_31[247], stage0_31[248], stage0_31[249], stage0_31[250], stage0_31[251]},
      {stage1_33[41],stage1_32[111],stage1_31[121],stage1_30[126],stage1_29[196]}
   );
   gpc615_5 gpc1177 (
      {stage0_29[291], stage0_29[292], stage0_29[293], stage0_29[294], stage0_29[295]},
      {stage0_30[441]},
      {stage0_31[252], stage0_31[253], stage0_31[254], stage0_31[255], stage0_31[256], stage0_31[257]},
      {stage1_33[42],stage1_32[112],stage1_31[122],stage1_30[127],stage1_29[197]}
   );
   gpc615_5 gpc1178 (
      {stage0_29[296], stage0_29[297], stage0_29[298], stage0_29[299], stage0_29[300]},
      {stage0_30[442]},
      {stage0_31[258], stage0_31[259], stage0_31[260], stage0_31[261], stage0_31[262], stage0_31[263]},
      {stage1_33[43],stage1_32[113],stage1_31[123],stage1_30[128],stage1_29[198]}
   );
   gpc615_5 gpc1179 (
      {stage0_29[301], stage0_29[302], stage0_29[303], stage0_29[304], stage0_29[305]},
      {stage0_30[443]},
      {stage0_31[264], stage0_31[265], stage0_31[266], stage0_31[267], stage0_31[268], stage0_31[269]},
      {stage1_33[44],stage1_32[114],stage1_31[124],stage1_30[129],stage1_29[199]}
   );
   gpc615_5 gpc1180 (
      {stage0_29[306], stage0_29[307], stage0_29[308], stage0_29[309], stage0_29[310]},
      {stage0_30[444]},
      {stage0_31[270], stage0_31[271], stage0_31[272], stage0_31[273], stage0_31[274], stage0_31[275]},
      {stage1_33[45],stage1_32[115],stage1_31[125],stage1_30[130],stage1_29[200]}
   );
   gpc615_5 gpc1181 (
      {stage0_29[311], stage0_29[312], stage0_29[313], stage0_29[314], stage0_29[315]},
      {stage0_30[445]},
      {stage0_31[276], stage0_31[277], stage0_31[278], stage0_31[279], stage0_31[280], stage0_31[281]},
      {stage1_33[46],stage1_32[116],stage1_31[126],stage1_30[131],stage1_29[201]}
   );
   gpc615_5 gpc1182 (
      {stage0_29[316], stage0_29[317], stage0_29[318], stage0_29[319], stage0_29[320]},
      {stage0_30[446]},
      {stage0_31[282], stage0_31[283], stage0_31[284], stage0_31[285], stage0_31[286], stage0_31[287]},
      {stage1_33[47],stage1_32[117],stage1_31[127],stage1_30[132],stage1_29[202]}
   );
   gpc615_5 gpc1183 (
      {stage0_29[321], stage0_29[322], stage0_29[323], stage0_29[324], stage0_29[325]},
      {stage0_30[447]},
      {stage0_31[288], stage0_31[289], stage0_31[290], stage0_31[291], stage0_31[292], stage0_31[293]},
      {stage1_33[48],stage1_32[118],stage1_31[128],stage1_30[133],stage1_29[203]}
   );
   gpc615_5 gpc1184 (
      {stage0_29[326], stage0_29[327], stage0_29[328], stage0_29[329], stage0_29[330]},
      {stage0_30[448]},
      {stage0_31[294], stage0_31[295], stage0_31[296], stage0_31[297], stage0_31[298], stage0_31[299]},
      {stage1_33[49],stage1_32[119],stage1_31[129],stage1_30[134],stage1_29[204]}
   );
   gpc615_5 gpc1185 (
      {stage0_29[331], stage0_29[332], stage0_29[333], stage0_29[334], stage0_29[335]},
      {stage0_30[449]},
      {stage0_31[300], stage0_31[301], stage0_31[302], stage0_31[303], stage0_31[304], stage0_31[305]},
      {stage1_33[50],stage1_32[120],stage1_31[130],stage1_30[135],stage1_29[205]}
   );
   gpc615_5 gpc1186 (
      {stage0_29[336], stage0_29[337], stage0_29[338], stage0_29[339], stage0_29[340]},
      {stage0_30[450]},
      {stage0_31[306], stage0_31[307], stage0_31[308], stage0_31[309], stage0_31[310], stage0_31[311]},
      {stage1_33[51],stage1_32[121],stage1_31[131],stage1_30[136],stage1_29[206]}
   );
   gpc615_5 gpc1187 (
      {stage0_29[341], stage0_29[342], stage0_29[343], stage0_29[344], stage0_29[345]},
      {stage0_30[451]},
      {stage0_31[312], stage0_31[313], stage0_31[314], stage0_31[315], stage0_31[316], stage0_31[317]},
      {stage1_33[52],stage1_32[122],stage1_31[132],stage1_30[137],stage1_29[207]}
   );
   gpc615_5 gpc1188 (
      {stage0_29[346], stage0_29[347], stage0_29[348], stage0_29[349], stage0_29[350]},
      {stage0_30[452]},
      {stage0_31[318], stage0_31[319], stage0_31[320], stage0_31[321], stage0_31[322], stage0_31[323]},
      {stage1_33[53],stage1_32[123],stage1_31[133],stage1_30[138],stage1_29[208]}
   );
   gpc615_5 gpc1189 (
      {stage0_29[351], stage0_29[352], stage0_29[353], stage0_29[354], stage0_29[355]},
      {stage0_30[453]},
      {stage0_31[324], stage0_31[325], stage0_31[326], stage0_31[327], stage0_31[328], stage0_31[329]},
      {stage1_33[54],stage1_32[124],stage1_31[134],stage1_30[139],stage1_29[209]}
   );
   gpc615_5 gpc1190 (
      {stage0_29[356], stage0_29[357], stage0_29[358], stage0_29[359], stage0_29[360]},
      {stage0_30[454]},
      {stage0_31[330], stage0_31[331], stage0_31[332], stage0_31[333], stage0_31[334], stage0_31[335]},
      {stage1_33[55],stage1_32[125],stage1_31[135],stage1_30[140],stage1_29[210]}
   );
   gpc615_5 gpc1191 (
      {stage0_29[361], stage0_29[362], stage0_29[363], stage0_29[364], stage0_29[365]},
      {stage0_30[455]},
      {stage0_31[336], stage0_31[337], stage0_31[338], stage0_31[339], stage0_31[340], stage0_31[341]},
      {stage1_33[56],stage1_32[126],stage1_31[136],stage1_30[141],stage1_29[211]}
   );
   gpc615_5 gpc1192 (
      {stage0_29[366], stage0_29[367], stage0_29[368], stage0_29[369], stage0_29[370]},
      {stage0_30[456]},
      {stage0_31[342], stage0_31[343], stage0_31[344], stage0_31[345], stage0_31[346], stage0_31[347]},
      {stage1_33[57],stage1_32[127],stage1_31[137],stage1_30[142],stage1_29[212]}
   );
   gpc615_5 gpc1193 (
      {stage0_29[371], stage0_29[372], stage0_29[373], stage0_29[374], stage0_29[375]},
      {stage0_30[457]},
      {stage0_31[348], stage0_31[349], stage0_31[350], stage0_31[351], stage0_31[352], stage0_31[353]},
      {stage1_33[58],stage1_32[128],stage1_31[138],stage1_30[143],stage1_29[213]}
   );
   gpc615_5 gpc1194 (
      {stage0_29[376], stage0_29[377], stage0_29[378], stage0_29[379], stage0_29[380]},
      {stage0_30[458]},
      {stage0_31[354], stage0_31[355], stage0_31[356], stage0_31[357], stage0_31[358], stage0_31[359]},
      {stage1_33[59],stage1_32[129],stage1_31[139],stage1_30[144],stage1_29[214]}
   );
   gpc615_5 gpc1195 (
      {stage0_29[381], stage0_29[382], stage0_29[383], stage0_29[384], stage0_29[385]},
      {stage0_30[459]},
      {stage0_31[360], stage0_31[361], stage0_31[362], stage0_31[363], stage0_31[364], stage0_31[365]},
      {stage1_33[60],stage1_32[130],stage1_31[140],stage1_30[145],stage1_29[215]}
   );
   gpc615_5 gpc1196 (
      {stage0_29[386], stage0_29[387], stage0_29[388], stage0_29[389], stage0_29[390]},
      {stage0_30[460]},
      {stage0_31[366], stage0_31[367], stage0_31[368], stage0_31[369], stage0_31[370], stage0_31[371]},
      {stage1_33[61],stage1_32[131],stage1_31[141],stage1_30[146],stage1_29[216]}
   );
   gpc615_5 gpc1197 (
      {stage0_29[391], stage0_29[392], stage0_29[393], stage0_29[394], stage0_29[395]},
      {stage0_30[461]},
      {stage0_31[372], stage0_31[373], stage0_31[374], stage0_31[375], stage0_31[376], stage0_31[377]},
      {stage1_33[62],stage1_32[132],stage1_31[142],stage1_30[147],stage1_29[217]}
   );
   gpc615_5 gpc1198 (
      {stage0_29[396], stage0_29[397], stage0_29[398], stage0_29[399], stage0_29[400]},
      {stage0_30[462]},
      {stage0_31[378], stage0_31[379], stage0_31[380], stage0_31[381], stage0_31[382], stage0_31[383]},
      {stage1_33[63],stage1_32[133],stage1_31[143],stage1_30[148],stage1_29[218]}
   );
   gpc615_5 gpc1199 (
      {stage0_29[401], stage0_29[402], stage0_29[403], stage0_29[404], stage0_29[405]},
      {stage0_30[463]},
      {stage0_31[384], stage0_31[385], stage0_31[386], stage0_31[387], stage0_31[388], stage0_31[389]},
      {stage1_33[64],stage1_32[134],stage1_31[144],stage1_30[149],stage1_29[219]}
   );
   gpc615_5 gpc1200 (
      {stage0_29[406], stage0_29[407], stage0_29[408], stage0_29[409], stage0_29[410]},
      {stage0_30[464]},
      {stage0_31[390], stage0_31[391], stage0_31[392], stage0_31[393], stage0_31[394], stage0_31[395]},
      {stage1_33[65],stage1_32[135],stage1_31[145],stage1_30[150],stage1_29[220]}
   );
   gpc615_5 gpc1201 (
      {stage0_29[411], stage0_29[412], stage0_29[413], stage0_29[414], stage0_29[415]},
      {stage0_30[465]},
      {stage0_31[396], stage0_31[397], stage0_31[398], stage0_31[399], stage0_31[400], stage0_31[401]},
      {stage1_33[66],stage1_32[136],stage1_31[146],stage1_30[151],stage1_29[221]}
   );
   gpc615_5 gpc1202 (
      {stage0_29[416], stage0_29[417], stage0_29[418], stage0_29[419], stage0_29[420]},
      {stage0_30[466]},
      {stage0_31[402], stage0_31[403], stage0_31[404], stage0_31[405], stage0_31[406], stage0_31[407]},
      {stage1_33[67],stage1_32[137],stage1_31[147],stage1_30[152],stage1_29[222]}
   );
   gpc615_5 gpc1203 (
      {stage0_29[421], stage0_29[422], stage0_29[423], stage0_29[424], stage0_29[425]},
      {stage0_30[467]},
      {stage0_31[408], stage0_31[409], stage0_31[410], stage0_31[411], stage0_31[412], stage0_31[413]},
      {stage1_33[68],stage1_32[138],stage1_31[148],stage1_30[153],stage1_29[223]}
   );
   gpc615_5 gpc1204 (
      {stage0_29[426], stage0_29[427], stage0_29[428], stage0_29[429], stage0_29[430]},
      {stage0_30[468]},
      {stage0_31[414], stage0_31[415], stage0_31[416], stage0_31[417], stage0_31[418], stage0_31[419]},
      {stage1_33[69],stage1_32[139],stage1_31[149],stage1_30[154],stage1_29[224]}
   );
   gpc615_5 gpc1205 (
      {stage0_29[431], stage0_29[432], stage0_29[433], stage0_29[434], stage0_29[435]},
      {stage0_30[469]},
      {stage0_31[420], stage0_31[421], stage0_31[422], stage0_31[423], stage0_31[424], stage0_31[425]},
      {stage1_33[70],stage1_32[140],stage1_31[150],stage1_30[155],stage1_29[225]}
   );
   gpc615_5 gpc1206 (
      {stage0_29[436], stage0_29[437], stage0_29[438], stage0_29[439], stage0_29[440]},
      {stage0_30[470]},
      {stage0_31[426], stage0_31[427], stage0_31[428], stage0_31[429], stage0_31[430], stage0_31[431]},
      {stage1_33[71],stage1_32[141],stage1_31[151],stage1_30[156],stage1_29[226]}
   );
   gpc615_5 gpc1207 (
      {stage0_29[441], stage0_29[442], stage0_29[443], stage0_29[444], stage0_29[445]},
      {stage0_30[471]},
      {stage0_31[432], stage0_31[433], stage0_31[434], stage0_31[435], stage0_31[436], stage0_31[437]},
      {stage1_33[72],stage1_32[142],stage1_31[152],stage1_30[157],stage1_29[227]}
   );
   gpc615_5 gpc1208 (
      {stage0_29[446], stage0_29[447], stage0_29[448], stage0_29[449], stage0_29[450]},
      {stage0_30[472]},
      {stage0_31[438], stage0_31[439], stage0_31[440], stage0_31[441], stage0_31[442], stage0_31[443]},
      {stage1_33[73],stage1_32[143],stage1_31[153],stage1_30[158],stage1_29[228]}
   );
   gpc615_5 gpc1209 (
      {stage0_29[451], stage0_29[452], stage0_29[453], stage0_29[454], stage0_29[455]},
      {stage0_30[473]},
      {stage0_31[444], stage0_31[445], stage0_31[446], stage0_31[447], stage0_31[448], stage0_31[449]},
      {stage1_33[74],stage1_32[144],stage1_31[154],stage1_30[159],stage1_29[229]}
   );
   gpc615_5 gpc1210 (
      {stage0_29[456], stage0_29[457], stage0_29[458], stage0_29[459], stage0_29[460]},
      {stage0_30[474]},
      {stage0_31[450], stage0_31[451], stage0_31[452], stage0_31[453], stage0_31[454], stage0_31[455]},
      {stage1_33[75],stage1_32[145],stage1_31[155],stage1_30[160],stage1_29[230]}
   );
   gpc615_5 gpc1211 (
      {stage0_29[461], stage0_29[462], stage0_29[463], stage0_29[464], stage0_29[465]},
      {stage0_30[475]},
      {stage0_31[456], stage0_31[457], stage0_31[458], stage0_31[459], stage0_31[460], stage0_31[461]},
      {stage1_33[76],stage1_32[146],stage1_31[156],stage1_30[161],stage1_29[231]}
   );
   gpc615_5 gpc1212 (
      {stage0_29[466], stage0_29[467], stage0_29[468], stage0_29[469], stage0_29[470]},
      {stage0_30[476]},
      {stage0_31[462], stage0_31[463], stage0_31[464], stage0_31[465], stage0_31[466], stage0_31[467]},
      {stage1_33[77],stage1_32[147],stage1_31[157],stage1_30[162],stage1_29[232]}
   );
   gpc615_5 gpc1213 (
      {stage0_29[471], stage0_29[472], stage0_29[473], stage0_29[474], stage0_29[475]},
      {stage0_30[477]},
      {stage0_31[468], stage0_31[469], stage0_31[470], stage0_31[471], stage0_31[472], stage0_31[473]},
      {stage1_33[78],stage1_32[148],stage1_31[158],stage1_30[163],stage1_29[233]}
   );
   gpc615_5 gpc1214 (
      {stage0_29[476], stage0_29[477], stage0_29[478], stage0_29[479], stage0_29[480]},
      {stage0_30[478]},
      {stage0_31[474], stage0_31[475], stage0_31[476], stage0_31[477], stage0_31[478], stage0_31[479]},
      {stage1_33[79],stage1_32[149],stage1_31[159],stage1_30[164],stage1_29[234]}
   );
   gpc615_5 gpc1215 (
      {stage0_29[481], stage0_29[482], stage0_29[483], stage0_29[484], stage0_29[485]},
      {stage0_30[479]},
      {stage0_31[480], stage0_31[481], stage0_31[482], stage0_31[483], stage0_31[484], stage0_31[485]},
      {stage1_33[80],stage1_32[150],stage1_31[160],stage1_30[165],stage1_29[235]}
   );
   gpc1_1 gpc1216 (
      {stage0_0[444]},
      {stage1_0[85]}
   );
   gpc1_1 gpc1217 (
      {stage0_0[445]},
      {stage1_0[86]}
   );
   gpc1_1 gpc1218 (
      {stage0_0[446]},
      {stage1_0[87]}
   );
   gpc1_1 gpc1219 (
      {stage0_0[447]},
      {stage1_0[88]}
   );
   gpc1_1 gpc1220 (
      {stage0_0[448]},
      {stage1_0[89]}
   );
   gpc1_1 gpc1221 (
      {stage0_0[449]},
      {stage1_0[90]}
   );
   gpc1_1 gpc1222 (
      {stage0_0[450]},
      {stage1_0[91]}
   );
   gpc1_1 gpc1223 (
      {stage0_0[451]},
      {stage1_0[92]}
   );
   gpc1_1 gpc1224 (
      {stage0_0[452]},
      {stage1_0[93]}
   );
   gpc1_1 gpc1225 (
      {stage0_0[453]},
      {stage1_0[94]}
   );
   gpc1_1 gpc1226 (
      {stage0_0[454]},
      {stage1_0[95]}
   );
   gpc1_1 gpc1227 (
      {stage0_0[455]},
      {stage1_0[96]}
   );
   gpc1_1 gpc1228 (
      {stage0_0[456]},
      {stage1_0[97]}
   );
   gpc1_1 gpc1229 (
      {stage0_0[457]},
      {stage1_0[98]}
   );
   gpc1_1 gpc1230 (
      {stage0_0[458]},
      {stage1_0[99]}
   );
   gpc1_1 gpc1231 (
      {stage0_0[459]},
      {stage1_0[100]}
   );
   gpc1_1 gpc1232 (
      {stage0_0[460]},
      {stage1_0[101]}
   );
   gpc1_1 gpc1233 (
      {stage0_0[461]},
      {stage1_0[102]}
   );
   gpc1_1 gpc1234 (
      {stage0_0[462]},
      {stage1_0[103]}
   );
   gpc1_1 gpc1235 (
      {stage0_0[463]},
      {stage1_0[104]}
   );
   gpc1_1 gpc1236 (
      {stage0_0[464]},
      {stage1_0[105]}
   );
   gpc1_1 gpc1237 (
      {stage0_0[465]},
      {stage1_0[106]}
   );
   gpc1_1 gpc1238 (
      {stage0_0[466]},
      {stage1_0[107]}
   );
   gpc1_1 gpc1239 (
      {stage0_0[467]},
      {stage1_0[108]}
   );
   gpc1_1 gpc1240 (
      {stage0_0[468]},
      {stage1_0[109]}
   );
   gpc1_1 gpc1241 (
      {stage0_0[469]},
      {stage1_0[110]}
   );
   gpc1_1 gpc1242 (
      {stage0_0[470]},
      {stage1_0[111]}
   );
   gpc1_1 gpc1243 (
      {stage0_0[471]},
      {stage1_0[112]}
   );
   gpc1_1 gpc1244 (
      {stage0_0[472]},
      {stage1_0[113]}
   );
   gpc1_1 gpc1245 (
      {stage0_0[473]},
      {stage1_0[114]}
   );
   gpc1_1 gpc1246 (
      {stage0_0[474]},
      {stage1_0[115]}
   );
   gpc1_1 gpc1247 (
      {stage0_0[475]},
      {stage1_0[116]}
   );
   gpc1_1 gpc1248 (
      {stage0_0[476]},
      {stage1_0[117]}
   );
   gpc1_1 gpc1249 (
      {stage0_0[477]},
      {stage1_0[118]}
   );
   gpc1_1 gpc1250 (
      {stage0_0[478]},
      {stage1_0[119]}
   );
   gpc1_1 gpc1251 (
      {stage0_0[479]},
      {stage1_0[120]}
   );
   gpc1_1 gpc1252 (
      {stage0_0[480]},
      {stage1_0[121]}
   );
   gpc1_1 gpc1253 (
      {stage0_0[481]},
      {stage1_0[122]}
   );
   gpc1_1 gpc1254 (
      {stage0_0[482]},
      {stage1_0[123]}
   );
   gpc1_1 gpc1255 (
      {stage0_0[483]},
      {stage1_0[124]}
   );
   gpc1_1 gpc1256 (
      {stage0_0[484]},
      {stage1_0[125]}
   );
   gpc1_1 gpc1257 (
      {stage0_0[485]},
      {stage1_0[126]}
   );
   gpc1_1 gpc1258 (
      {stage0_1[484]},
      {stage1_1[136]}
   );
   gpc1_1 gpc1259 (
      {stage0_1[485]},
      {stage1_1[137]}
   );
   gpc1_1 gpc1260 (
      {stage0_2[415]},
      {stage1_2[157]}
   );
   gpc1_1 gpc1261 (
      {stage0_2[416]},
      {stage1_2[158]}
   );
   gpc1_1 gpc1262 (
      {stage0_2[417]},
      {stage1_2[159]}
   );
   gpc1_1 gpc1263 (
      {stage0_2[418]},
      {stage1_2[160]}
   );
   gpc1_1 gpc1264 (
      {stage0_2[419]},
      {stage1_2[161]}
   );
   gpc1_1 gpc1265 (
      {stage0_2[420]},
      {stage1_2[162]}
   );
   gpc1_1 gpc1266 (
      {stage0_2[421]},
      {stage1_2[163]}
   );
   gpc1_1 gpc1267 (
      {stage0_2[422]},
      {stage1_2[164]}
   );
   gpc1_1 gpc1268 (
      {stage0_2[423]},
      {stage1_2[165]}
   );
   gpc1_1 gpc1269 (
      {stage0_2[424]},
      {stage1_2[166]}
   );
   gpc1_1 gpc1270 (
      {stage0_2[425]},
      {stage1_2[167]}
   );
   gpc1_1 gpc1271 (
      {stage0_2[426]},
      {stage1_2[168]}
   );
   gpc1_1 gpc1272 (
      {stage0_2[427]},
      {stage1_2[169]}
   );
   gpc1_1 gpc1273 (
      {stage0_2[428]},
      {stage1_2[170]}
   );
   gpc1_1 gpc1274 (
      {stage0_2[429]},
      {stage1_2[171]}
   );
   gpc1_1 gpc1275 (
      {stage0_2[430]},
      {stage1_2[172]}
   );
   gpc1_1 gpc1276 (
      {stage0_2[431]},
      {stage1_2[173]}
   );
   gpc1_1 gpc1277 (
      {stage0_2[432]},
      {stage1_2[174]}
   );
   gpc1_1 gpc1278 (
      {stage0_2[433]},
      {stage1_2[175]}
   );
   gpc1_1 gpc1279 (
      {stage0_2[434]},
      {stage1_2[176]}
   );
   gpc1_1 gpc1280 (
      {stage0_2[435]},
      {stage1_2[177]}
   );
   gpc1_1 gpc1281 (
      {stage0_2[436]},
      {stage1_2[178]}
   );
   gpc1_1 gpc1282 (
      {stage0_2[437]},
      {stage1_2[179]}
   );
   gpc1_1 gpc1283 (
      {stage0_2[438]},
      {stage1_2[180]}
   );
   gpc1_1 gpc1284 (
      {stage0_2[439]},
      {stage1_2[181]}
   );
   gpc1_1 gpc1285 (
      {stage0_2[440]},
      {stage1_2[182]}
   );
   gpc1_1 gpc1286 (
      {stage0_2[441]},
      {stage1_2[183]}
   );
   gpc1_1 gpc1287 (
      {stage0_2[442]},
      {stage1_2[184]}
   );
   gpc1_1 gpc1288 (
      {stage0_2[443]},
      {stage1_2[185]}
   );
   gpc1_1 gpc1289 (
      {stage0_2[444]},
      {stage1_2[186]}
   );
   gpc1_1 gpc1290 (
      {stage0_2[445]},
      {stage1_2[187]}
   );
   gpc1_1 gpc1291 (
      {stage0_2[446]},
      {stage1_2[188]}
   );
   gpc1_1 gpc1292 (
      {stage0_2[447]},
      {stage1_2[189]}
   );
   gpc1_1 gpc1293 (
      {stage0_2[448]},
      {stage1_2[190]}
   );
   gpc1_1 gpc1294 (
      {stage0_2[449]},
      {stage1_2[191]}
   );
   gpc1_1 gpc1295 (
      {stage0_2[450]},
      {stage1_2[192]}
   );
   gpc1_1 gpc1296 (
      {stage0_2[451]},
      {stage1_2[193]}
   );
   gpc1_1 gpc1297 (
      {stage0_2[452]},
      {stage1_2[194]}
   );
   gpc1_1 gpc1298 (
      {stage0_2[453]},
      {stage1_2[195]}
   );
   gpc1_1 gpc1299 (
      {stage0_2[454]},
      {stage1_2[196]}
   );
   gpc1_1 gpc1300 (
      {stage0_2[455]},
      {stage1_2[197]}
   );
   gpc1_1 gpc1301 (
      {stage0_2[456]},
      {stage1_2[198]}
   );
   gpc1_1 gpc1302 (
      {stage0_2[457]},
      {stage1_2[199]}
   );
   gpc1_1 gpc1303 (
      {stage0_2[458]},
      {stage1_2[200]}
   );
   gpc1_1 gpc1304 (
      {stage0_2[459]},
      {stage1_2[201]}
   );
   gpc1_1 gpc1305 (
      {stage0_2[460]},
      {stage1_2[202]}
   );
   gpc1_1 gpc1306 (
      {stage0_2[461]},
      {stage1_2[203]}
   );
   gpc1_1 gpc1307 (
      {stage0_2[462]},
      {stage1_2[204]}
   );
   gpc1_1 gpc1308 (
      {stage0_2[463]},
      {stage1_2[205]}
   );
   gpc1_1 gpc1309 (
      {stage0_2[464]},
      {stage1_2[206]}
   );
   gpc1_1 gpc1310 (
      {stage0_2[465]},
      {stage1_2[207]}
   );
   gpc1_1 gpc1311 (
      {stage0_2[466]},
      {stage1_2[208]}
   );
   gpc1_1 gpc1312 (
      {stage0_2[467]},
      {stage1_2[209]}
   );
   gpc1_1 gpc1313 (
      {stage0_2[468]},
      {stage1_2[210]}
   );
   gpc1_1 gpc1314 (
      {stage0_2[469]},
      {stage1_2[211]}
   );
   gpc1_1 gpc1315 (
      {stage0_2[470]},
      {stage1_2[212]}
   );
   gpc1_1 gpc1316 (
      {stage0_2[471]},
      {stage1_2[213]}
   );
   gpc1_1 gpc1317 (
      {stage0_2[472]},
      {stage1_2[214]}
   );
   gpc1_1 gpc1318 (
      {stage0_2[473]},
      {stage1_2[215]}
   );
   gpc1_1 gpc1319 (
      {stage0_2[474]},
      {stage1_2[216]}
   );
   gpc1_1 gpc1320 (
      {stage0_2[475]},
      {stage1_2[217]}
   );
   gpc1_1 gpc1321 (
      {stage0_2[476]},
      {stage1_2[218]}
   );
   gpc1_1 gpc1322 (
      {stage0_2[477]},
      {stage1_2[219]}
   );
   gpc1_1 gpc1323 (
      {stage0_2[478]},
      {stage1_2[220]}
   );
   gpc1_1 gpc1324 (
      {stage0_2[479]},
      {stage1_2[221]}
   );
   gpc1_1 gpc1325 (
      {stage0_2[480]},
      {stage1_2[222]}
   );
   gpc1_1 gpc1326 (
      {stage0_2[481]},
      {stage1_2[223]}
   );
   gpc1_1 gpc1327 (
      {stage0_2[482]},
      {stage1_2[224]}
   );
   gpc1_1 gpc1328 (
      {stage0_2[483]},
      {stage1_2[225]}
   );
   gpc1_1 gpc1329 (
      {stage0_2[484]},
      {stage1_2[226]}
   );
   gpc1_1 gpc1330 (
      {stage0_2[485]},
      {stage1_2[227]}
   );
   gpc1_1 gpc1331 (
      {stage0_3[484]},
      {stage1_3[186]}
   );
   gpc1_1 gpc1332 (
      {stage0_3[485]},
      {stage1_3[187]}
   );
   gpc1_1 gpc1333 (
      {stage0_4[485]},
      {stage1_4[225]}
   );
   gpc1_1 gpc1334 (
      {stage0_5[474]},
      {stage1_5[206]}
   );
   gpc1_1 gpc1335 (
      {stage0_5[475]},
      {stage1_5[207]}
   );
   gpc1_1 gpc1336 (
      {stage0_5[476]},
      {stage1_5[208]}
   );
   gpc1_1 gpc1337 (
      {stage0_5[477]},
      {stage1_5[209]}
   );
   gpc1_1 gpc1338 (
      {stage0_5[478]},
      {stage1_5[210]}
   );
   gpc1_1 gpc1339 (
      {stage0_5[479]},
      {stage1_5[211]}
   );
   gpc1_1 gpc1340 (
      {stage0_5[480]},
      {stage1_5[212]}
   );
   gpc1_1 gpc1341 (
      {stage0_5[481]},
      {stage1_5[213]}
   );
   gpc1_1 gpc1342 (
      {stage0_5[482]},
      {stage1_5[214]}
   );
   gpc1_1 gpc1343 (
      {stage0_5[483]},
      {stage1_5[215]}
   );
   gpc1_1 gpc1344 (
      {stage0_5[484]},
      {stage1_5[216]}
   );
   gpc1_1 gpc1345 (
      {stage0_5[485]},
      {stage1_5[217]}
   );
   gpc1_1 gpc1346 (
      {stage0_6[410]},
      {stage1_6[171]}
   );
   gpc1_1 gpc1347 (
      {stage0_6[411]},
      {stage1_6[172]}
   );
   gpc1_1 gpc1348 (
      {stage0_6[412]},
      {stage1_6[173]}
   );
   gpc1_1 gpc1349 (
      {stage0_6[413]},
      {stage1_6[174]}
   );
   gpc1_1 gpc1350 (
      {stage0_6[414]},
      {stage1_6[175]}
   );
   gpc1_1 gpc1351 (
      {stage0_6[415]},
      {stage1_6[176]}
   );
   gpc1_1 gpc1352 (
      {stage0_6[416]},
      {stage1_6[177]}
   );
   gpc1_1 gpc1353 (
      {stage0_6[417]},
      {stage1_6[178]}
   );
   gpc1_1 gpc1354 (
      {stage0_6[418]},
      {stage1_6[179]}
   );
   gpc1_1 gpc1355 (
      {stage0_6[419]},
      {stage1_6[180]}
   );
   gpc1_1 gpc1356 (
      {stage0_6[420]},
      {stage1_6[181]}
   );
   gpc1_1 gpc1357 (
      {stage0_6[421]},
      {stage1_6[182]}
   );
   gpc1_1 gpc1358 (
      {stage0_6[422]},
      {stage1_6[183]}
   );
   gpc1_1 gpc1359 (
      {stage0_6[423]},
      {stage1_6[184]}
   );
   gpc1_1 gpc1360 (
      {stage0_6[424]},
      {stage1_6[185]}
   );
   gpc1_1 gpc1361 (
      {stage0_6[425]},
      {stage1_6[186]}
   );
   gpc1_1 gpc1362 (
      {stage0_6[426]},
      {stage1_6[187]}
   );
   gpc1_1 gpc1363 (
      {stage0_6[427]},
      {stage1_6[188]}
   );
   gpc1_1 gpc1364 (
      {stage0_6[428]},
      {stage1_6[189]}
   );
   gpc1_1 gpc1365 (
      {stage0_6[429]},
      {stage1_6[190]}
   );
   gpc1_1 gpc1366 (
      {stage0_6[430]},
      {stage1_6[191]}
   );
   gpc1_1 gpc1367 (
      {stage0_6[431]},
      {stage1_6[192]}
   );
   gpc1_1 gpc1368 (
      {stage0_6[432]},
      {stage1_6[193]}
   );
   gpc1_1 gpc1369 (
      {stage0_6[433]},
      {stage1_6[194]}
   );
   gpc1_1 gpc1370 (
      {stage0_6[434]},
      {stage1_6[195]}
   );
   gpc1_1 gpc1371 (
      {stage0_6[435]},
      {stage1_6[196]}
   );
   gpc1_1 gpc1372 (
      {stage0_6[436]},
      {stage1_6[197]}
   );
   gpc1_1 gpc1373 (
      {stage0_6[437]},
      {stage1_6[198]}
   );
   gpc1_1 gpc1374 (
      {stage0_6[438]},
      {stage1_6[199]}
   );
   gpc1_1 gpc1375 (
      {stage0_6[439]},
      {stage1_6[200]}
   );
   gpc1_1 gpc1376 (
      {stage0_6[440]},
      {stage1_6[201]}
   );
   gpc1_1 gpc1377 (
      {stage0_6[441]},
      {stage1_6[202]}
   );
   gpc1_1 gpc1378 (
      {stage0_6[442]},
      {stage1_6[203]}
   );
   gpc1_1 gpc1379 (
      {stage0_6[443]},
      {stage1_6[204]}
   );
   gpc1_1 gpc1380 (
      {stage0_6[444]},
      {stage1_6[205]}
   );
   gpc1_1 gpc1381 (
      {stage0_6[445]},
      {stage1_6[206]}
   );
   gpc1_1 gpc1382 (
      {stage0_6[446]},
      {stage1_6[207]}
   );
   gpc1_1 gpc1383 (
      {stage0_6[447]},
      {stage1_6[208]}
   );
   gpc1_1 gpc1384 (
      {stage0_6[448]},
      {stage1_6[209]}
   );
   gpc1_1 gpc1385 (
      {stage0_6[449]},
      {stage1_6[210]}
   );
   gpc1_1 gpc1386 (
      {stage0_6[450]},
      {stage1_6[211]}
   );
   gpc1_1 gpc1387 (
      {stage0_6[451]},
      {stage1_6[212]}
   );
   gpc1_1 gpc1388 (
      {stage0_6[452]},
      {stage1_6[213]}
   );
   gpc1_1 gpc1389 (
      {stage0_6[453]},
      {stage1_6[214]}
   );
   gpc1_1 gpc1390 (
      {stage0_6[454]},
      {stage1_6[215]}
   );
   gpc1_1 gpc1391 (
      {stage0_6[455]},
      {stage1_6[216]}
   );
   gpc1_1 gpc1392 (
      {stage0_6[456]},
      {stage1_6[217]}
   );
   gpc1_1 gpc1393 (
      {stage0_6[457]},
      {stage1_6[218]}
   );
   gpc1_1 gpc1394 (
      {stage0_6[458]},
      {stage1_6[219]}
   );
   gpc1_1 gpc1395 (
      {stage0_6[459]},
      {stage1_6[220]}
   );
   gpc1_1 gpc1396 (
      {stage0_6[460]},
      {stage1_6[221]}
   );
   gpc1_1 gpc1397 (
      {stage0_6[461]},
      {stage1_6[222]}
   );
   gpc1_1 gpc1398 (
      {stage0_6[462]},
      {stage1_6[223]}
   );
   gpc1_1 gpc1399 (
      {stage0_6[463]},
      {stage1_6[224]}
   );
   gpc1_1 gpc1400 (
      {stage0_6[464]},
      {stage1_6[225]}
   );
   gpc1_1 gpc1401 (
      {stage0_6[465]},
      {stage1_6[226]}
   );
   gpc1_1 gpc1402 (
      {stage0_6[466]},
      {stage1_6[227]}
   );
   gpc1_1 gpc1403 (
      {stage0_6[467]},
      {stage1_6[228]}
   );
   gpc1_1 gpc1404 (
      {stage0_6[468]},
      {stage1_6[229]}
   );
   gpc1_1 gpc1405 (
      {stage0_6[469]},
      {stage1_6[230]}
   );
   gpc1_1 gpc1406 (
      {stage0_6[470]},
      {stage1_6[231]}
   );
   gpc1_1 gpc1407 (
      {stage0_6[471]},
      {stage1_6[232]}
   );
   gpc1_1 gpc1408 (
      {stage0_6[472]},
      {stage1_6[233]}
   );
   gpc1_1 gpc1409 (
      {stage0_6[473]},
      {stage1_6[234]}
   );
   gpc1_1 gpc1410 (
      {stage0_6[474]},
      {stage1_6[235]}
   );
   gpc1_1 gpc1411 (
      {stage0_6[475]},
      {stage1_6[236]}
   );
   gpc1_1 gpc1412 (
      {stage0_6[476]},
      {stage1_6[237]}
   );
   gpc1_1 gpc1413 (
      {stage0_6[477]},
      {stage1_6[238]}
   );
   gpc1_1 gpc1414 (
      {stage0_6[478]},
      {stage1_6[239]}
   );
   gpc1_1 gpc1415 (
      {stage0_6[479]},
      {stage1_6[240]}
   );
   gpc1_1 gpc1416 (
      {stage0_6[480]},
      {stage1_6[241]}
   );
   gpc1_1 gpc1417 (
      {stage0_6[481]},
      {stage1_6[242]}
   );
   gpc1_1 gpc1418 (
      {stage0_6[482]},
      {stage1_6[243]}
   );
   gpc1_1 gpc1419 (
      {stage0_6[483]},
      {stage1_6[244]}
   );
   gpc1_1 gpc1420 (
      {stage0_6[484]},
      {stage1_6[245]}
   );
   gpc1_1 gpc1421 (
      {stage0_6[485]},
      {stage1_6[246]}
   );
   gpc1_1 gpc1422 (
      {stage0_7[436]},
      {stage1_7[174]}
   );
   gpc1_1 gpc1423 (
      {stage0_7[437]},
      {stage1_7[175]}
   );
   gpc1_1 gpc1424 (
      {stage0_7[438]},
      {stage1_7[176]}
   );
   gpc1_1 gpc1425 (
      {stage0_7[439]},
      {stage1_7[177]}
   );
   gpc1_1 gpc1426 (
      {stage0_7[440]},
      {stage1_7[178]}
   );
   gpc1_1 gpc1427 (
      {stage0_7[441]},
      {stage1_7[179]}
   );
   gpc1_1 gpc1428 (
      {stage0_7[442]},
      {stage1_7[180]}
   );
   gpc1_1 gpc1429 (
      {stage0_7[443]},
      {stage1_7[181]}
   );
   gpc1_1 gpc1430 (
      {stage0_7[444]},
      {stage1_7[182]}
   );
   gpc1_1 gpc1431 (
      {stage0_7[445]},
      {stage1_7[183]}
   );
   gpc1_1 gpc1432 (
      {stage0_7[446]},
      {stage1_7[184]}
   );
   gpc1_1 gpc1433 (
      {stage0_7[447]},
      {stage1_7[185]}
   );
   gpc1_1 gpc1434 (
      {stage0_7[448]},
      {stage1_7[186]}
   );
   gpc1_1 gpc1435 (
      {stage0_7[449]},
      {stage1_7[187]}
   );
   gpc1_1 gpc1436 (
      {stage0_7[450]},
      {stage1_7[188]}
   );
   gpc1_1 gpc1437 (
      {stage0_7[451]},
      {stage1_7[189]}
   );
   gpc1_1 gpc1438 (
      {stage0_7[452]},
      {stage1_7[190]}
   );
   gpc1_1 gpc1439 (
      {stage0_7[453]},
      {stage1_7[191]}
   );
   gpc1_1 gpc1440 (
      {stage0_7[454]},
      {stage1_7[192]}
   );
   gpc1_1 gpc1441 (
      {stage0_7[455]},
      {stage1_7[193]}
   );
   gpc1_1 gpc1442 (
      {stage0_7[456]},
      {stage1_7[194]}
   );
   gpc1_1 gpc1443 (
      {stage0_7[457]},
      {stage1_7[195]}
   );
   gpc1_1 gpc1444 (
      {stage0_7[458]},
      {stage1_7[196]}
   );
   gpc1_1 gpc1445 (
      {stage0_7[459]},
      {stage1_7[197]}
   );
   gpc1_1 gpc1446 (
      {stage0_7[460]},
      {stage1_7[198]}
   );
   gpc1_1 gpc1447 (
      {stage0_7[461]},
      {stage1_7[199]}
   );
   gpc1_1 gpc1448 (
      {stage0_7[462]},
      {stage1_7[200]}
   );
   gpc1_1 gpc1449 (
      {stage0_7[463]},
      {stage1_7[201]}
   );
   gpc1_1 gpc1450 (
      {stage0_7[464]},
      {stage1_7[202]}
   );
   gpc1_1 gpc1451 (
      {stage0_7[465]},
      {stage1_7[203]}
   );
   gpc1_1 gpc1452 (
      {stage0_7[466]},
      {stage1_7[204]}
   );
   gpc1_1 gpc1453 (
      {stage0_7[467]},
      {stage1_7[205]}
   );
   gpc1_1 gpc1454 (
      {stage0_7[468]},
      {stage1_7[206]}
   );
   gpc1_1 gpc1455 (
      {stage0_7[469]},
      {stage1_7[207]}
   );
   gpc1_1 gpc1456 (
      {stage0_7[470]},
      {stage1_7[208]}
   );
   gpc1_1 gpc1457 (
      {stage0_7[471]},
      {stage1_7[209]}
   );
   gpc1_1 gpc1458 (
      {stage0_7[472]},
      {stage1_7[210]}
   );
   gpc1_1 gpc1459 (
      {stage0_7[473]},
      {stage1_7[211]}
   );
   gpc1_1 gpc1460 (
      {stage0_7[474]},
      {stage1_7[212]}
   );
   gpc1_1 gpc1461 (
      {stage0_7[475]},
      {stage1_7[213]}
   );
   gpc1_1 gpc1462 (
      {stage0_7[476]},
      {stage1_7[214]}
   );
   gpc1_1 gpc1463 (
      {stage0_7[477]},
      {stage1_7[215]}
   );
   gpc1_1 gpc1464 (
      {stage0_7[478]},
      {stage1_7[216]}
   );
   gpc1_1 gpc1465 (
      {stage0_7[479]},
      {stage1_7[217]}
   );
   gpc1_1 gpc1466 (
      {stage0_7[480]},
      {stage1_7[218]}
   );
   gpc1_1 gpc1467 (
      {stage0_7[481]},
      {stage1_7[219]}
   );
   gpc1_1 gpc1468 (
      {stage0_7[482]},
      {stage1_7[220]}
   );
   gpc1_1 gpc1469 (
      {stage0_7[483]},
      {stage1_7[221]}
   );
   gpc1_1 gpc1470 (
      {stage0_7[484]},
      {stage1_7[222]}
   );
   gpc1_1 gpc1471 (
      {stage0_7[485]},
      {stage1_7[223]}
   );
   gpc1_1 gpc1472 (
      {stage0_9[478]},
      {stage1_9[206]}
   );
   gpc1_1 gpc1473 (
      {stage0_9[479]},
      {stage1_9[207]}
   );
   gpc1_1 gpc1474 (
      {stage0_9[480]},
      {stage1_9[208]}
   );
   gpc1_1 gpc1475 (
      {stage0_9[481]},
      {stage1_9[209]}
   );
   gpc1_1 gpc1476 (
      {stage0_9[482]},
      {stage1_9[210]}
   );
   gpc1_1 gpc1477 (
      {stage0_9[483]},
      {stage1_9[211]}
   );
   gpc1_1 gpc1478 (
      {stage0_9[484]},
      {stage1_9[212]}
   );
   gpc1_1 gpc1479 (
      {stage0_9[485]},
      {stage1_9[213]}
   );
   gpc1_1 gpc1480 (
      {stage0_10[475]},
      {stage1_10[177]}
   );
   gpc1_1 gpc1481 (
      {stage0_10[476]},
      {stage1_10[178]}
   );
   gpc1_1 gpc1482 (
      {stage0_10[477]},
      {stage1_10[179]}
   );
   gpc1_1 gpc1483 (
      {stage0_10[478]},
      {stage1_10[180]}
   );
   gpc1_1 gpc1484 (
      {stage0_10[479]},
      {stage1_10[181]}
   );
   gpc1_1 gpc1485 (
      {stage0_10[480]},
      {stage1_10[182]}
   );
   gpc1_1 gpc1486 (
      {stage0_10[481]},
      {stage1_10[183]}
   );
   gpc1_1 gpc1487 (
      {stage0_10[482]},
      {stage1_10[184]}
   );
   gpc1_1 gpc1488 (
      {stage0_10[483]},
      {stage1_10[185]}
   );
   gpc1_1 gpc1489 (
      {stage0_10[484]},
      {stage1_10[186]}
   );
   gpc1_1 gpc1490 (
      {stage0_10[485]},
      {stage1_10[187]}
   );
   gpc1_1 gpc1491 (
      {stage0_11[451]},
      {stage1_11[185]}
   );
   gpc1_1 gpc1492 (
      {stage0_11[452]},
      {stage1_11[186]}
   );
   gpc1_1 gpc1493 (
      {stage0_11[453]},
      {stage1_11[187]}
   );
   gpc1_1 gpc1494 (
      {stage0_11[454]},
      {stage1_11[188]}
   );
   gpc1_1 gpc1495 (
      {stage0_11[455]},
      {stage1_11[189]}
   );
   gpc1_1 gpc1496 (
      {stage0_11[456]},
      {stage1_11[190]}
   );
   gpc1_1 gpc1497 (
      {stage0_11[457]},
      {stage1_11[191]}
   );
   gpc1_1 gpc1498 (
      {stage0_11[458]},
      {stage1_11[192]}
   );
   gpc1_1 gpc1499 (
      {stage0_11[459]},
      {stage1_11[193]}
   );
   gpc1_1 gpc1500 (
      {stage0_11[460]},
      {stage1_11[194]}
   );
   gpc1_1 gpc1501 (
      {stage0_11[461]},
      {stage1_11[195]}
   );
   gpc1_1 gpc1502 (
      {stage0_11[462]},
      {stage1_11[196]}
   );
   gpc1_1 gpc1503 (
      {stage0_11[463]},
      {stage1_11[197]}
   );
   gpc1_1 gpc1504 (
      {stage0_11[464]},
      {stage1_11[198]}
   );
   gpc1_1 gpc1505 (
      {stage0_11[465]},
      {stage1_11[199]}
   );
   gpc1_1 gpc1506 (
      {stage0_11[466]},
      {stage1_11[200]}
   );
   gpc1_1 gpc1507 (
      {stage0_11[467]},
      {stage1_11[201]}
   );
   gpc1_1 gpc1508 (
      {stage0_11[468]},
      {stage1_11[202]}
   );
   gpc1_1 gpc1509 (
      {stage0_11[469]},
      {stage1_11[203]}
   );
   gpc1_1 gpc1510 (
      {stage0_11[470]},
      {stage1_11[204]}
   );
   gpc1_1 gpc1511 (
      {stage0_11[471]},
      {stage1_11[205]}
   );
   gpc1_1 gpc1512 (
      {stage0_11[472]},
      {stage1_11[206]}
   );
   gpc1_1 gpc1513 (
      {stage0_11[473]},
      {stage1_11[207]}
   );
   gpc1_1 gpc1514 (
      {stage0_11[474]},
      {stage1_11[208]}
   );
   gpc1_1 gpc1515 (
      {stage0_11[475]},
      {stage1_11[209]}
   );
   gpc1_1 gpc1516 (
      {stage0_11[476]},
      {stage1_11[210]}
   );
   gpc1_1 gpc1517 (
      {stage0_11[477]},
      {stage1_11[211]}
   );
   gpc1_1 gpc1518 (
      {stage0_11[478]},
      {stage1_11[212]}
   );
   gpc1_1 gpc1519 (
      {stage0_11[479]},
      {stage1_11[213]}
   );
   gpc1_1 gpc1520 (
      {stage0_11[480]},
      {stage1_11[214]}
   );
   gpc1_1 gpc1521 (
      {stage0_11[481]},
      {stage1_11[215]}
   );
   gpc1_1 gpc1522 (
      {stage0_11[482]},
      {stage1_11[216]}
   );
   gpc1_1 gpc1523 (
      {stage0_11[483]},
      {stage1_11[217]}
   );
   gpc1_1 gpc1524 (
      {stage0_11[484]},
      {stage1_11[218]}
   );
   gpc1_1 gpc1525 (
      {stage0_11[485]},
      {stage1_11[219]}
   );
   gpc1_1 gpc1526 (
      {stage0_12[408]},
      {stage1_12[204]}
   );
   gpc1_1 gpc1527 (
      {stage0_12[409]},
      {stage1_12[205]}
   );
   gpc1_1 gpc1528 (
      {stage0_12[410]},
      {stage1_12[206]}
   );
   gpc1_1 gpc1529 (
      {stage0_12[411]},
      {stage1_12[207]}
   );
   gpc1_1 gpc1530 (
      {stage0_12[412]},
      {stage1_12[208]}
   );
   gpc1_1 gpc1531 (
      {stage0_12[413]},
      {stage1_12[209]}
   );
   gpc1_1 gpc1532 (
      {stage0_12[414]},
      {stage1_12[210]}
   );
   gpc1_1 gpc1533 (
      {stage0_12[415]},
      {stage1_12[211]}
   );
   gpc1_1 gpc1534 (
      {stage0_12[416]},
      {stage1_12[212]}
   );
   gpc1_1 gpc1535 (
      {stage0_12[417]},
      {stage1_12[213]}
   );
   gpc1_1 gpc1536 (
      {stage0_12[418]},
      {stage1_12[214]}
   );
   gpc1_1 gpc1537 (
      {stage0_12[419]},
      {stage1_12[215]}
   );
   gpc1_1 gpc1538 (
      {stage0_12[420]},
      {stage1_12[216]}
   );
   gpc1_1 gpc1539 (
      {stage0_12[421]},
      {stage1_12[217]}
   );
   gpc1_1 gpc1540 (
      {stage0_12[422]},
      {stage1_12[218]}
   );
   gpc1_1 gpc1541 (
      {stage0_12[423]},
      {stage1_12[219]}
   );
   gpc1_1 gpc1542 (
      {stage0_12[424]},
      {stage1_12[220]}
   );
   gpc1_1 gpc1543 (
      {stage0_12[425]},
      {stage1_12[221]}
   );
   gpc1_1 gpc1544 (
      {stage0_12[426]},
      {stage1_12[222]}
   );
   gpc1_1 gpc1545 (
      {stage0_12[427]},
      {stage1_12[223]}
   );
   gpc1_1 gpc1546 (
      {stage0_12[428]},
      {stage1_12[224]}
   );
   gpc1_1 gpc1547 (
      {stage0_12[429]},
      {stage1_12[225]}
   );
   gpc1_1 gpc1548 (
      {stage0_12[430]},
      {stage1_12[226]}
   );
   gpc1_1 gpc1549 (
      {stage0_12[431]},
      {stage1_12[227]}
   );
   gpc1_1 gpc1550 (
      {stage0_12[432]},
      {stage1_12[228]}
   );
   gpc1_1 gpc1551 (
      {stage0_12[433]},
      {stage1_12[229]}
   );
   gpc1_1 gpc1552 (
      {stage0_12[434]},
      {stage1_12[230]}
   );
   gpc1_1 gpc1553 (
      {stage0_12[435]},
      {stage1_12[231]}
   );
   gpc1_1 gpc1554 (
      {stage0_12[436]},
      {stage1_12[232]}
   );
   gpc1_1 gpc1555 (
      {stage0_12[437]},
      {stage1_12[233]}
   );
   gpc1_1 gpc1556 (
      {stage0_12[438]},
      {stage1_12[234]}
   );
   gpc1_1 gpc1557 (
      {stage0_12[439]},
      {stage1_12[235]}
   );
   gpc1_1 gpc1558 (
      {stage0_12[440]},
      {stage1_12[236]}
   );
   gpc1_1 gpc1559 (
      {stage0_12[441]},
      {stage1_12[237]}
   );
   gpc1_1 gpc1560 (
      {stage0_12[442]},
      {stage1_12[238]}
   );
   gpc1_1 gpc1561 (
      {stage0_12[443]},
      {stage1_12[239]}
   );
   gpc1_1 gpc1562 (
      {stage0_12[444]},
      {stage1_12[240]}
   );
   gpc1_1 gpc1563 (
      {stage0_12[445]},
      {stage1_12[241]}
   );
   gpc1_1 gpc1564 (
      {stage0_12[446]},
      {stage1_12[242]}
   );
   gpc1_1 gpc1565 (
      {stage0_12[447]},
      {stage1_12[243]}
   );
   gpc1_1 gpc1566 (
      {stage0_12[448]},
      {stage1_12[244]}
   );
   gpc1_1 gpc1567 (
      {stage0_12[449]},
      {stage1_12[245]}
   );
   gpc1_1 gpc1568 (
      {stage0_12[450]},
      {stage1_12[246]}
   );
   gpc1_1 gpc1569 (
      {stage0_12[451]},
      {stage1_12[247]}
   );
   gpc1_1 gpc1570 (
      {stage0_12[452]},
      {stage1_12[248]}
   );
   gpc1_1 gpc1571 (
      {stage0_12[453]},
      {stage1_12[249]}
   );
   gpc1_1 gpc1572 (
      {stage0_12[454]},
      {stage1_12[250]}
   );
   gpc1_1 gpc1573 (
      {stage0_12[455]},
      {stage1_12[251]}
   );
   gpc1_1 gpc1574 (
      {stage0_12[456]},
      {stage1_12[252]}
   );
   gpc1_1 gpc1575 (
      {stage0_12[457]},
      {stage1_12[253]}
   );
   gpc1_1 gpc1576 (
      {stage0_12[458]},
      {stage1_12[254]}
   );
   gpc1_1 gpc1577 (
      {stage0_12[459]},
      {stage1_12[255]}
   );
   gpc1_1 gpc1578 (
      {stage0_12[460]},
      {stage1_12[256]}
   );
   gpc1_1 gpc1579 (
      {stage0_12[461]},
      {stage1_12[257]}
   );
   gpc1_1 gpc1580 (
      {stage0_12[462]},
      {stage1_12[258]}
   );
   gpc1_1 gpc1581 (
      {stage0_12[463]},
      {stage1_12[259]}
   );
   gpc1_1 gpc1582 (
      {stage0_12[464]},
      {stage1_12[260]}
   );
   gpc1_1 gpc1583 (
      {stage0_12[465]},
      {stage1_12[261]}
   );
   gpc1_1 gpc1584 (
      {stage0_12[466]},
      {stage1_12[262]}
   );
   gpc1_1 gpc1585 (
      {stage0_12[467]},
      {stage1_12[263]}
   );
   gpc1_1 gpc1586 (
      {stage0_12[468]},
      {stage1_12[264]}
   );
   gpc1_1 gpc1587 (
      {stage0_12[469]},
      {stage1_12[265]}
   );
   gpc1_1 gpc1588 (
      {stage0_12[470]},
      {stage1_12[266]}
   );
   gpc1_1 gpc1589 (
      {stage0_12[471]},
      {stage1_12[267]}
   );
   gpc1_1 gpc1590 (
      {stage0_12[472]},
      {stage1_12[268]}
   );
   gpc1_1 gpc1591 (
      {stage0_12[473]},
      {stage1_12[269]}
   );
   gpc1_1 gpc1592 (
      {stage0_12[474]},
      {stage1_12[270]}
   );
   gpc1_1 gpc1593 (
      {stage0_12[475]},
      {stage1_12[271]}
   );
   gpc1_1 gpc1594 (
      {stage0_12[476]},
      {stage1_12[272]}
   );
   gpc1_1 gpc1595 (
      {stage0_12[477]},
      {stage1_12[273]}
   );
   gpc1_1 gpc1596 (
      {stage0_12[478]},
      {stage1_12[274]}
   );
   gpc1_1 gpc1597 (
      {stage0_12[479]},
      {stage1_12[275]}
   );
   gpc1_1 gpc1598 (
      {stage0_12[480]},
      {stage1_12[276]}
   );
   gpc1_1 gpc1599 (
      {stage0_12[481]},
      {stage1_12[277]}
   );
   gpc1_1 gpc1600 (
      {stage0_12[482]},
      {stage1_12[278]}
   );
   gpc1_1 gpc1601 (
      {stage0_12[483]},
      {stage1_12[279]}
   );
   gpc1_1 gpc1602 (
      {stage0_12[484]},
      {stage1_12[280]}
   );
   gpc1_1 gpc1603 (
      {stage0_12[485]},
      {stage1_12[281]}
   );
   gpc1_1 gpc1604 (
      {stage0_13[476]},
      {stage1_13[195]}
   );
   gpc1_1 gpc1605 (
      {stage0_13[477]},
      {stage1_13[196]}
   );
   gpc1_1 gpc1606 (
      {stage0_13[478]},
      {stage1_13[197]}
   );
   gpc1_1 gpc1607 (
      {stage0_13[479]},
      {stage1_13[198]}
   );
   gpc1_1 gpc1608 (
      {stage0_13[480]},
      {stage1_13[199]}
   );
   gpc1_1 gpc1609 (
      {stage0_13[481]},
      {stage1_13[200]}
   );
   gpc1_1 gpc1610 (
      {stage0_13[482]},
      {stage1_13[201]}
   );
   gpc1_1 gpc1611 (
      {stage0_13[483]},
      {stage1_13[202]}
   );
   gpc1_1 gpc1612 (
      {stage0_13[484]},
      {stage1_13[203]}
   );
   gpc1_1 gpc1613 (
      {stage0_13[485]},
      {stage1_13[204]}
   );
   gpc1_1 gpc1614 (
      {stage0_14[349]},
      {stage1_14[160]}
   );
   gpc1_1 gpc1615 (
      {stage0_14[350]},
      {stage1_14[161]}
   );
   gpc1_1 gpc1616 (
      {stage0_14[351]},
      {stage1_14[162]}
   );
   gpc1_1 gpc1617 (
      {stage0_14[352]},
      {stage1_14[163]}
   );
   gpc1_1 gpc1618 (
      {stage0_14[353]},
      {stage1_14[164]}
   );
   gpc1_1 gpc1619 (
      {stage0_14[354]},
      {stage1_14[165]}
   );
   gpc1_1 gpc1620 (
      {stage0_14[355]},
      {stage1_14[166]}
   );
   gpc1_1 gpc1621 (
      {stage0_14[356]},
      {stage1_14[167]}
   );
   gpc1_1 gpc1622 (
      {stage0_14[357]},
      {stage1_14[168]}
   );
   gpc1_1 gpc1623 (
      {stage0_14[358]},
      {stage1_14[169]}
   );
   gpc1_1 gpc1624 (
      {stage0_14[359]},
      {stage1_14[170]}
   );
   gpc1_1 gpc1625 (
      {stage0_14[360]},
      {stage1_14[171]}
   );
   gpc1_1 gpc1626 (
      {stage0_14[361]},
      {stage1_14[172]}
   );
   gpc1_1 gpc1627 (
      {stage0_14[362]},
      {stage1_14[173]}
   );
   gpc1_1 gpc1628 (
      {stage0_14[363]},
      {stage1_14[174]}
   );
   gpc1_1 gpc1629 (
      {stage0_14[364]},
      {stage1_14[175]}
   );
   gpc1_1 gpc1630 (
      {stage0_14[365]},
      {stage1_14[176]}
   );
   gpc1_1 gpc1631 (
      {stage0_14[366]},
      {stage1_14[177]}
   );
   gpc1_1 gpc1632 (
      {stage0_14[367]},
      {stage1_14[178]}
   );
   gpc1_1 gpc1633 (
      {stage0_14[368]},
      {stage1_14[179]}
   );
   gpc1_1 gpc1634 (
      {stage0_14[369]},
      {stage1_14[180]}
   );
   gpc1_1 gpc1635 (
      {stage0_14[370]},
      {stage1_14[181]}
   );
   gpc1_1 gpc1636 (
      {stage0_14[371]},
      {stage1_14[182]}
   );
   gpc1_1 gpc1637 (
      {stage0_14[372]},
      {stage1_14[183]}
   );
   gpc1_1 gpc1638 (
      {stage0_14[373]},
      {stage1_14[184]}
   );
   gpc1_1 gpc1639 (
      {stage0_14[374]},
      {stage1_14[185]}
   );
   gpc1_1 gpc1640 (
      {stage0_14[375]},
      {stage1_14[186]}
   );
   gpc1_1 gpc1641 (
      {stage0_14[376]},
      {stage1_14[187]}
   );
   gpc1_1 gpc1642 (
      {stage0_14[377]},
      {stage1_14[188]}
   );
   gpc1_1 gpc1643 (
      {stage0_14[378]},
      {stage1_14[189]}
   );
   gpc1_1 gpc1644 (
      {stage0_14[379]},
      {stage1_14[190]}
   );
   gpc1_1 gpc1645 (
      {stage0_14[380]},
      {stage1_14[191]}
   );
   gpc1_1 gpc1646 (
      {stage0_14[381]},
      {stage1_14[192]}
   );
   gpc1_1 gpc1647 (
      {stage0_14[382]},
      {stage1_14[193]}
   );
   gpc1_1 gpc1648 (
      {stage0_14[383]},
      {stage1_14[194]}
   );
   gpc1_1 gpc1649 (
      {stage0_14[384]},
      {stage1_14[195]}
   );
   gpc1_1 gpc1650 (
      {stage0_14[385]},
      {stage1_14[196]}
   );
   gpc1_1 gpc1651 (
      {stage0_14[386]},
      {stage1_14[197]}
   );
   gpc1_1 gpc1652 (
      {stage0_14[387]},
      {stage1_14[198]}
   );
   gpc1_1 gpc1653 (
      {stage0_14[388]},
      {stage1_14[199]}
   );
   gpc1_1 gpc1654 (
      {stage0_14[389]},
      {stage1_14[200]}
   );
   gpc1_1 gpc1655 (
      {stage0_14[390]},
      {stage1_14[201]}
   );
   gpc1_1 gpc1656 (
      {stage0_14[391]},
      {stage1_14[202]}
   );
   gpc1_1 gpc1657 (
      {stage0_14[392]},
      {stage1_14[203]}
   );
   gpc1_1 gpc1658 (
      {stage0_14[393]},
      {stage1_14[204]}
   );
   gpc1_1 gpc1659 (
      {stage0_14[394]},
      {stage1_14[205]}
   );
   gpc1_1 gpc1660 (
      {stage0_14[395]},
      {stage1_14[206]}
   );
   gpc1_1 gpc1661 (
      {stage0_14[396]},
      {stage1_14[207]}
   );
   gpc1_1 gpc1662 (
      {stage0_14[397]},
      {stage1_14[208]}
   );
   gpc1_1 gpc1663 (
      {stage0_14[398]},
      {stage1_14[209]}
   );
   gpc1_1 gpc1664 (
      {stage0_14[399]},
      {stage1_14[210]}
   );
   gpc1_1 gpc1665 (
      {stage0_14[400]},
      {stage1_14[211]}
   );
   gpc1_1 gpc1666 (
      {stage0_14[401]},
      {stage1_14[212]}
   );
   gpc1_1 gpc1667 (
      {stage0_14[402]},
      {stage1_14[213]}
   );
   gpc1_1 gpc1668 (
      {stage0_14[403]},
      {stage1_14[214]}
   );
   gpc1_1 gpc1669 (
      {stage0_14[404]},
      {stage1_14[215]}
   );
   gpc1_1 gpc1670 (
      {stage0_14[405]},
      {stage1_14[216]}
   );
   gpc1_1 gpc1671 (
      {stage0_14[406]},
      {stage1_14[217]}
   );
   gpc1_1 gpc1672 (
      {stage0_14[407]},
      {stage1_14[218]}
   );
   gpc1_1 gpc1673 (
      {stage0_14[408]},
      {stage1_14[219]}
   );
   gpc1_1 gpc1674 (
      {stage0_14[409]},
      {stage1_14[220]}
   );
   gpc1_1 gpc1675 (
      {stage0_14[410]},
      {stage1_14[221]}
   );
   gpc1_1 gpc1676 (
      {stage0_14[411]},
      {stage1_14[222]}
   );
   gpc1_1 gpc1677 (
      {stage0_14[412]},
      {stage1_14[223]}
   );
   gpc1_1 gpc1678 (
      {stage0_14[413]},
      {stage1_14[224]}
   );
   gpc1_1 gpc1679 (
      {stage0_14[414]},
      {stage1_14[225]}
   );
   gpc1_1 gpc1680 (
      {stage0_14[415]},
      {stage1_14[226]}
   );
   gpc1_1 gpc1681 (
      {stage0_14[416]},
      {stage1_14[227]}
   );
   gpc1_1 gpc1682 (
      {stage0_14[417]},
      {stage1_14[228]}
   );
   gpc1_1 gpc1683 (
      {stage0_14[418]},
      {stage1_14[229]}
   );
   gpc1_1 gpc1684 (
      {stage0_14[419]},
      {stage1_14[230]}
   );
   gpc1_1 gpc1685 (
      {stage0_14[420]},
      {stage1_14[231]}
   );
   gpc1_1 gpc1686 (
      {stage0_14[421]},
      {stage1_14[232]}
   );
   gpc1_1 gpc1687 (
      {stage0_14[422]},
      {stage1_14[233]}
   );
   gpc1_1 gpc1688 (
      {stage0_14[423]},
      {stage1_14[234]}
   );
   gpc1_1 gpc1689 (
      {stage0_14[424]},
      {stage1_14[235]}
   );
   gpc1_1 gpc1690 (
      {stage0_14[425]},
      {stage1_14[236]}
   );
   gpc1_1 gpc1691 (
      {stage0_14[426]},
      {stage1_14[237]}
   );
   gpc1_1 gpc1692 (
      {stage0_14[427]},
      {stage1_14[238]}
   );
   gpc1_1 gpc1693 (
      {stage0_14[428]},
      {stage1_14[239]}
   );
   gpc1_1 gpc1694 (
      {stage0_14[429]},
      {stage1_14[240]}
   );
   gpc1_1 gpc1695 (
      {stage0_14[430]},
      {stage1_14[241]}
   );
   gpc1_1 gpc1696 (
      {stage0_14[431]},
      {stage1_14[242]}
   );
   gpc1_1 gpc1697 (
      {stage0_14[432]},
      {stage1_14[243]}
   );
   gpc1_1 gpc1698 (
      {stage0_14[433]},
      {stage1_14[244]}
   );
   gpc1_1 gpc1699 (
      {stage0_14[434]},
      {stage1_14[245]}
   );
   gpc1_1 gpc1700 (
      {stage0_14[435]},
      {stage1_14[246]}
   );
   gpc1_1 gpc1701 (
      {stage0_14[436]},
      {stage1_14[247]}
   );
   gpc1_1 gpc1702 (
      {stage0_14[437]},
      {stage1_14[248]}
   );
   gpc1_1 gpc1703 (
      {stage0_14[438]},
      {stage1_14[249]}
   );
   gpc1_1 gpc1704 (
      {stage0_14[439]},
      {stage1_14[250]}
   );
   gpc1_1 gpc1705 (
      {stage0_14[440]},
      {stage1_14[251]}
   );
   gpc1_1 gpc1706 (
      {stage0_14[441]},
      {stage1_14[252]}
   );
   gpc1_1 gpc1707 (
      {stage0_14[442]},
      {stage1_14[253]}
   );
   gpc1_1 gpc1708 (
      {stage0_14[443]},
      {stage1_14[254]}
   );
   gpc1_1 gpc1709 (
      {stage0_14[444]},
      {stage1_14[255]}
   );
   gpc1_1 gpc1710 (
      {stage0_14[445]},
      {stage1_14[256]}
   );
   gpc1_1 gpc1711 (
      {stage0_14[446]},
      {stage1_14[257]}
   );
   gpc1_1 gpc1712 (
      {stage0_14[447]},
      {stage1_14[258]}
   );
   gpc1_1 gpc1713 (
      {stage0_14[448]},
      {stage1_14[259]}
   );
   gpc1_1 gpc1714 (
      {stage0_14[449]},
      {stage1_14[260]}
   );
   gpc1_1 gpc1715 (
      {stage0_14[450]},
      {stage1_14[261]}
   );
   gpc1_1 gpc1716 (
      {stage0_14[451]},
      {stage1_14[262]}
   );
   gpc1_1 gpc1717 (
      {stage0_14[452]},
      {stage1_14[263]}
   );
   gpc1_1 gpc1718 (
      {stage0_14[453]},
      {stage1_14[264]}
   );
   gpc1_1 gpc1719 (
      {stage0_14[454]},
      {stage1_14[265]}
   );
   gpc1_1 gpc1720 (
      {stage0_14[455]},
      {stage1_14[266]}
   );
   gpc1_1 gpc1721 (
      {stage0_14[456]},
      {stage1_14[267]}
   );
   gpc1_1 gpc1722 (
      {stage0_14[457]},
      {stage1_14[268]}
   );
   gpc1_1 gpc1723 (
      {stage0_14[458]},
      {stage1_14[269]}
   );
   gpc1_1 gpc1724 (
      {stage0_14[459]},
      {stage1_14[270]}
   );
   gpc1_1 gpc1725 (
      {stage0_14[460]},
      {stage1_14[271]}
   );
   gpc1_1 gpc1726 (
      {stage0_14[461]},
      {stage1_14[272]}
   );
   gpc1_1 gpc1727 (
      {stage0_14[462]},
      {stage1_14[273]}
   );
   gpc1_1 gpc1728 (
      {stage0_14[463]},
      {stage1_14[274]}
   );
   gpc1_1 gpc1729 (
      {stage0_14[464]},
      {stage1_14[275]}
   );
   gpc1_1 gpc1730 (
      {stage0_14[465]},
      {stage1_14[276]}
   );
   gpc1_1 gpc1731 (
      {stage0_14[466]},
      {stage1_14[277]}
   );
   gpc1_1 gpc1732 (
      {stage0_14[467]},
      {stage1_14[278]}
   );
   gpc1_1 gpc1733 (
      {stage0_14[468]},
      {stage1_14[279]}
   );
   gpc1_1 gpc1734 (
      {stage0_14[469]},
      {stage1_14[280]}
   );
   gpc1_1 gpc1735 (
      {stage0_14[470]},
      {stage1_14[281]}
   );
   gpc1_1 gpc1736 (
      {stage0_14[471]},
      {stage1_14[282]}
   );
   gpc1_1 gpc1737 (
      {stage0_14[472]},
      {stage1_14[283]}
   );
   gpc1_1 gpc1738 (
      {stage0_14[473]},
      {stage1_14[284]}
   );
   gpc1_1 gpc1739 (
      {stage0_14[474]},
      {stage1_14[285]}
   );
   gpc1_1 gpc1740 (
      {stage0_14[475]},
      {stage1_14[286]}
   );
   gpc1_1 gpc1741 (
      {stage0_14[476]},
      {stage1_14[287]}
   );
   gpc1_1 gpc1742 (
      {stage0_14[477]},
      {stage1_14[288]}
   );
   gpc1_1 gpc1743 (
      {stage0_14[478]},
      {stage1_14[289]}
   );
   gpc1_1 gpc1744 (
      {stage0_14[479]},
      {stage1_14[290]}
   );
   gpc1_1 gpc1745 (
      {stage0_14[480]},
      {stage1_14[291]}
   );
   gpc1_1 gpc1746 (
      {stage0_14[481]},
      {stage1_14[292]}
   );
   gpc1_1 gpc1747 (
      {stage0_14[482]},
      {stage1_14[293]}
   );
   gpc1_1 gpc1748 (
      {stage0_14[483]},
      {stage1_14[294]}
   );
   gpc1_1 gpc1749 (
      {stage0_14[484]},
      {stage1_14[295]}
   );
   gpc1_1 gpc1750 (
      {stage0_14[485]},
      {stage1_14[296]}
   );
   gpc1_1 gpc1751 (
      {stage0_15[480]},
      {stage1_15[166]}
   );
   gpc1_1 gpc1752 (
      {stage0_15[481]},
      {stage1_15[167]}
   );
   gpc1_1 gpc1753 (
      {stage0_15[482]},
      {stage1_15[168]}
   );
   gpc1_1 gpc1754 (
      {stage0_15[483]},
      {stage1_15[169]}
   );
   gpc1_1 gpc1755 (
      {stage0_15[484]},
      {stage1_15[170]}
   );
   gpc1_1 gpc1756 (
      {stage0_15[485]},
      {stage1_15[171]}
   );
   gpc1_1 gpc1757 (
      {stage0_16[411]},
      {stage1_16[190]}
   );
   gpc1_1 gpc1758 (
      {stage0_16[412]},
      {stage1_16[191]}
   );
   gpc1_1 gpc1759 (
      {stage0_16[413]},
      {stage1_16[192]}
   );
   gpc1_1 gpc1760 (
      {stage0_16[414]},
      {stage1_16[193]}
   );
   gpc1_1 gpc1761 (
      {stage0_16[415]},
      {stage1_16[194]}
   );
   gpc1_1 gpc1762 (
      {stage0_16[416]},
      {stage1_16[195]}
   );
   gpc1_1 gpc1763 (
      {stage0_16[417]},
      {stage1_16[196]}
   );
   gpc1_1 gpc1764 (
      {stage0_16[418]},
      {stage1_16[197]}
   );
   gpc1_1 gpc1765 (
      {stage0_16[419]},
      {stage1_16[198]}
   );
   gpc1_1 gpc1766 (
      {stage0_16[420]},
      {stage1_16[199]}
   );
   gpc1_1 gpc1767 (
      {stage0_16[421]},
      {stage1_16[200]}
   );
   gpc1_1 gpc1768 (
      {stage0_16[422]},
      {stage1_16[201]}
   );
   gpc1_1 gpc1769 (
      {stage0_16[423]},
      {stage1_16[202]}
   );
   gpc1_1 gpc1770 (
      {stage0_16[424]},
      {stage1_16[203]}
   );
   gpc1_1 gpc1771 (
      {stage0_16[425]},
      {stage1_16[204]}
   );
   gpc1_1 gpc1772 (
      {stage0_16[426]},
      {stage1_16[205]}
   );
   gpc1_1 gpc1773 (
      {stage0_16[427]},
      {stage1_16[206]}
   );
   gpc1_1 gpc1774 (
      {stage0_16[428]},
      {stage1_16[207]}
   );
   gpc1_1 gpc1775 (
      {stage0_16[429]},
      {stage1_16[208]}
   );
   gpc1_1 gpc1776 (
      {stage0_16[430]},
      {stage1_16[209]}
   );
   gpc1_1 gpc1777 (
      {stage0_16[431]},
      {stage1_16[210]}
   );
   gpc1_1 gpc1778 (
      {stage0_16[432]},
      {stage1_16[211]}
   );
   gpc1_1 gpc1779 (
      {stage0_16[433]},
      {stage1_16[212]}
   );
   gpc1_1 gpc1780 (
      {stage0_16[434]},
      {stage1_16[213]}
   );
   gpc1_1 gpc1781 (
      {stage0_16[435]},
      {stage1_16[214]}
   );
   gpc1_1 gpc1782 (
      {stage0_16[436]},
      {stage1_16[215]}
   );
   gpc1_1 gpc1783 (
      {stage0_16[437]},
      {stage1_16[216]}
   );
   gpc1_1 gpc1784 (
      {stage0_16[438]},
      {stage1_16[217]}
   );
   gpc1_1 gpc1785 (
      {stage0_16[439]},
      {stage1_16[218]}
   );
   gpc1_1 gpc1786 (
      {stage0_16[440]},
      {stage1_16[219]}
   );
   gpc1_1 gpc1787 (
      {stage0_16[441]},
      {stage1_16[220]}
   );
   gpc1_1 gpc1788 (
      {stage0_16[442]},
      {stage1_16[221]}
   );
   gpc1_1 gpc1789 (
      {stage0_16[443]},
      {stage1_16[222]}
   );
   gpc1_1 gpc1790 (
      {stage0_16[444]},
      {stage1_16[223]}
   );
   gpc1_1 gpc1791 (
      {stage0_16[445]},
      {stage1_16[224]}
   );
   gpc1_1 gpc1792 (
      {stage0_16[446]},
      {stage1_16[225]}
   );
   gpc1_1 gpc1793 (
      {stage0_16[447]},
      {stage1_16[226]}
   );
   gpc1_1 gpc1794 (
      {stage0_16[448]},
      {stage1_16[227]}
   );
   gpc1_1 gpc1795 (
      {stage0_16[449]},
      {stage1_16[228]}
   );
   gpc1_1 gpc1796 (
      {stage0_16[450]},
      {stage1_16[229]}
   );
   gpc1_1 gpc1797 (
      {stage0_16[451]},
      {stage1_16[230]}
   );
   gpc1_1 gpc1798 (
      {stage0_16[452]},
      {stage1_16[231]}
   );
   gpc1_1 gpc1799 (
      {stage0_16[453]},
      {stage1_16[232]}
   );
   gpc1_1 gpc1800 (
      {stage0_16[454]},
      {stage1_16[233]}
   );
   gpc1_1 gpc1801 (
      {stage0_16[455]},
      {stage1_16[234]}
   );
   gpc1_1 gpc1802 (
      {stage0_16[456]},
      {stage1_16[235]}
   );
   gpc1_1 gpc1803 (
      {stage0_16[457]},
      {stage1_16[236]}
   );
   gpc1_1 gpc1804 (
      {stage0_16[458]},
      {stage1_16[237]}
   );
   gpc1_1 gpc1805 (
      {stage0_16[459]},
      {stage1_16[238]}
   );
   gpc1_1 gpc1806 (
      {stage0_16[460]},
      {stage1_16[239]}
   );
   gpc1_1 gpc1807 (
      {stage0_16[461]},
      {stage1_16[240]}
   );
   gpc1_1 gpc1808 (
      {stage0_16[462]},
      {stage1_16[241]}
   );
   gpc1_1 gpc1809 (
      {stage0_16[463]},
      {stage1_16[242]}
   );
   gpc1_1 gpc1810 (
      {stage0_16[464]},
      {stage1_16[243]}
   );
   gpc1_1 gpc1811 (
      {stage0_16[465]},
      {stage1_16[244]}
   );
   gpc1_1 gpc1812 (
      {stage0_16[466]},
      {stage1_16[245]}
   );
   gpc1_1 gpc1813 (
      {stage0_16[467]},
      {stage1_16[246]}
   );
   gpc1_1 gpc1814 (
      {stage0_16[468]},
      {stage1_16[247]}
   );
   gpc1_1 gpc1815 (
      {stage0_16[469]},
      {stage1_16[248]}
   );
   gpc1_1 gpc1816 (
      {stage0_16[470]},
      {stage1_16[249]}
   );
   gpc1_1 gpc1817 (
      {stage0_16[471]},
      {stage1_16[250]}
   );
   gpc1_1 gpc1818 (
      {stage0_16[472]},
      {stage1_16[251]}
   );
   gpc1_1 gpc1819 (
      {stage0_16[473]},
      {stage1_16[252]}
   );
   gpc1_1 gpc1820 (
      {stage0_16[474]},
      {stage1_16[253]}
   );
   gpc1_1 gpc1821 (
      {stage0_16[475]},
      {stage1_16[254]}
   );
   gpc1_1 gpc1822 (
      {stage0_16[476]},
      {stage1_16[255]}
   );
   gpc1_1 gpc1823 (
      {stage0_16[477]},
      {stage1_16[256]}
   );
   gpc1_1 gpc1824 (
      {stage0_16[478]},
      {stage1_16[257]}
   );
   gpc1_1 gpc1825 (
      {stage0_16[479]},
      {stage1_16[258]}
   );
   gpc1_1 gpc1826 (
      {stage0_16[480]},
      {stage1_16[259]}
   );
   gpc1_1 gpc1827 (
      {stage0_16[481]},
      {stage1_16[260]}
   );
   gpc1_1 gpc1828 (
      {stage0_16[482]},
      {stage1_16[261]}
   );
   gpc1_1 gpc1829 (
      {stage0_16[483]},
      {stage1_16[262]}
   );
   gpc1_1 gpc1830 (
      {stage0_16[484]},
      {stage1_16[263]}
   );
   gpc1_1 gpc1831 (
      {stage0_16[485]},
      {stage1_16[264]}
   );
   gpc1_1 gpc1832 (
      {stage0_17[402]},
      {stage1_17[187]}
   );
   gpc1_1 gpc1833 (
      {stage0_17[403]},
      {stage1_17[188]}
   );
   gpc1_1 gpc1834 (
      {stage0_17[404]},
      {stage1_17[189]}
   );
   gpc1_1 gpc1835 (
      {stage0_17[405]},
      {stage1_17[190]}
   );
   gpc1_1 gpc1836 (
      {stage0_17[406]},
      {stage1_17[191]}
   );
   gpc1_1 gpc1837 (
      {stage0_17[407]},
      {stage1_17[192]}
   );
   gpc1_1 gpc1838 (
      {stage0_17[408]},
      {stage1_17[193]}
   );
   gpc1_1 gpc1839 (
      {stage0_17[409]},
      {stage1_17[194]}
   );
   gpc1_1 gpc1840 (
      {stage0_17[410]},
      {stage1_17[195]}
   );
   gpc1_1 gpc1841 (
      {stage0_17[411]},
      {stage1_17[196]}
   );
   gpc1_1 gpc1842 (
      {stage0_17[412]},
      {stage1_17[197]}
   );
   gpc1_1 gpc1843 (
      {stage0_17[413]},
      {stage1_17[198]}
   );
   gpc1_1 gpc1844 (
      {stage0_17[414]},
      {stage1_17[199]}
   );
   gpc1_1 gpc1845 (
      {stage0_17[415]},
      {stage1_17[200]}
   );
   gpc1_1 gpc1846 (
      {stage0_17[416]},
      {stage1_17[201]}
   );
   gpc1_1 gpc1847 (
      {stage0_17[417]},
      {stage1_17[202]}
   );
   gpc1_1 gpc1848 (
      {stage0_17[418]},
      {stage1_17[203]}
   );
   gpc1_1 gpc1849 (
      {stage0_17[419]},
      {stage1_17[204]}
   );
   gpc1_1 gpc1850 (
      {stage0_17[420]},
      {stage1_17[205]}
   );
   gpc1_1 gpc1851 (
      {stage0_17[421]},
      {stage1_17[206]}
   );
   gpc1_1 gpc1852 (
      {stage0_17[422]},
      {stage1_17[207]}
   );
   gpc1_1 gpc1853 (
      {stage0_17[423]},
      {stage1_17[208]}
   );
   gpc1_1 gpc1854 (
      {stage0_17[424]},
      {stage1_17[209]}
   );
   gpc1_1 gpc1855 (
      {stage0_17[425]},
      {stage1_17[210]}
   );
   gpc1_1 gpc1856 (
      {stage0_17[426]},
      {stage1_17[211]}
   );
   gpc1_1 gpc1857 (
      {stage0_17[427]},
      {stage1_17[212]}
   );
   gpc1_1 gpc1858 (
      {stage0_17[428]},
      {stage1_17[213]}
   );
   gpc1_1 gpc1859 (
      {stage0_17[429]},
      {stage1_17[214]}
   );
   gpc1_1 gpc1860 (
      {stage0_17[430]},
      {stage1_17[215]}
   );
   gpc1_1 gpc1861 (
      {stage0_17[431]},
      {stage1_17[216]}
   );
   gpc1_1 gpc1862 (
      {stage0_17[432]},
      {stage1_17[217]}
   );
   gpc1_1 gpc1863 (
      {stage0_17[433]},
      {stage1_17[218]}
   );
   gpc1_1 gpc1864 (
      {stage0_17[434]},
      {stage1_17[219]}
   );
   gpc1_1 gpc1865 (
      {stage0_17[435]},
      {stage1_17[220]}
   );
   gpc1_1 gpc1866 (
      {stage0_17[436]},
      {stage1_17[221]}
   );
   gpc1_1 gpc1867 (
      {stage0_17[437]},
      {stage1_17[222]}
   );
   gpc1_1 gpc1868 (
      {stage0_17[438]},
      {stage1_17[223]}
   );
   gpc1_1 gpc1869 (
      {stage0_17[439]},
      {stage1_17[224]}
   );
   gpc1_1 gpc1870 (
      {stage0_17[440]},
      {stage1_17[225]}
   );
   gpc1_1 gpc1871 (
      {stage0_17[441]},
      {stage1_17[226]}
   );
   gpc1_1 gpc1872 (
      {stage0_17[442]},
      {stage1_17[227]}
   );
   gpc1_1 gpc1873 (
      {stage0_17[443]},
      {stage1_17[228]}
   );
   gpc1_1 gpc1874 (
      {stage0_17[444]},
      {stage1_17[229]}
   );
   gpc1_1 gpc1875 (
      {stage0_17[445]},
      {stage1_17[230]}
   );
   gpc1_1 gpc1876 (
      {stage0_17[446]},
      {stage1_17[231]}
   );
   gpc1_1 gpc1877 (
      {stage0_17[447]},
      {stage1_17[232]}
   );
   gpc1_1 gpc1878 (
      {stage0_17[448]},
      {stage1_17[233]}
   );
   gpc1_1 gpc1879 (
      {stage0_17[449]},
      {stage1_17[234]}
   );
   gpc1_1 gpc1880 (
      {stage0_17[450]},
      {stage1_17[235]}
   );
   gpc1_1 gpc1881 (
      {stage0_17[451]},
      {stage1_17[236]}
   );
   gpc1_1 gpc1882 (
      {stage0_17[452]},
      {stage1_17[237]}
   );
   gpc1_1 gpc1883 (
      {stage0_17[453]},
      {stage1_17[238]}
   );
   gpc1_1 gpc1884 (
      {stage0_17[454]},
      {stage1_17[239]}
   );
   gpc1_1 gpc1885 (
      {stage0_17[455]},
      {stage1_17[240]}
   );
   gpc1_1 gpc1886 (
      {stage0_17[456]},
      {stage1_17[241]}
   );
   gpc1_1 gpc1887 (
      {stage0_17[457]},
      {stage1_17[242]}
   );
   gpc1_1 gpc1888 (
      {stage0_17[458]},
      {stage1_17[243]}
   );
   gpc1_1 gpc1889 (
      {stage0_17[459]},
      {stage1_17[244]}
   );
   gpc1_1 gpc1890 (
      {stage0_17[460]},
      {stage1_17[245]}
   );
   gpc1_1 gpc1891 (
      {stage0_17[461]},
      {stage1_17[246]}
   );
   gpc1_1 gpc1892 (
      {stage0_17[462]},
      {stage1_17[247]}
   );
   gpc1_1 gpc1893 (
      {stage0_17[463]},
      {stage1_17[248]}
   );
   gpc1_1 gpc1894 (
      {stage0_17[464]},
      {stage1_17[249]}
   );
   gpc1_1 gpc1895 (
      {stage0_17[465]},
      {stage1_17[250]}
   );
   gpc1_1 gpc1896 (
      {stage0_17[466]},
      {stage1_17[251]}
   );
   gpc1_1 gpc1897 (
      {stage0_17[467]},
      {stage1_17[252]}
   );
   gpc1_1 gpc1898 (
      {stage0_17[468]},
      {stage1_17[253]}
   );
   gpc1_1 gpc1899 (
      {stage0_17[469]},
      {stage1_17[254]}
   );
   gpc1_1 gpc1900 (
      {stage0_17[470]},
      {stage1_17[255]}
   );
   gpc1_1 gpc1901 (
      {stage0_17[471]},
      {stage1_17[256]}
   );
   gpc1_1 gpc1902 (
      {stage0_17[472]},
      {stage1_17[257]}
   );
   gpc1_1 gpc1903 (
      {stage0_17[473]},
      {stage1_17[258]}
   );
   gpc1_1 gpc1904 (
      {stage0_17[474]},
      {stage1_17[259]}
   );
   gpc1_1 gpc1905 (
      {stage0_17[475]},
      {stage1_17[260]}
   );
   gpc1_1 gpc1906 (
      {stage0_17[476]},
      {stage1_17[261]}
   );
   gpc1_1 gpc1907 (
      {stage0_17[477]},
      {stage1_17[262]}
   );
   gpc1_1 gpc1908 (
      {stage0_17[478]},
      {stage1_17[263]}
   );
   gpc1_1 gpc1909 (
      {stage0_17[479]},
      {stage1_17[264]}
   );
   gpc1_1 gpc1910 (
      {stage0_17[480]},
      {stage1_17[265]}
   );
   gpc1_1 gpc1911 (
      {stage0_17[481]},
      {stage1_17[266]}
   );
   gpc1_1 gpc1912 (
      {stage0_17[482]},
      {stage1_17[267]}
   );
   gpc1_1 gpc1913 (
      {stage0_17[483]},
      {stage1_17[268]}
   );
   gpc1_1 gpc1914 (
      {stage0_17[484]},
      {stage1_17[269]}
   );
   gpc1_1 gpc1915 (
      {stage0_17[485]},
      {stage1_17[270]}
   );
   gpc1_1 gpc1916 (
      {stage0_18[447]},
      {stage1_18[162]}
   );
   gpc1_1 gpc1917 (
      {stage0_18[448]},
      {stage1_18[163]}
   );
   gpc1_1 gpc1918 (
      {stage0_18[449]},
      {stage1_18[164]}
   );
   gpc1_1 gpc1919 (
      {stage0_18[450]},
      {stage1_18[165]}
   );
   gpc1_1 gpc1920 (
      {stage0_18[451]},
      {stage1_18[166]}
   );
   gpc1_1 gpc1921 (
      {stage0_18[452]},
      {stage1_18[167]}
   );
   gpc1_1 gpc1922 (
      {stage0_18[453]},
      {stage1_18[168]}
   );
   gpc1_1 gpc1923 (
      {stage0_18[454]},
      {stage1_18[169]}
   );
   gpc1_1 gpc1924 (
      {stage0_18[455]},
      {stage1_18[170]}
   );
   gpc1_1 gpc1925 (
      {stage0_18[456]},
      {stage1_18[171]}
   );
   gpc1_1 gpc1926 (
      {stage0_18[457]},
      {stage1_18[172]}
   );
   gpc1_1 gpc1927 (
      {stage0_18[458]},
      {stage1_18[173]}
   );
   gpc1_1 gpc1928 (
      {stage0_18[459]},
      {stage1_18[174]}
   );
   gpc1_1 gpc1929 (
      {stage0_18[460]},
      {stage1_18[175]}
   );
   gpc1_1 gpc1930 (
      {stage0_18[461]},
      {stage1_18[176]}
   );
   gpc1_1 gpc1931 (
      {stage0_18[462]},
      {stage1_18[177]}
   );
   gpc1_1 gpc1932 (
      {stage0_18[463]},
      {stage1_18[178]}
   );
   gpc1_1 gpc1933 (
      {stage0_18[464]},
      {stage1_18[179]}
   );
   gpc1_1 gpc1934 (
      {stage0_18[465]},
      {stage1_18[180]}
   );
   gpc1_1 gpc1935 (
      {stage0_18[466]},
      {stage1_18[181]}
   );
   gpc1_1 gpc1936 (
      {stage0_18[467]},
      {stage1_18[182]}
   );
   gpc1_1 gpc1937 (
      {stage0_18[468]},
      {stage1_18[183]}
   );
   gpc1_1 gpc1938 (
      {stage0_18[469]},
      {stage1_18[184]}
   );
   gpc1_1 gpc1939 (
      {stage0_18[470]},
      {stage1_18[185]}
   );
   gpc1_1 gpc1940 (
      {stage0_18[471]},
      {stage1_18[186]}
   );
   gpc1_1 gpc1941 (
      {stage0_18[472]},
      {stage1_18[187]}
   );
   gpc1_1 gpc1942 (
      {stage0_18[473]},
      {stage1_18[188]}
   );
   gpc1_1 gpc1943 (
      {stage0_18[474]},
      {stage1_18[189]}
   );
   gpc1_1 gpc1944 (
      {stage0_18[475]},
      {stage1_18[190]}
   );
   gpc1_1 gpc1945 (
      {stage0_18[476]},
      {stage1_18[191]}
   );
   gpc1_1 gpc1946 (
      {stage0_18[477]},
      {stage1_18[192]}
   );
   gpc1_1 gpc1947 (
      {stage0_18[478]},
      {stage1_18[193]}
   );
   gpc1_1 gpc1948 (
      {stage0_18[479]},
      {stage1_18[194]}
   );
   gpc1_1 gpc1949 (
      {stage0_18[480]},
      {stage1_18[195]}
   );
   gpc1_1 gpc1950 (
      {stage0_18[481]},
      {stage1_18[196]}
   );
   gpc1_1 gpc1951 (
      {stage0_18[482]},
      {stage1_18[197]}
   );
   gpc1_1 gpc1952 (
      {stage0_18[483]},
      {stage1_18[198]}
   );
   gpc1_1 gpc1953 (
      {stage0_18[484]},
      {stage1_18[199]}
   );
   gpc1_1 gpc1954 (
      {stage0_18[485]},
      {stage1_18[200]}
   );
   gpc1_1 gpc1955 (
      {stage0_19[347]},
      {stage1_19[161]}
   );
   gpc1_1 gpc1956 (
      {stage0_19[348]},
      {stage1_19[162]}
   );
   gpc1_1 gpc1957 (
      {stage0_19[349]},
      {stage1_19[163]}
   );
   gpc1_1 gpc1958 (
      {stage0_19[350]},
      {stage1_19[164]}
   );
   gpc1_1 gpc1959 (
      {stage0_19[351]},
      {stage1_19[165]}
   );
   gpc1_1 gpc1960 (
      {stage0_19[352]},
      {stage1_19[166]}
   );
   gpc1_1 gpc1961 (
      {stage0_19[353]},
      {stage1_19[167]}
   );
   gpc1_1 gpc1962 (
      {stage0_19[354]},
      {stage1_19[168]}
   );
   gpc1_1 gpc1963 (
      {stage0_19[355]},
      {stage1_19[169]}
   );
   gpc1_1 gpc1964 (
      {stage0_19[356]},
      {stage1_19[170]}
   );
   gpc1_1 gpc1965 (
      {stage0_19[357]},
      {stage1_19[171]}
   );
   gpc1_1 gpc1966 (
      {stage0_19[358]},
      {stage1_19[172]}
   );
   gpc1_1 gpc1967 (
      {stage0_19[359]},
      {stage1_19[173]}
   );
   gpc1_1 gpc1968 (
      {stage0_19[360]},
      {stage1_19[174]}
   );
   gpc1_1 gpc1969 (
      {stage0_19[361]},
      {stage1_19[175]}
   );
   gpc1_1 gpc1970 (
      {stage0_19[362]},
      {stage1_19[176]}
   );
   gpc1_1 gpc1971 (
      {stage0_19[363]},
      {stage1_19[177]}
   );
   gpc1_1 gpc1972 (
      {stage0_19[364]},
      {stage1_19[178]}
   );
   gpc1_1 gpc1973 (
      {stage0_19[365]},
      {stage1_19[179]}
   );
   gpc1_1 gpc1974 (
      {stage0_19[366]},
      {stage1_19[180]}
   );
   gpc1_1 gpc1975 (
      {stage0_19[367]},
      {stage1_19[181]}
   );
   gpc1_1 gpc1976 (
      {stage0_19[368]},
      {stage1_19[182]}
   );
   gpc1_1 gpc1977 (
      {stage0_19[369]},
      {stage1_19[183]}
   );
   gpc1_1 gpc1978 (
      {stage0_19[370]},
      {stage1_19[184]}
   );
   gpc1_1 gpc1979 (
      {stage0_19[371]},
      {stage1_19[185]}
   );
   gpc1_1 gpc1980 (
      {stage0_19[372]},
      {stage1_19[186]}
   );
   gpc1_1 gpc1981 (
      {stage0_19[373]},
      {stage1_19[187]}
   );
   gpc1_1 gpc1982 (
      {stage0_19[374]},
      {stage1_19[188]}
   );
   gpc1_1 gpc1983 (
      {stage0_19[375]},
      {stage1_19[189]}
   );
   gpc1_1 gpc1984 (
      {stage0_19[376]},
      {stage1_19[190]}
   );
   gpc1_1 gpc1985 (
      {stage0_19[377]},
      {stage1_19[191]}
   );
   gpc1_1 gpc1986 (
      {stage0_19[378]},
      {stage1_19[192]}
   );
   gpc1_1 gpc1987 (
      {stage0_19[379]},
      {stage1_19[193]}
   );
   gpc1_1 gpc1988 (
      {stage0_19[380]},
      {stage1_19[194]}
   );
   gpc1_1 gpc1989 (
      {stage0_19[381]},
      {stage1_19[195]}
   );
   gpc1_1 gpc1990 (
      {stage0_19[382]},
      {stage1_19[196]}
   );
   gpc1_1 gpc1991 (
      {stage0_19[383]},
      {stage1_19[197]}
   );
   gpc1_1 gpc1992 (
      {stage0_19[384]},
      {stage1_19[198]}
   );
   gpc1_1 gpc1993 (
      {stage0_19[385]},
      {stage1_19[199]}
   );
   gpc1_1 gpc1994 (
      {stage0_19[386]},
      {stage1_19[200]}
   );
   gpc1_1 gpc1995 (
      {stage0_19[387]},
      {stage1_19[201]}
   );
   gpc1_1 gpc1996 (
      {stage0_19[388]},
      {stage1_19[202]}
   );
   gpc1_1 gpc1997 (
      {stage0_19[389]},
      {stage1_19[203]}
   );
   gpc1_1 gpc1998 (
      {stage0_19[390]},
      {stage1_19[204]}
   );
   gpc1_1 gpc1999 (
      {stage0_19[391]},
      {stage1_19[205]}
   );
   gpc1_1 gpc2000 (
      {stage0_19[392]},
      {stage1_19[206]}
   );
   gpc1_1 gpc2001 (
      {stage0_19[393]},
      {stage1_19[207]}
   );
   gpc1_1 gpc2002 (
      {stage0_19[394]},
      {stage1_19[208]}
   );
   gpc1_1 gpc2003 (
      {stage0_19[395]},
      {stage1_19[209]}
   );
   gpc1_1 gpc2004 (
      {stage0_19[396]},
      {stage1_19[210]}
   );
   gpc1_1 gpc2005 (
      {stage0_19[397]},
      {stage1_19[211]}
   );
   gpc1_1 gpc2006 (
      {stage0_19[398]},
      {stage1_19[212]}
   );
   gpc1_1 gpc2007 (
      {stage0_19[399]},
      {stage1_19[213]}
   );
   gpc1_1 gpc2008 (
      {stage0_19[400]},
      {stage1_19[214]}
   );
   gpc1_1 gpc2009 (
      {stage0_19[401]},
      {stage1_19[215]}
   );
   gpc1_1 gpc2010 (
      {stage0_19[402]},
      {stage1_19[216]}
   );
   gpc1_1 gpc2011 (
      {stage0_19[403]},
      {stage1_19[217]}
   );
   gpc1_1 gpc2012 (
      {stage0_19[404]},
      {stage1_19[218]}
   );
   gpc1_1 gpc2013 (
      {stage0_19[405]},
      {stage1_19[219]}
   );
   gpc1_1 gpc2014 (
      {stage0_19[406]},
      {stage1_19[220]}
   );
   gpc1_1 gpc2015 (
      {stage0_19[407]},
      {stage1_19[221]}
   );
   gpc1_1 gpc2016 (
      {stage0_19[408]},
      {stage1_19[222]}
   );
   gpc1_1 gpc2017 (
      {stage0_19[409]},
      {stage1_19[223]}
   );
   gpc1_1 gpc2018 (
      {stage0_19[410]},
      {stage1_19[224]}
   );
   gpc1_1 gpc2019 (
      {stage0_19[411]},
      {stage1_19[225]}
   );
   gpc1_1 gpc2020 (
      {stage0_19[412]},
      {stage1_19[226]}
   );
   gpc1_1 gpc2021 (
      {stage0_19[413]},
      {stage1_19[227]}
   );
   gpc1_1 gpc2022 (
      {stage0_19[414]},
      {stage1_19[228]}
   );
   gpc1_1 gpc2023 (
      {stage0_19[415]},
      {stage1_19[229]}
   );
   gpc1_1 gpc2024 (
      {stage0_19[416]},
      {stage1_19[230]}
   );
   gpc1_1 gpc2025 (
      {stage0_19[417]},
      {stage1_19[231]}
   );
   gpc1_1 gpc2026 (
      {stage0_19[418]},
      {stage1_19[232]}
   );
   gpc1_1 gpc2027 (
      {stage0_19[419]},
      {stage1_19[233]}
   );
   gpc1_1 gpc2028 (
      {stage0_19[420]},
      {stage1_19[234]}
   );
   gpc1_1 gpc2029 (
      {stage0_19[421]},
      {stage1_19[235]}
   );
   gpc1_1 gpc2030 (
      {stage0_19[422]},
      {stage1_19[236]}
   );
   gpc1_1 gpc2031 (
      {stage0_19[423]},
      {stage1_19[237]}
   );
   gpc1_1 gpc2032 (
      {stage0_19[424]},
      {stage1_19[238]}
   );
   gpc1_1 gpc2033 (
      {stage0_19[425]},
      {stage1_19[239]}
   );
   gpc1_1 gpc2034 (
      {stage0_19[426]},
      {stage1_19[240]}
   );
   gpc1_1 gpc2035 (
      {stage0_19[427]},
      {stage1_19[241]}
   );
   gpc1_1 gpc2036 (
      {stage0_19[428]},
      {stage1_19[242]}
   );
   gpc1_1 gpc2037 (
      {stage0_19[429]},
      {stage1_19[243]}
   );
   gpc1_1 gpc2038 (
      {stage0_19[430]},
      {stage1_19[244]}
   );
   gpc1_1 gpc2039 (
      {stage0_19[431]},
      {stage1_19[245]}
   );
   gpc1_1 gpc2040 (
      {stage0_19[432]},
      {stage1_19[246]}
   );
   gpc1_1 gpc2041 (
      {stage0_19[433]},
      {stage1_19[247]}
   );
   gpc1_1 gpc2042 (
      {stage0_19[434]},
      {stage1_19[248]}
   );
   gpc1_1 gpc2043 (
      {stage0_19[435]},
      {stage1_19[249]}
   );
   gpc1_1 gpc2044 (
      {stage0_19[436]},
      {stage1_19[250]}
   );
   gpc1_1 gpc2045 (
      {stage0_19[437]},
      {stage1_19[251]}
   );
   gpc1_1 gpc2046 (
      {stage0_19[438]},
      {stage1_19[252]}
   );
   gpc1_1 gpc2047 (
      {stage0_19[439]},
      {stage1_19[253]}
   );
   gpc1_1 gpc2048 (
      {stage0_19[440]},
      {stage1_19[254]}
   );
   gpc1_1 gpc2049 (
      {stage0_19[441]},
      {stage1_19[255]}
   );
   gpc1_1 gpc2050 (
      {stage0_19[442]},
      {stage1_19[256]}
   );
   gpc1_1 gpc2051 (
      {stage0_19[443]},
      {stage1_19[257]}
   );
   gpc1_1 gpc2052 (
      {stage0_19[444]},
      {stage1_19[258]}
   );
   gpc1_1 gpc2053 (
      {stage0_19[445]},
      {stage1_19[259]}
   );
   gpc1_1 gpc2054 (
      {stage0_19[446]},
      {stage1_19[260]}
   );
   gpc1_1 gpc2055 (
      {stage0_19[447]},
      {stage1_19[261]}
   );
   gpc1_1 gpc2056 (
      {stage0_19[448]},
      {stage1_19[262]}
   );
   gpc1_1 gpc2057 (
      {stage0_19[449]},
      {stage1_19[263]}
   );
   gpc1_1 gpc2058 (
      {stage0_19[450]},
      {stage1_19[264]}
   );
   gpc1_1 gpc2059 (
      {stage0_19[451]},
      {stage1_19[265]}
   );
   gpc1_1 gpc2060 (
      {stage0_19[452]},
      {stage1_19[266]}
   );
   gpc1_1 gpc2061 (
      {stage0_19[453]},
      {stage1_19[267]}
   );
   gpc1_1 gpc2062 (
      {stage0_19[454]},
      {stage1_19[268]}
   );
   gpc1_1 gpc2063 (
      {stage0_19[455]},
      {stage1_19[269]}
   );
   gpc1_1 gpc2064 (
      {stage0_19[456]},
      {stage1_19[270]}
   );
   gpc1_1 gpc2065 (
      {stage0_19[457]},
      {stage1_19[271]}
   );
   gpc1_1 gpc2066 (
      {stage0_19[458]},
      {stage1_19[272]}
   );
   gpc1_1 gpc2067 (
      {stage0_19[459]},
      {stage1_19[273]}
   );
   gpc1_1 gpc2068 (
      {stage0_19[460]},
      {stage1_19[274]}
   );
   gpc1_1 gpc2069 (
      {stage0_19[461]},
      {stage1_19[275]}
   );
   gpc1_1 gpc2070 (
      {stage0_19[462]},
      {stage1_19[276]}
   );
   gpc1_1 gpc2071 (
      {stage0_19[463]},
      {stage1_19[277]}
   );
   gpc1_1 gpc2072 (
      {stage0_19[464]},
      {stage1_19[278]}
   );
   gpc1_1 gpc2073 (
      {stage0_19[465]},
      {stage1_19[279]}
   );
   gpc1_1 gpc2074 (
      {stage0_19[466]},
      {stage1_19[280]}
   );
   gpc1_1 gpc2075 (
      {stage0_19[467]},
      {stage1_19[281]}
   );
   gpc1_1 gpc2076 (
      {stage0_19[468]},
      {stage1_19[282]}
   );
   gpc1_1 gpc2077 (
      {stage0_19[469]},
      {stage1_19[283]}
   );
   gpc1_1 gpc2078 (
      {stage0_19[470]},
      {stage1_19[284]}
   );
   gpc1_1 gpc2079 (
      {stage0_19[471]},
      {stage1_19[285]}
   );
   gpc1_1 gpc2080 (
      {stage0_19[472]},
      {stage1_19[286]}
   );
   gpc1_1 gpc2081 (
      {stage0_19[473]},
      {stage1_19[287]}
   );
   gpc1_1 gpc2082 (
      {stage0_19[474]},
      {stage1_19[288]}
   );
   gpc1_1 gpc2083 (
      {stage0_19[475]},
      {stage1_19[289]}
   );
   gpc1_1 gpc2084 (
      {stage0_19[476]},
      {stage1_19[290]}
   );
   gpc1_1 gpc2085 (
      {stage0_19[477]},
      {stage1_19[291]}
   );
   gpc1_1 gpc2086 (
      {stage0_19[478]},
      {stage1_19[292]}
   );
   gpc1_1 gpc2087 (
      {stage0_19[479]},
      {stage1_19[293]}
   );
   gpc1_1 gpc2088 (
      {stage0_19[480]},
      {stage1_19[294]}
   );
   gpc1_1 gpc2089 (
      {stage0_19[481]},
      {stage1_19[295]}
   );
   gpc1_1 gpc2090 (
      {stage0_19[482]},
      {stage1_19[296]}
   );
   gpc1_1 gpc2091 (
      {stage0_19[483]},
      {stage1_19[297]}
   );
   gpc1_1 gpc2092 (
      {stage0_19[484]},
      {stage1_19[298]}
   );
   gpc1_1 gpc2093 (
      {stage0_19[485]},
      {stage1_19[299]}
   );
   gpc1_1 gpc2094 (
      {stage0_20[478]},
      {stage1_20[181]}
   );
   gpc1_1 gpc2095 (
      {stage0_20[479]},
      {stage1_20[182]}
   );
   gpc1_1 gpc2096 (
      {stage0_20[480]},
      {stage1_20[183]}
   );
   gpc1_1 gpc2097 (
      {stage0_20[481]},
      {stage1_20[184]}
   );
   gpc1_1 gpc2098 (
      {stage0_20[482]},
      {stage1_20[185]}
   );
   gpc1_1 gpc2099 (
      {stage0_20[483]},
      {stage1_20[186]}
   );
   gpc1_1 gpc2100 (
      {stage0_20[484]},
      {stage1_20[187]}
   );
   gpc1_1 gpc2101 (
      {stage0_20[485]},
      {stage1_20[188]}
   );
   gpc1_1 gpc2102 (
      {stage0_22[422]},
      {stage1_22[187]}
   );
   gpc1_1 gpc2103 (
      {stage0_22[423]},
      {stage1_22[188]}
   );
   gpc1_1 gpc2104 (
      {stage0_22[424]},
      {stage1_22[189]}
   );
   gpc1_1 gpc2105 (
      {stage0_22[425]},
      {stage1_22[190]}
   );
   gpc1_1 gpc2106 (
      {stage0_22[426]},
      {stage1_22[191]}
   );
   gpc1_1 gpc2107 (
      {stage0_22[427]},
      {stage1_22[192]}
   );
   gpc1_1 gpc2108 (
      {stage0_22[428]},
      {stage1_22[193]}
   );
   gpc1_1 gpc2109 (
      {stage0_22[429]},
      {stage1_22[194]}
   );
   gpc1_1 gpc2110 (
      {stage0_22[430]},
      {stage1_22[195]}
   );
   gpc1_1 gpc2111 (
      {stage0_22[431]},
      {stage1_22[196]}
   );
   gpc1_1 gpc2112 (
      {stage0_22[432]},
      {stage1_22[197]}
   );
   gpc1_1 gpc2113 (
      {stage0_22[433]},
      {stage1_22[198]}
   );
   gpc1_1 gpc2114 (
      {stage0_22[434]},
      {stage1_22[199]}
   );
   gpc1_1 gpc2115 (
      {stage0_22[435]},
      {stage1_22[200]}
   );
   gpc1_1 gpc2116 (
      {stage0_22[436]},
      {stage1_22[201]}
   );
   gpc1_1 gpc2117 (
      {stage0_22[437]},
      {stage1_22[202]}
   );
   gpc1_1 gpc2118 (
      {stage0_22[438]},
      {stage1_22[203]}
   );
   gpc1_1 gpc2119 (
      {stage0_22[439]},
      {stage1_22[204]}
   );
   gpc1_1 gpc2120 (
      {stage0_22[440]},
      {stage1_22[205]}
   );
   gpc1_1 gpc2121 (
      {stage0_22[441]},
      {stage1_22[206]}
   );
   gpc1_1 gpc2122 (
      {stage0_22[442]},
      {stage1_22[207]}
   );
   gpc1_1 gpc2123 (
      {stage0_22[443]},
      {stage1_22[208]}
   );
   gpc1_1 gpc2124 (
      {stage0_22[444]},
      {stage1_22[209]}
   );
   gpc1_1 gpc2125 (
      {stage0_22[445]},
      {stage1_22[210]}
   );
   gpc1_1 gpc2126 (
      {stage0_22[446]},
      {stage1_22[211]}
   );
   gpc1_1 gpc2127 (
      {stage0_22[447]},
      {stage1_22[212]}
   );
   gpc1_1 gpc2128 (
      {stage0_22[448]},
      {stage1_22[213]}
   );
   gpc1_1 gpc2129 (
      {stage0_22[449]},
      {stage1_22[214]}
   );
   gpc1_1 gpc2130 (
      {stage0_22[450]},
      {stage1_22[215]}
   );
   gpc1_1 gpc2131 (
      {stage0_22[451]},
      {stage1_22[216]}
   );
   gpc1_1 gpc2132 (
      {stage0_22[452]},
      {stage1_22[217]}
   );
   gpc1_1 gpc2133 (
      {stage0_22[453]},
      {stage1_22[218]}
   );
   gpc1_1 gpc2134 (
      {stage0_22[454]},
      {stage1_22[219]}
   );
   gpc1_1 gpc2135 (
      {stage0_22[455]},
      {stage1_22[220]}
   );
   gpc1_1 gpc2136 (
      {stage0_22[456]},
      {stage1_22[221]}
   );
   gpc1_1 gpc2137 (
      {stage0_22[457]},
      {stage1_22[222]}
   );
   gpc1_1 gpc2138 (
      {stage0_22[458]},
      {stage1_22[223]}
   );
   gpc1_1 gpc2139 (
      {stage0_22[459]},
      {stage1_22[224]}
   );
   gpc1_1 gpc2140 (
      {stage0_22[460]},
      {stage1_22[225]}
   );
   gpc1_1 gpc2141 (
      {stage0_22[461]},
      {stage1_22[226]}
   );
   gpc1_1 gpc2142 (
      {stage0_22[462]},
      {stage1_22[227]}
   );
   gpc1_1 gpc2143 (
      {stage0_22[463]},
      {stage1_22[228]}
   );
   gpc1_1 gpc2144 (
      {stage0_22[464]},
      {stage1_22[229]}
   );
   gpc1_1 gpc2145 (
      {stage0_22[465]},
      {stage1_22[230]}
   );
   gpc1_1 gpc2146 (
      {stage0_22[466]},
      {stage1_22[231]}
   );
   gpc1_1 gpc2147 (
      {stage0_22[467]},
      {stage1_22[232]}
   );
   gpc1_1 gpc2148 (
      {stage0_22[468]},
      {stage1_22[233]}
   );
   gpc1_1 gpc2149 (
      {stage0_22[469]},
      {stage1_22[234]}
   );
   gpc1_1 gpc2150 (
      {stage0_22[470]},
      {stage1_22[235]}
   );
   gpc1_1 gpc2151 (
      {stage0_22[471]},
      {stage1_22[236]}
   );
   gpc1_1 gpc2152 (
      {stage0_22[472]},
      {stage1_22[237]}
   );
   gpc1_1 gpc2153 (
      {stage0_22[473]},
      {stage1_22[238]}
   );
   gpc1_1 gpc2154 (
      {stage0_22[474]},
      {stage1_22[239]}
   );
   gpc1_1 gpc2155 (
      {stage0_22[475]},
      {stage1_22[240]}
   );
   gpc1_1 gpc2156 (
      {stage0_22[476]},
      {stage1_22[241]}
   );
   gpc1_1 gpc2157 (
      {stage0_22[477]},
      {stage1_22[242]}
   );
   gpc1_1 gpc2158 (
      {stage0_22[478]},
      {stage1_22[243]}
   );
   gpc1_1 gpc2159 (
      {stage0_22[479]},
      {stage1_22[244]}
   );
   gpc1_1 gpc2160 (
      {stage0_22[480]},
      {stage1_22[245]}
   );
   gpc1_1 gpc2161 (
      {stage0_22[481]},
      {stage1_22[246]}
   );
   gpc1_1 gpc2162 (
      {stage0_22[482]},
      {stage1_22[247]}
   );
   gpc1_1 gpc2163 (
      {stage0_22[483]},
      {stage1_22[248]}
   );
   gpc1_1 gpc2164 (
      {stage0_22[484]},
      {stage1_22[249]}
   );
   gpc1_1 gpc2165 (
      {stage0_22[485]},
      {stage1_22[250]}
   );
   gpc1_1 gpc2166 (
      {stage0_23[474]},
      {stage1_23[166]}
   );
   gpc1_1 gpc2167 (
      {stage0_23[475]},
      {stage1_23[167]}
   );
   gpc1_1 gpc2168 (
      {stage0_23[476]},
      {stage1_23[168]}
   );
   gpc1_1 gpc2169 (
      {stage0_23[477]},
      {stage1_23[169]}
   );
   gpc1_1 gpc2170 (
      {stage0_23[478]},
      {stage1_23[170]}
   );
   gpc1_1 gpc2171 (
      {stage0_23[479]},
      {stage1_23[171]}
   );
   gpc1_1 gpc2172 (
      {stage0_23[480]},
      {stage1_23[172]}
   );
   gpc1_1 gpc2173 (
      {stage0_23[481]},
      {stage1_23[173]}
   );
   gpc1_1 gpc2174 (
      {stage0_23[482]},
      {stage1_23[174]}
   );
   gpc1_1 gpc2175 (
      {stage0_23[483]},
      {stage1_23[175]}
   );
   gpc1_1 gpc2176 (
      {stage0_23[484]},
      {stage1_23[176]}
   );
   gpc1_1 gpc2177 (
      {stage0_23[485]},
      {stage1_23[177]}
   );
   gpc1_1 gpc2178 (
      {stage0_26[445]},
      {stage1_26[174]}
   );
   gpc1_1 gpc2179 (
      {stage0_26[446]},
      {stage1_26[175]}
   );
   gpc1_1 gpc2180 (
      {stage0_26[447]},
      {stage1_26[176]}
   );
   gpc1_1 gpc2181 (
      {stage0_26[448]},
      {stage1_26[177]}
   );
   gpc1_1 gpc2182 (
      {stage0_26[449]},
      {stage1_26[178]}
   );
   gpc1_1 gpc2183 (
      {stage0_26[450]},
      {stage1_26[179]}
   );
   gpc1_1 gpc2184 (
      {stage0_26[451]},
      {stage1_26[180]}
   );
   gpc1_1 gpc2185 (
      {stage0_26[452]},
      {stage1_26[181]}
   );
   gpc1_1 gpc2186 (
      {stage0_26[453]},
      {stage1_26[182]}
   );
   gpc1_1 gpc2187 (
      {stage0_26[454]},
      {stage1_26[183]}
   );
   gpc1_1 gpc2188 (
      {stage0_26[455]},
      {stage1_26[184]}
   );
   gpc1_1 gpc2189 (
      {stage0_26[456]},
      {stage1_26[185]}
   );
   gpc1_1 gpc2190 (
      {stage0_26[457]},
      {stage1_26[186]}
   );
   gpc1_1 gpc2191 (
      {stage0_26[458]},
      {stage1_26[187]}
   );
   gpc1_1 gpc2192 (
      {stage0_26[459]},
      {stage1_26[188]}
   );
   gpc1_1 gpc2193 (
      {stage0_26[460]},
      {stage1_26[189]}
   );
   gpc1_1 gpc2194 (
      {stage0_26[461]},
      {stage1_26[190]}
   );
   gpc1_1 gpc2195 (
      {stage0_26[462]},
      {stage1_26[191]}
   );
   gpc1_1 gpc2196 (
      {stage0_26[463]},
      {stage1_26[192]}
   );
   gpc1_1 gpc2197 (
      {stage0_26[464]},
      {stage1_26[193]}
   );
   gpc1_1 gpc2198 (
      {stage0_26[465]},
      {stage1_26[194]}
   );
   gpc1_1 gpc2199 (
      {stage0_26[466]},
      {stage1_26[195]}
   );
   gpc1_1 gpc2200 (
      {stage0_26[467]},
      {stage1_26[196]}
   );
   gpc1_1 gpc2201 (
      {stage0_26[468]},
      {stage1_26[197]}
   );
   gpc1_1 gpc2202 (
      {stage0_26[469]},
      {stage1_26[198]}
   );
   gpc1_1 gpc2203 (
      {stage0_26[470]},
      {stage1_26[199]}
   );
   gpc1_1 gpc2204 (
      {stage0_26[471]},
      {stage1_26[200]}
   );
   gpc1_1 gpc2205 (
      {stage0_26[472]},
      {stage1_26[201]}
   );
   gpc1_1 gpc2206 (
      {stage0_26[473]},
      {stage1_26[202]}
   );
   gpc1_1 gpc2207 (
      {stage0_26[474]},
      {stage1_26[203]}
   );
   gpc1_1 gpc2208 (
      {stage0_26[475]},
      {stage1_26[204]}
   );
   gpc1_1 gpc2209 (
      {stage0_26[476]},
      {stage1_26[205]}
   );
   gpc1_1 gpc2210 (
      {stage0_26[477]},
      {stage1_26[206]}
   );
   gpc1_1 gpc2211 (
      {stage0_26[478]},
      {stage1_26[207]}
   );
   gpc1_1 gpc2212 (
      {stage0_26[479]},
      {stage1_26[208]}
   );
   gpc1_1 gpc2213 (
      {stage0_26[480]},
      {stage1_26[209]}
   );
   gpc1_1 gpc2214 (
      {stage0_26[481]},
      {stage1_26[210]}
   );
   gpc1_1 gpc2215 (
      {stage0_26[482]},
      {stage1_26[211]}
   );
   gpc1_1 gpc2216 (
      {stage0_26[483]},
      {stage1_26[212]}
   );
   gpc1_1 gpc2217 (
      {stage0_26[484]},
      {stage1_26[213]}
   );
   gpc1_1 gpc2218 (
      {stage0_26[485]},
      {stage1_26[214]}
   );
   gpc1_1 gpc2219 (
      {stage0_27[483]},
      {stage1_27[156]}
   );
   gpc1_1 gpc2220 (
      {stage0_27[484]},
      {stage1_27[157]}
   );
   gpc1_1 gpc2221 (
      {stage0_27[485]},
      {stage1_27[158]}
   );
   gpc1_1 gpc2222 (
      {stage0_28[450]},
      {stage1_28[216]}
   );
   gpc1_1 gpc2223 (
      {stage0_28[451]},
      {stage1_28[217]}
   );
   gpc1_1 gpc2224 (
      {stage0_28[452]},
      {stage1_28[218]}
   );
   gpc1_1 gpc2225 (
      {stage0_28[453]},
      {stage1_28[219]}
   );
   gpc1_1 gpc2226 (
      {stage0_28[454]},
      {stage1_28[220]}
   );
   gpc1_1 gpc2227 (
      {stage0_28[455]},
      {stage1_28[221]}
   );
   gpc1_1 gpc2228 (
      {stage0_28[456]},
      {stage1_28[222]}
   );
   gpc1_1 gpc2229 (
      {stage0_28[457]},
      {stage1_28[223]}
   );
   gpc1_1 gpc2230 (
      {stage0_28[458]},
      {stage1_28[224]}
   );
   gpc1_1 gpc2231 (
      {stage0_28[459]},
      {stage1_28[225]}
   );
   gpc1_1 gpc2232 (
      {stage0_28[460]},
      {stage1_28[226]}
   );
   gpc1_1 gpc2233 (
      {stage0_28[461]},
      {stage1_28[227]}
   );
   gpc1_1 gpc2234 (
      {stage0_28[462]},
      {stage1_28[228]}
   );
   gpc1_1 gpc2235 (
      {stage0_28[463]},
      {stage1_28[229]}
   );
   gpc1_1 gpc2236 (
      {stage0_28[464]},
      {stage1_28[230]}
   );
   gpc1_1 gpc2237 (
      {stage0_28[465]},
      {stage1_28[231]}
   );
   gpc1_1 gpc2238 (
      {stage0_28[466]},
      {stage1_28[232]}
   );
   gpc1_1 gpc2239 (
      {stage0_28[467]},
      {stage1_28[233]}
   );
   gpc1_1 gpc2240 (
      {stage0_28[468]},
      {stage1_28[234]}
   );
   gpc1_1 gpc2241 (
      {stage0_28[469]},
      {stage1_28[235]}
   );
   gpc1_1 gpc2242 (
      {stage0_28[470]},
      {stage1_28[236]}
   );
   gpc1_1 gpc2243 (
      {stage0_28[471]},
      {stage1_28[237]}
   );
   gpc1_1 gpc2244 (
      {stage0_28[472]},
      {stage1_28[238]}
   );
   gpc1_1 gpc2245 (
      {stage0_28[473]},
      {stage1_28[239]}
   );
   gpc1_1 gpc2246 (
      {stage0_28[474]},
      {stage1_28[240]}
   );
   gpc1_1 gpc2247 (
      {stage0_28[475]},
      {stage1_28[241]}
   );
   gpc1_1 gpc2248 (
      {stage0_28[476]},
      {stage1_28[242]}
   );
   gpc1_1 gpc2249 (
      {stage0_28[477]},
      {stage1_28[243]}
   );
   gpc1_1 gpc2250 (
      {stage0_28[478]},
      {stage1_28[244]}
   );
   gpc1_1 gpc2251 (
      {stage0_28[479]},
      {stage1_28[245]}
   );
   gpc1_1 gpc2252 (
      {stage0_28[480]},
      {stage1_28[246]}
   );
   gpc1_1 gpc2253 (
      {stage0_28[481]},
      {stage1_28[247]}
   );
   gpc1_1 gpc2254 (
      {stage0_28[482]},
      {stage1_28[248]}
   );
   gpc1_1 gpc2255 (
      {stage0_28[483]},
      {stage1_28[249]}
   );
   gpc1_1 gpc2256 (
      {stage0_28[484]},
      {stage1_28[250]}
   );
   gpc1_1 gpc2257 (
      {stage0_28[485]},
      {stage1_28[251]}
   );
   gpc1_1 gpc2258 (
      {stage0_30[480]},
      {stage1_30[166]}
   );
   gpc1_1 gpc2259 (
      {stage0_30[481]},
      {stage1_30[167]}
   );
   gpc1_1 gpc2260 (
      {stage0_30[482]},
      {stage1_30[168]}
   );
   gpc1_1 gpc2261 (
      {stage0_30[483]},
      {stage1_30[169]}
   );
   gpc1_1 gpc2262 (
      {stage0_30[484]},
      {stage1_30[170]}
   );
   gpc1_1 gpc2263 (
      {stage0_30[485]},
      {stage1_30[171]}
   );
   gpc1163_5 gpc2264 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc2265 (
      {stage1_0[3], stage1_0[4], stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc2266 (
      {stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc2267 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc606_5 gpc2268 (
      {stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc2269 (
      {stage1_0[27], stage1_0[28], stage1_0[29], stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc2270 (
      {stage1_0[33], stage1_0[34], stage1_0[35], stage1_0[36], stage1_0[37], stage1_0[38]},
      {stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc606_5 gpc2271 (
      {stage1_0[39], stage1_0[40], stage1_0[41], stage1_0[42], stage1_0[43], stage1_0[44]},
      {stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc606_5 gpc2272 (
      {stage1_0[45], stage1_0[46], stage1_0[47], stage1_0[48], stage1_0[49], stage1_0[50]},
      {stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc606_5 gpc2273 (
      {stage1_0[51], stage1_0[52], stage1_0[53], stage1_0[54], stage1_0[55], stage1_0[56]},
      {stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc2274 (
      {stage1_0[57], stage1_0[58], stage1_0[59], stage1_0[60], stage1_0[61], stage1_0[62]},
      {stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59], stage1_2[60]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc606_5 gpc2275 (
      {stage1_0[63], stage1_0[64], stage1_0[65], stage1_0[66], stage1_0[67], stage1_0[68]},
      {stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65], stage1_2[66]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc2276 (
      {stage1_0[69], stage1_0[70], stage1_0[71], stage1_0[72], stage1_0[73], stage1_0[74]},
      {stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71], stage1_2[72]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc2277 (
      {stage1_0[75], stage1_0[76], stage1_0[77], stage1_0[78], stage1_0[79], stage1_0[80]},
      {stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77], stage1_2[78]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc606_5 gpc2278 (
      {stage1_0[81], stage1_0[82], stage1_0[83], stage1_0[84], stage1_0[85], stage1_0[86]},
      {stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82], stage1_2[83], stage1_2[84]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc606_5 gpc2279 (
      {stage1_0[87], stage1_0[88], stage1_0[89], stage1_0[90], stage1_0[91], stage1_0[92]},
      {stage1_2[85], stage1_2[86], stage1_2[87], stage1_2[88], stage1_2[89], stage1_2[90]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc606_5 gpc2280 (
      {stage1_0[93], stage1_0[94], stage1_0[95], stage1_0[96], stage1_0[97], stage1_0[98]},
      {stage1_2[91], stage1_2[92], stage1_2[93], stage1_2[94], stage1_2[95], stage1_2[96]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc606_5 gpc2281 (
      {stage1_0[99], stage1_0[100], stage1_0[101], stage1_0[102], stage1_0[103], stage1_0[104]},
      {stage1_2[97], stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101], stage1_2[102]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc606_5 gpc2282 (
      {stage1_0[105], stage1_0[106], stage1_0[107], stage1_0[108], stage1_0[109], stage1_0[110]},
      {stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106], stage1_2[107], stage1_2[108]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc606_5 gpc2283 (
      {stage1_0[111], stage1_0[112], stage1_0[113], stage1_0[114], stage1_0[115], stage1_0[116]},
      {stage1_2[109], stage1_2[110], stage1_2[111], stage1_2[112], stage1_2[113], stage1_2[114]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc615_5 gpc2284 (
      {stage1_0[117], stage1_0[118], stage1_0[119], stage1_0[120], stage1_0[121]},
      {stage1_1[6]},
      {stage1_2[115], stage1_2[116], stage1_2[117], stage1_2[118], stage1_2[119], stage1_2[120]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc615_5 gpc2285 (
      {stage1_0[122], stage1_0[123], stage1_0[124], stage1_0[125], stage1_0[126]},
      {stage1_1[7]},
      {stage1_2[121], stage1_2[122], stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc606_5 gpc2286 (
      {stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13]},
      {stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6]},
      {stage2_5[0],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc606_5 gpc2287 (
      {stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19]},
      {stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage2_5[1],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc2288 (
      {stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25]},
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18]},
      {stage2_5[2],stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24]}
   );
   gpc606_5 gpc2289 (
      {stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31]},
      {stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24]},
      {stage2_5[3],stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25]}
   );
   gpc606_5 gpc2290 (
      {stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37]},
      {stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30]},
      {stage2_5[4],stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26]}
   );
   gpc606_5 gpc2291 (
      {stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41], stage1_1[42], stage1_1[43]},
      {stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage2_5[5],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc2292 (
      {stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47], stage1_1[48], stage1_1[49]},
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42]},
      {stage2_5[6],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc2293 (
      {stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53], stage1_1[54], stage1_1[55]},
      {stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage2_5[7],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc2294 (
      {stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59], stage1_1[60], stage1_1[61]},
      {stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54]},
      {stage2_5[8],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc2295 (
      {stage1_2[127], stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131], stage1_2[132]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[9],stage2_4[31],stage2_3[31],stage2_2[31]}
   );
   gpc606_5 gpc2296 (
      {stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137], stage1_2[138]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[10],stage2_4[32],stage2_3[32],stage2_2[32]}
   );
   gpc606_5 gpc2297 (
      {stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142], stage1_2[143], stage1_2[144]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[11],stage2_4[33],stage2_3[33],stage2_2[33]}
   );
   gpc606_5 gpc2298 (
      {stage1_2[145], stage1_2[146], stage1_2[147], stage1_2[148], stage1_2[149], stage1_2[150]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[12],stage2_4[34],stage2_3[34],stage2_2[34]}
   );
   gpc606_5 gpc2299 (
      {stage1_2[151], stage1_2[152], stage1_2[153], stage1_2[154], stage1_2[155], stage1_2[156]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[13],stage2_4[35],stage2_3[35],stage2_2[35]}
   );
   gpc606_5 gpc2300 (
      {stage1_2[157], stage1_2[158], stage1_2[159], stage1_2[160], stage1_2[161], stage1_2[162]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[14],stage2_4[36],stage2_3[36],stage2_2[36]}
   );
   gpc606_5 gpc2301 (
      {stage1_2[163], stage1_2[164], stage1_2[165], stage1_2[166], stage1_2[167], stage1_2[168]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[15],stage2_4[37],stage2_3[37],stage2_2[37]}
   );
   gpc606_5 gpc2302 (
      {stage1_2[169], stage1_2[170], stage1_2[171], stage1_2[172], stage1_2[173], stage1_2[174]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[16],stage2_4[38],stage2_3[38],stage2_2[38]}
   );
   gpc606_5 gpc2303 (
      {stage1_2[175], stage1_2[176], stage1_2[177], stage1_2[178], stage1_2[179], stage1_2[180]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[17],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc606_5 gpc2304 (
      {stage1_2[181], stage1_2[182], stage1_2[183], stage1_2[184], stage1_2[185], stage1_2[186]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[18],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc606_5 gpc2305 (
      {stage1_2[187], stage1_2[188], stage1_2[189], stage1_2[190], stage1_2[191], stage1_2[192]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[19],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc606_5 gpc2306 (
      {stage1_2[193], stage1_2[194], stage1_2[195], stage1_2[196], stage1_2[197], stage1_2[198]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[20],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc606_5 gpc2307 (
      {stage1_2[199], stage1_2[200], stage1_2[201], stage1_2[202], stage1_2[203], stage1_2[204]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[21],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc2308 (
      {stage1_2[205], stage1_2[206], stage1_2[207], stage1_2[208], stage1_2[209]},
      {stage1_3[55]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[22],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc615_5 gpc2309 (
      {stage1_2[210], stage1_2[211], stage1_2[212], stage1_2[213], stage1_2[214]},
      {stage1_3[56]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[23],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc615_5 gpc2310 (
      {stage1_2[215], stage1_2[216], stage1_2[217], stage1_2[218], stage1_2[219]},
      {stage1_3[57]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[24],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc615_5 gpc2311 (
      {stage1_2[220], stage1_2[221], stage1_2[222], stage1_2[223], stage1_2[224]},
      {stage1_3[58]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[25],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc606_5 gpc2312 (
      {stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[17],stage2_5[26],stage2_4[48],stage2_3[48]}
   );
   gpc606_5 gpc2313 (
      {stage1_3[65], stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[18],stage2_5[27],stage2_4[49],stage2_3[49]}
   );
   gpc606_5 gpc2314 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[19],stage2_5[28],stage2_4[50],stage2_3[50]}
   );
   gpc606_5 gpc2315 (
      {stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[20],stage2_5[29],stage2_4[51],stage2_3[51]}
   );
   gpc606_5 gpc2316 (
      {stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87], stage1_3[88]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[21],stage2_5[30],stage2_4[52],stage2_3[52]}
   );
   gpc615_5 gpc2317 (
      {stage1_3[89], stage1_3[90], stage1_3[91], stage1_3[92], stage1_3[93]},
      {stage1_4[102]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[22],stage2_5[31],stage2_4[53],stage2_3[53]}
   );
   gpc615_5 gpc2318 (
      {stage1_3[94], stage1_3[95], stage1_3[96], stage1_3[97], stage1_3[98]},
      {stage1_4[103]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[23],stage2_5[32],stage2_4[54],stage2_3[54]}
   );
   gpc615_5 gpc2319 (
      {stage1_3[99], stage1_3[100], stage1_3[101], stage1_3[102], stage1_3[103]},
      {stage1_4[104]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[24],stage2_5[33],stage2_4[55],stage2_3[55]}
   );
   gpc615_5 gpc2320 (
      {stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107], stage1_3[108]},
      {stage1_4[105]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[25],stage2_5[34],stage2_4[56],stage2_3[56]}
   );
   gpc615_5 gpc2321 (
      {stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112], stage1_3[113]},
      {stage1_4[106]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[26],stage2_5[35],stage2_4[57],stage2_3[57]}
   );
   gpc615_5 gpc2322 (
      {stage1_3[114], stage1_3[115], stage1_3[116], stage1_3[117], stage1_3[118]},
      {stage1_4[107]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[27],stage2_5[36],stage2_4[58],stage2_3[58]}
   );
   gpc615_5 gpc2323 (
      {stage1_3[119], stage1_3[120], stage1_3[121], stage1_3[122], stage1_3[123]},
      {stage1_4[108]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[28],stage2_5[37],stage2_4[59],stage2_3[59]}
   );
   gpc615_5 gpc2324 (
      {stage1_3[124], stage1_3[125], stage1_3[126], stage1_3[127], stage1_3[128]},
      {stage1_4[109]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[29],stage2_5[38],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc2325 (
      {stage1_3[129], stage1_3[130], stage1_3[131], stage1_3[132], stage1_3[133]},
      {stage1_4[110]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[30],stage2_5[39],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc2326 (
      {stage1_3[134], stage1_3[135], stage1_3[136], stage1_3[137], stage1_3[138]},
      {stage1_4[111]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[31],stage2_5[40],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc2327 (
      {stage1_3[139], stage1_3[140], stage1_3[141], stage1_3[142], stage1_3[143]},
      {stage1_4[112]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[32],stage2_5[41],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc2328 (
      {stage1_3[144], stage1_3[145], stage1_3[146], stage1_3[147], stage1_3[148]},
      {stage1_4[113]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[33],stage2_5[42],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc2329 (
      {stage1_3[149], stage1_3[150], stage1_3[151], stage1_3[152], stage1_3[153]},
      {stage1_4[114]},
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage2_7[17],stage2_6[34],stage2_5[43],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc2330 (
      {stage1_3[154], stage1_3[155], stage1_3[156], stage1_3[157], stage1_3[158]},
      {stage1_4[115]},
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage2_7[18],stage2_6[35],stage2_5[44],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc2331 (
      {stage1_3[159], stage1_3[160], stage1_3[161], stage1_3[162], stage1_3[163]},
      {stage1_4[116]},
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage2_7[19],stage2_6[36],stage2_5[45],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc2332 (
      {stage1_3[164], stage1_3[165], stage1_3[166], stage1_3[167], stage1_3[168]},
      {stage1_4[117]},
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage2_7[20],stage2_6[37],stage2_5[46],stage2_4[68],stage2_3[68]}
   );
   gpc1163_5 gpc2333 (
      {stage1_4[118], stage1_4[119], stage1_4[120]},
      {stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[21],stage2_6[38],stage2_5[47],stage2_4[69]}
   );
   gpc615_5 gpc2334 (
      {stage1_4[121], stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125]},
      {stage1_5[132]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[22],stage2_6[39],stage2_5[48],stage2_4[70]}
   );
   gpc615_5 gpc2335 (
      {stage1_4[126], stage1_4[127], stage1_4[128], stage1_4[129], stage1_4[130]},
      {stage1_5[133]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[2],stage2_7[23],stage2_6[40],stage2_5[49],stage2_4[71]}
   );
   gpc615_5 gpc2336 (
      {stage1_4[131], stage1_4[132], stage1_4[133], stage1_4[134], stage1_4[135]},
      {stage1_5[134]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[3],stage2_7[24],stage2_6[41],stage2_5[50],stage2_4[72]}
   );
   gpc615_5 gpc2337 (
      {stage1_4[136], stage1_4[137], stage1_4[138], stage1_4[139], stage1_4[140]},
      {stage1_5[135]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[4],stage2_7[25],stage2_6[42],stage2_5[51],stage2_4[73]}
   );
   gpc615_5 gpc2338 (
      {stage1_4[141], stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145]},
      {stage1_5[136]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[5],stage2_7[26],stage2_6[43],stage2_5[52],stage2_4[74]}
   );
   gpc615_5 gpc2339 (
      {stage1_4[146], stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150]},
      {stage1_5[137]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[6],stage2_7[27],stage2_6[44],stage2_5[53],stage2_4[75]}
   );
   gpc615_5 gpc2340 (
      {stage1_4[151], stage1_4[152], stage1_4[153], stage1_4[154], stage1_4[155]},
      {stage1_5[138]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[7],stage2_7[28],stage2_6[45],stage2_5[54],stage2_4[76]}
   );
   gpc615_5 gpc2341 (
      {stage1_4[156], stage1_4[157], stage1_4[158], stage1_4[159], stage1_4[160]},
      {stage1_5[139]},
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage2_8[8],stage2_7[29],stage2_6[46],stage2_5[55],stage2_4[77]}
   );
   gpc615_5 gpc2342 (
      {stage1_4[161], stage1_4[162], stage1_4[163], stage1_4[164], stage1_4[165]},
      {stage1_5[140]},
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54]},
      {stage2_8[9],stage2_7[30],stage2_6[47],stage2_5[56],stage2_4[78]}
   );
   gpc615_5 gpc2343 (
      {stage1_4[166], stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170]},
      {stage1_5[141]},
      {stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage2_8[10],stage2_7[31],stage2_6[48],stage2_5[57],stage2_4[79]}
   );
   gpc615_5 gpc2344 (
      {stage1_4[171], stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175]},
      {stage1_5[142]},
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66]},
      {stage2_8[11],stage2_7[32],stage2_6[49],stage2_5[58],stage2_4[80]}
   );
   gpc615_5 gpc2345 (
      {stage1_4[176], stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180]},
      {stage1_5[143]},
      {stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71], stage1_6[72]},
      {stage2_8[12],stage2_7[33],stage2_6[50],stage2_5[59],stage2_4[81]}
   );
   gpc615_5 gpc2346 (
      {stage1_4[181], stage1_4[182], stage1_4[183], stage1_4[184], stage1_4[185]},
      {stage1_5[144]},
      {stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78]},
      {stage2_8[13],stage2_7[34],stage2_6[51],stage2_5[60],stage2_4[82]}
   );
   gpc615_5 gpc2347 (
      {stage1_4[186], stage1_4[187], stage1_4[188], stage1_4[189], stage1_4[190]},
      {stage1_5[145]},
      {stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84]},
      {stage2_8[14],stage2_7[35],stage2_6[52],stage2_5[61],stage2_4[83]}
   );
   gpc615_5 gpc2348 (
      {stage1_4[191], stage1_4[192], stage1_4[193], stage1_4[194], stage1_4[195]},
      {stage1_5[146]},
      {stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage2_8[15],stage2_7[36],stage2_6[53],stage2_5[62],stage2_4[84]}
   );
   gpc615_5 gpc2349 (
      {stage1_4[196], stage1_4[197], stage1_4[198], stage1_4[199], stage1_4[200]},
      {stage1_5[147]},
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95], stage1_6[96]},
      {stage2_8[16],stage2_7[37],stage2_6[54],stage2_5[63],stage2_4[85]}
   );
   gpc615_5 gpc2350 (
      {stage1_4[201], stage1_4[202], stage1_4[203], stage1_4[204], stage1_4[205]},
      {stage1_5[148]},
      {stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101], stage1_6[102]},
      {stage2_8[17],stage2_7[38],stage2_6[55],stage2_5[64],stage2_4[86]}
   );
   gpc615_5 gpc2351 (
      {stage1_4[206], stage1_4[207], stage1_4[208], stage1_4[209], stage1_4[210]},
      {stage1_5[149]},
      {stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107], stage1_6[108]},
      {stage2_8[18],stage2_7[39],stage2_6[56],stage2_5[65],stage2_4[87]}
   );
   gpc615_5 gpc2352 (
      {stage1_4[211], stage1_4[212], stage1_4[213], stage1_4[214], stage1_4[215]},
      {stage1_5[150]},
      {stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114]},
      {stage2_8[19],stage2_7[40],stage2_6[57],stage2_5[66],stage2_4[88]}
   );
   gpc615_5 gpc2353 (
      {stage1_4[216], stage1_4[217], stage1_4[218], stage1_4[219], stage1_4[220]},
      {stage1_5[151]},
      {stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119], stage1_6[120]},
      {stage2_8[20],stage2_7[41],stage2_6[58],stage2_5[67],stage2_4[89]}
   );
   gpc615_5 gpc2354 (
      {stage1_4[221], stage1_4[222], stage1_4[223], stage1_4[224], stage1_4[225]},
      {stage1_5[152]},
      {stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125], stage1_6[126]},
      {stage2_8[21],stage2_7[42],stage2_6[59],stage2_5[68],stage2_4[90]}
   );
   gpc606_5 gpc2355 (
      {stage1_5[153], stage1_5[154], stage1_5[155], stage1_5[156], stage1_5[157], stage1_5[158]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[22],stage2_7[43],stage2_6[60],stage2_5[69]}
   );
   gpc606_5 gpc2356 (
      {stage1_5[159], stage1_5[160], stage1_5[161], stage1_5[162], stage1_5[163], stage1_5[164]},
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage2_9[1],stage2_8[23],stage2_7[44],stage2_6[61],stage2_5[70]}
   );
   gpc606_5 gpc2357 (
      {stage1_5[165], stage1_5[166], stage1_5[167], stage1_5[168], stage1_5[169], stage1_5[170]},
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18]},
      {stage2_9[2],stage2_8[24],stage2_7[45],stage2_6[62],stage2_5[71]}
   );
   gpc606_5 gpc2358 (
      {stage1_5[171], stage1_5[172], stage1_5[173], stage1_5[174], stage1_5[175], stage1_5[176]},
      {stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24]},
      {stage2_9[3],stage2_8[25],stage2_7[46],stage2_6[63],stage2_5[72]}
   );
   gpc606_5 gpc2359 (
      {stage1_5[177], stage1_5[178], stage1_5[179], stage1_5[180], stage1_5[181], stage1_5[182]},
      {stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30]},
      {stage2_9[4],stage2_8[26],stage2_7[47],stage2_6[64],stage2_5[73]}
   );
   gpc606_5 gpc2360 (
      {stage1_5[183], stage1_5[184], stage1_5[185], stage1_5[186], stage1_5[187], stage1_5[188]},
      {stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36]},
      {stage2_9[5],stage2_8[27],stage2_7[48],stage2_6[65],stage2_5[74]}
   );
   gpc606_5 gpc2361 (
      {stage1_5[189], stage1_5[190], stage1_5[191], stage1_5[192], stage1_5[193], stage1_5[194]},
      {stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42]},
      {stage2_9[6],stage2_8[28],stage2_7[49],stage2_6[66],stage2_5[75]}
   );
   gpc606_5 gpc2362 (
      {stage1_5[195], stage1_5[196], stage1_5[197], stage1_5[198], stage1_5[199], stage1_5[200]},
      {stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage2_9[7],stage2_8[29],stage2_7[50],stage2_6[67],stage2_5[76]}
   );
   gpc606_5 gpc2363 (
      {stage1_5[201], stage1_5[202], stage1_5[203], stage1_5[204], stage1_5[205], stage1_5[206]},
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53], stage1_7[54]},
      {stage2_9[8],stage2_8[30],stage2_7[51],stage2_6[68],stage2_5[77]}
   );
   gpc606_5 gpc2364 (
      {stage1_5[207], stage1_5[208], stage1_5[209], stage1_5[210], stage1_5[211], stage1_5[212]},
      {stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60]},
      {stage2_9[9],stage2_8[31],stage2_7[52],stage2_6[69],stage2_5[78]}
   );
   gpc615_5 gpc2365 (
      {stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131]},
      {stage1_7[61]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[10],stage2_8[32],stage2_7[53],stage2_6[70]}
   );
   gpc615_5 gpc2366 (
      {stage1_6[132], stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136]},
      {stage1_7[62]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[11],stage2_8[33],stage2_7[54],stage2_6[71]}
   );
   gpc615_5 gpc2367 (
      {stage1_6[137], stage1_6[138], stage1_6[139], stage1_6[140], stage1_6[141]},
      {stage1_7[63]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[12],stage2_8[34],stage2_7[55],stage2_6[72]}
   );
   gpc615_5 gpc2368 (
      {stage1_6[142], stage1_6[143], stage1_6[144], stage1_6[145], stage1_6[146]},
      {stage1_7[64]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[13],stage2_8[35],stage2_7[56],stage2_6[73]}
   );
   gpc615_5 gpc2369 (
      {stage1_6[147], stage1_6[148], stage1_6[149], stage1_6[150], stage1_6[151]},
      {stage1_7[65]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[14],stage2_8[36],stage2_7[57],stage2_6[74]}
   );
   gpc615_5 gpc2370 (
      {stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155], stage1_6[156]},
      {stage1_7[66]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[15],stage2_8[37],stage2_7[58],stage2_6[75]}
   );
   gpc615_5 gpc2371 (
      {stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161]},
      {stage1_7[67]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[16],stage2_8[38],stage2_7[59],stage2_6[76]}
   );
   gpc615_5 gpc2372 (
      {stage1_6[162], stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166]},
      {stage1_7[68]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[17],stage2_8[39],stage2_7[60],stage2_6[77]}
   );
   gpc615_5 gpc2373 (
      {stage1_6[167], stage1_6[168], stage1_6[169], stage1_6[170], stage1_6[171]},
      {stage1_7[69]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[18],stage2_8[40],stage2_7[61],stage2_6[78]}
   );
   gpc615_5 gpc2374 (
      {stage1_6[172], stage1_6[173], stage1_6[174], stage1_6[175], stage1_6[176]},
      {stage1_7[70]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[19],stage2_8[41],stage2_7[62],stage2_6[79]}
   );
   gpc615_5 gpc2375 (
      {stage1_6[177], stage1_6[178], stage1_6[179], stage1_6[180], stage1_6[181]},
      {stage1_7[71]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[20],stage2_8[42],stage2_7[63],stage2_6[80]}
   );
   gpc615_5 gpc2376 (
      {stage1_6[182], stage1_6[183], stage1_6[184], stage1_6[185], stage1_6[186]},
      {stage1_7[72]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[21],stage2_8[43],stage2_7[64],stage2_6[81]}
   );
   gpc615_5 gpc2377 (
      {stage1_6[187], stage1_6[188], stage1_6[189], stage1_6[190], stage1_6[191]},
      {stage1_7[73]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[22],stage2_8[44],stage2_7[65],stage2_6[82]}
   );
   gpc615_5 gpc2378 (
      {stage1_6[192], stage1_6[193], stage1_6[194], stage1_6[195], stage1_6[196]},
      {stage1_7[74]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[23],stage2_8[45],stage2_7[66],stage2_6[83]}
   );
   gpc615_5 gpc2379 (
      {stage1_6[197], stage1_6[198], stage1_6[199], stage1_6[200], stage1_6[201]},
      {stage1_7[75]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[24],stage2_8[46],stage2_7[67],stage2_6[84]}
   );
   gpc615_5 gpc2380 (
      {stage1_6[202], stage1_6[203], stage1_6[204], stage1_6[205], stage1_6[206]},
      {stage1_7[76]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[25],stage2_8[47],stage2_7[68],stage2_6[85]}
   );
   gpc615_5 gpc2381 (
      {stage1_6[207], stage1_6[208], stage1_6[209], stage1_6[210], stage1_6[211]},
      {stage1_7[77]},
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage2_10[16],stage2_9[26],stage2_8[48],stage2_7[69],stage2_6[86]}
   );
   gpc615_5 gpc2382 (
      {stage1_6[212], stage1_6[213], stage1_6[214], stage1_6[215], stage1_6[216]},
      {stage1_7[78]},
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage2_10[17],stage2_9[27],stage2_8[49],stage2_7[70],stage2_6[87]}
   );
   gpc615_5 gpc2383 (
      {stage1_6[217], stage1_6[218], stage1_6[219], stage1_6[220], stage1_6[221]},
      {stage1_7[79]},
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage2_10[18],stage2_9[28],stage2_8[50],stage2_7[71],stage2_6[88]}
   );
   gpc615_5 gpc2384 (
      {stage1_6[222], stage1_6[223], stage1_6[224], stage1_6[225], stage1_6[226]},
      {stage1_7[80]},
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage2_10[19],stage2_9[29],stage2_8[51],stage2_7[72],stage2_6[89]}
   );
   gpc615_5 gpc2385 (
      {stage1_6[227], stage1_6[228], stage1_6[229], stage1_6[230], stage1_6[231]},
      {stage1_7[81]},
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage2_10[20],stage2_9[30],stage2_8[52],stage2_7[73],stage2_6[90]}
   );
   gpc615_5 gpc2386 (
      {stage1_6[232], stage1_6[233], stage1_6[234], stage1_6[235], stage1_6[236]},
      {stage1_7[82]},
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage2_10[21],stage2_9[31],stage2_8[53],stage2_7[74],stage2_6[91]}
   );
   gpc615_5 gpc2387 (
      {stage1_6[237], stage1_6[238], stage1_6[239], stage1_6[240], stage1_6[241]},
      {stage1_7[83]},
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage2_10[22],stage2_9[32],stage2_8[54],stage2_7[75],stage2_6[92]}
   );
   gpc615_5 gpc2388 (
      {stage1_6[242], stage1_6[243], stage1_6[244], stage1_6[245], stage1_6[246]},
      {stage1_7[84]},
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage2_10[23],stage2_9[33],stage2_8[55],stage2_7[76],stage2_6[93]}
   );
   gpc615_5 gpc2389 (
      {stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage1_8[144]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[24],stage2_9[34],stage2_8[56],stage2_7[77]}
   );
   gpc615_5 gpc2390 (
      {stage1_7[90], stage1_7[91], stage1_7[92], stage1_7[93], stage1_7[94]},
      {stage1_8[145]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[25],stage2_9[35],stage2_8[57],stage2_7[78]}
   );
   gpc615_5 gpc2391 (
      {stage1_7[95], stage1_7[96], stage1_7[97], stage1_7[98], stage1_7[99]},
      {stage1_8[146]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[26],stage2_9[36],stage2_8[58],stage2_7[79]}
   );
   gpc615_5 gpc2392 (
      {stage1_7[100], stage1_7[101], stage1_7[102], stage1_7[103], stage1_7[104]},
      {stage1_8[147]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[27],stage2_9[37],stage2_8[59],stage2_7[80]}
   );
   gpc615_5 gpc2393 (
      {stage1_7[105], stage1_7[106], stage1_7[107], stage1_7[108], stage1_7[109]},
      {stage1_8[148]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[28],stage2_9[38],stage2_8[60],stage2_7[81]}
   );
   gpc615_5 gpc2394 (
      {stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113], stage1_7[114]},
      {stage1_8[149]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[29],stage2_9[39],stage2_8[61],stage2_7[82]}
   );
   gpc615_5 gpc2395 (
      {stage1_7[115], stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119]},
      {stage1_8[150]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[30],stage2_9[40],stage2_8[62],stage2_7[83]}
   );
   gpc615_5 gpc2396 (
      {stage1_7[120], stage1_7[121], stage1_7[122], stage1_7[123], stage1_7[124]},
      {stage1_8[151]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[31],stage2_9[41],stage2_8[63],stage2_7[84]}
   );
   gpc615_5 gpc2397 (
      {stage1_7[125], stage1_7[126], stage1_7[127], stage1_7[128], stage1_7[129]},
      {stage1_8[152]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[32],stage2_9[42],stage2_8[64],stage2_7[85]}
   );
   gpc615_5 gpc2398 (
      {stage1_7[130], stage1_7[131], stage1_7[132], stage1_7[133], stage1_7[134]},
      {stage1_8[153]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[33],stage2_9[43],stage2_8[65],stage2_7[86]}
   );
   gpc615_5 gpc2399 (
      {stage1_7[135], stage1_7[136], stage1_7[137], stage1_7[138], stage1_7[139]},
      {stage1_8[154]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[34],stage2_9[44],stage2_8[66],stage2_7[87]}
   );
   gpc615_5 gpc2400 (
      {stage1_7[140], stage1_7[141], stage1_7[142], stage1_7[143], stage1_7[144]},
      {stage1_8[155]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[35],stage2_9[45],stage2_8[67],stage2_7[88]}
   );
   gpc615_5 gpc2401 (
      {stage1_7[145], stage1_7[146], stage1_7[147], stage1_7[148], stage1_7[149]},
      {stage1_8[156]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[36],stage2_9[46],stage2_8[68],stage2_7[89]}
   );
   gpc615_5 gpc2402 (
      {stage1_7[150], stage1_7[151], stage1_7[152], stage1_7[153], stage1_7[154]},
      {stage1_8[157]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[37],stage2_9[47],stage2_8[69],stage2_7[90]}
   );
   gpc615_5 gpc2403 (
      {stage1_7[155], stage1_7[156], stage1_7[157], stage1_7[158], stage1_7[159]},
      {stage1_8[158]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[38],stage2_9[48],stage2_8[70],stage2_7[91]}
   );
   gpc615_5 gpc2404 (
      {stage1_7[160], stage1_7[161], stage1_7[162], stage1_7[163], stage1_7[164]},
      {stage1_8[159]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[39],stage2_9[49],stage2_8[71],stage2_7[92]}
   );
   gpc615_5 gpc2405 (
      {stage1_7[165], stage1_7[166], stage1_7[167], stage1_7[168], stage1_7[169]},
      {stage1_8[160]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[40],stage2_9[50],stage2_8[72],stage2_7[93]}
   );
   gpc615_5 gpc2406 (
      {stage1_7[170], stage1_7[171], stage1_7[172], stage1_7[173], stage1_7[174]},
      {stage1_8[161]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[41],stage2_9[51],stage2_8[73],stage2_7[94]}
   );
   gpc615_5 gpc2407 (
      {stage1_7[175], stage1_7[176], stage1_7[177], stage1_7[178], stage1_7[179]},
      {stage1_8[162]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[42],stage2_9[52],stage2_8[74],stage2_7[95]}
   );
   gpc615_5 gpc2408 (
      {stage1_7[180], stage1_7[181], stage1_7[182], stage1_7[183], stage1_7[184]},
      {stage1_8[163]},
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage2_11[19],stage2_10[43],stage2_9[53],stage2_8[75],stage2_7[96]}
   );
   gpc615_5 gpc2409 (
      {stage1_7[185], stage1_7[186], stage1_7[187], stage1_7[188], stage1_7[189]},
      {stage1_8[164]},
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage2_11[20],stage2_10[44],stage2_9[54],stage2_8[76],stage2_7[97]}
   );
   gpc615_5 gpc2410 (
      {stage1_7[190], stage1_7[191], stage1_7[192], stage1_7[193], stage1_7[194]},
      {stage1_8[165]},
      {stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131]},
      {stage2_11[21],stage2_10[45],stage2_9[55],stage2_8[77],stage2_7[98]}
   );
   gpc615_5 gpc2411 (
      {stage1_7[195], stage1_7[196], stage1_7[197], stage1_7[198], stage1_7[199]},
      {stage1_8[166]},
      {stage1_9[132], stage1_9[133], stage1_9[134], stage1_9[135], stage1_9[136], stage1_9[137]},
      {stage2_11[22],stage2_10[46],stage2_9[56],stage2_8[78],stage2_7[99]}
   );
   gpc615_5 gpc2412 (
      {stage1_7[200], stage1_7[201], stage1_7[202], stage1_7[203], stage1_7[204]},
      {stage1_8[167]},
      {stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142], stage1_9[143]},
      {stage2_11[23],stage2_10[47],stage2_9[57],stage2_8[79],stage2_7[100]}
   );
   gpc615_5 gpc2413 (
      {stage1_7[205], stage1_7[206], stage1_7[207], stage1_7[208], stage1_7[209]},
      {stage1_8[168]},
      {stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148], stage1_9[149]},
      {stage2_11[24],stage2_10[48],stage2_9[58],stage2_8[80],stage2_7[101]}
   );
   gpc615_5 gpc2414 (
      {stage1_7[210], stage1_7[211], stage1_7[212], stage1_7[213], stage1_7[214]},
      {stage1_8[169]},
      {stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154], stage1_9[155]},
      {stage2_11[25],stage2_10[49],stage2_9[59],stage2_8[81],stage2_7[102]}
   );
   gpc623_5 gpc2415 (
      {stage1_7[215], stage1_7[216], stage1_7[217]},
      {stage1_8[170], stage1_8[171]},
      {stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160], stage1_9[161]},
      {stage2_11[26],stage2_10[50],stage2_9[60],stage2_8[82],stage2_7[103]}
   );
   gpc1415_5 gpc2416 (
      {stage1_8[172], stage1_8[173], stage1_8[174], stage1_8[175], stage1_8[176]},
      {stage1_9[162]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[27],stage2_10[51],stage2_9[61],stage2_8[83]}
   );
   gpc606_5 gpc2417 (
      {stage1_8[177], stage1_8[178], stage1_8[179], stage1_8[180], stage1_8[181], stage1_8[182]},
      {stage1_10[4], stage1_10[5], stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9]},
      {stage2_12[1],stage2_11[28],stage2_10[52],stage2_9[62],stage2_8[84]}
   );
   gpc606_5 gpc2418 (
      {stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166], stage1_9[167], stage1_9[168]},
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6]},
      {stage2_13[0],stage2_12[2],stage2_11[29],stage2_10[53],stage2_9[63]}
   );
   gpc606_5 gpc2419 (
      {stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172], stage1_9[173], stage1_9[174]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[1],stage2_12[3],stage2_11[30],stage2_10[54],stage2_9[64]}
   );
   gpc606_5 gpc2420 (
      {stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178], stage1_9[179], stage1_9[180]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[2],stage2_12[4],stage2_11[31],stage2_10[55],stage2_9[65]}
   );
   gpc615_5 gpc2421 (
      {stage1_9[181], stage1_9[182], stage1_9[183], stage1_9[184], stage1_9[185]},
      {stage1_10[10]},
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage2_13[3],stage2_12[5],stage2_11[32],stage2_10[56],stage2_9[66]}
   );
   gpc615_5 gpc2422 (
      {stage1_9[186], stage1_9[187], stage1_9[188], stage1_9[189], stage1_9[190]},
      {stage1_10[11]},
      {stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29], stage1_11[30]},
      {stage2_13[4],stage2_12[6],stage2_11[33],stage2_10[57],stage2_9[67]}
   );
   gpc615_5 gpc2423 (
      {stage1_9[191], stage1_9[192], stage1_9[193], stage1_9[194], stage1_9[195]},
      {stage1_10[12]},
      {stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35], stage1_11[36]},
      {stage2_13[5],stage2_12[7],stage2_11[34],stage2_10[58],stage2_9[68]}
   );
   gpc615_5 gpc2424 (
      {stage1_9[196], stage1_9[197], stage1_9[198], stage1_9[199], stage1_9[200]},
      {stage1_10[13]},
      {stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage2_13[6],stage2_12[8],stage2_11[35],stage2_10[59],stage2_9[69]}
   );
   gpc615_5 gpc2425 (
      {stage1_9[201], stage1_9[202], stage1_9[203], stage1_9[204], stage1_9[205]},
      {stage1_10[14]},
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage2_13[7],stage2_12[9],stage2_11[36],stage2_10[60],stage2_9[70]}
   );
   gpc615_5 gpc2426 (
      {stage1_9[206], stage1_9[207], stage1_9[208], stage1_9[209], stage1_9[210]},
      {stage1_10[15]},
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53], stage1_11[54]},
      {stage2_13[8],stage2_12[10],stage2_11[37],stage2_10[61],stage2_9[71]}
   );
   gpc117_4 gpc2427 (
      {stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22]},
      {stage1_11[55]},
      {stage1_12[0]},
      {stage2_13[9],stage2_12[11],stage2_11[38],stage2_10[62]}
   );
   gpc117_4 gpc2428 (
      {stage1_10[23], stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage1_11[56]},
      {stage1_12[1]},
      {stage2_13[10],stage2_12[12],stage2_11[39],stage2_10[63]}
   );
   gpc117_4 gpc2429 (
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36]},
      {stage1_11[57]},
      {stage1_12[2]},
      {stage2_13[11],stage2_12[13],stage2_11[40],stage2_10[64]}
   );
   gpc117_4 gpc2430 (
      {stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41], stage1_10[42], stage1_10[43]},
      {stage1_11[58]},
      {stage1_12[3]},
      {stage2_13[12],stage2_12[14],stage2_11[41],stage2_10[65]}
   );
   gpc117_4 gpc2431 (
      {stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50]},
      {stage1_11[59]},
      {stage1_12[4]},
      {stage2_13[13],stage2_12[15],stage2_11[42],stage2_10[66]}
   );
   gpc117_4 gpc2432 (
      {stage1_10[51], stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57]},
      {stage1_11[60]},
      {stage1_12[5]},
      {stage2_13[14],stage2_12[16],stage2_11[43],stage2_10[67]}
   );
   gpc117_4 gpc2433 (
      {stage1_10[58], stage1_10[59], stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64]},
      {stage1_11[61]},
      {stage1_12[6]},
      {stage2_13[15],stage2_12[17],stage2_11[44],stage2_10[68]}
   );
   gpc117_4 gpc2434 (
      {stage1_10[65], stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage1_11[62]},
      {stage1_12[7]},
      {stage2_13[16],stage2_12[18],stage2_11[45],stage2_10[69]}
   );
   gpc117_4 gpc2435 (
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77], stage1_10[78]},
      {stage1_11[63]},
      {stage1_12[8]},
      {stage2_13[17],stage2_12[19],stage2_11[46],stage2_10[70]}
   );
   gpc117_4 gpc2436 (
      {stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83], stage1_10[84], stage1_10[85]},
      {stage1_11[64]},
      {stage1_12[9]},
      {stage2_13[18],stage2_12[20],stage2_11[47],stage2_10[71]}
   );
   gpc117_4 gpc2437 (
      {stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89], stage1_10[90], stage1_10[91], stage1_10[92]},
      {stage1_11[65]},
      {stage1_12[10]},
      {stage2_13[19],stage2_12[21],stage2_11[48],stage2_10[72]}
   );
   gpc117_4 gpc2438 (
      {stage1_10[93], stage1_10[94], stage1_10[95], stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99]},
      {stage1_11[66]},
      {stage1_12[11]},
      {stage2_13[20],stage2_12[22],stage2_11[49],stage2_10[73]}
   );
   gpc117_4 gpc2439 (
      {stage1_10[100], stage1_10[101], stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106]},
      {stage1_11[67]},
      {stage1_12[12]},
      {stage2_13[21],stage2_12[23],stage2_11[50],stage2_10[74]}
   );
   gpc117_4 gpc2440 (
      {stage1_10[107], stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage1_11[68]},
      {stage1_12[13]},
      {stage2_13[22],stage2_12[24],stage2_11[51],stage2_10[75]}
   );
   gpc117_4 gpc2441 (
      {stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119], stage1_10[120]},
      {stage1_11[69]},
      {stage1_12[14]},
      {stage2_13[23],stage2_12[25],stage2_11[52],stage2_10[76]}
   );
   gpc117_4 gpc2442 (
      {stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124], stage1_10[125], stage1_10[126], stage1_10[127]},
      {stage1_11[70]},
      {stage1_12[15]},
      {stage2_13[24],stage2_12[26],stage2_11[53],stage2_10[77]}
   );
   gpc117_4 gpc2443 (
      {stage1_10[128], stage1_10[129], stage1_10[130], stage1_10[131], stage1_10[132], stage1_10[133], stage1_10[134]},
      {stage1_11[71]},
      {stage1_12[16]},
      {stage2_13[25],stage2_12[27],stage2_11[54],stage2_10[78]}
   );
   gpc117_4 gpc2444 (
      {stage1_10[135], stage1_10[136], stage1_10[137], stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141]},
      {stage1_11[72]},
      {stage1_12[17]},
      {stage2_13[26],stage2_12[28],stage2_11[55],stage2_10[79]}
   );
   gpc117_4 gpc2445 (
      {stage1_10[142], stage1_10[143], stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148]},
      {stage1_11[73]},
      {stage1_12[18]},
      {stage2_13[27],stage2_12[29],stage2_11[56],stage2_10[80]}
   );
   gpc117_4 gpc2446 (
      {stage1_10[149], stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154], stage1_10[155]},
      {stage1_11[74]},
      {stage1_12[19]},
      {stage2_13[28],stage2_12[30],stage2_11[57],stage2_10[81]}
   );
   gpc606_5 gpc2447 (
      {stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160], stage1_10[161]},
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage2_14[0],stage2_13[29],stage2_12[31],stage2_11[58],stage2_10[82]}
   );
   gpc606_5 gpc2448 (
      {stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166], stage1_10[167]},
      {stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31]},
      {stage2_14[1],stage2_13[30],stage2_12[32],stage2_11[59],stage2_10[83]}
   );
   gpc606_5 gpc2449 (
      {stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171], stage1_10[172], stage1_10[173]},
      {stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35], stage1_12[36], stage1_12[37]},
      {stage2_14[2],stage2_13[31],stage2_12[33],stage2_11[60],stage2_10[84]}
   );
   gpc606_5 gpc2450 (
      {stage1_10[174], stage1_10[175], stage1_10[176], stage1_10[177], stage1_10[178], stage1_10[179]},
      {stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41], stage1_12[42], stage1_12[43]},
      {stage2_14[3],stage2_13[32],stage2_12[34],stage2_11[61],stage2_10[85]}
   );
   gpc606_5 gpc2451 (
      {stage1_10[180], stage1_10[181], stage1_10[182], stage1_10[183], stage1_10[184], stage1_10[185]},
      {stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47], stage1_12[48], stage1_12[49]},
      {stage2_14[4],stage2_13[33],stage2_12[35],stage2_11[62],stage2_10[86]}
   );
   gpc615_5 gpc2452 (
      {stage1_11[75], stage1_11[76], stage1_11[77], stage1_11[78], stage1_11[79]},
      {stage1_12[50]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[5],stage2_13[34],stage2_12[36],stage2_11[63]}
   );
   gpc615_5 gpc2453 (
      {stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83], stage1_11[84]},
      {stage1_12[51]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[6],stage2_13[35],stage2_12[37],stage2_11[64]}
   );
   gpc615_5 gpc2454 (
      {stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage1_12[52]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[7],stage2_13[36],stage2_12[38],stage2_11[65]}
   );
   gpc615_5 gpc2455 (
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94]},
      {stage1_12[53]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[8],stage2_13[37],stage2_12[39],stage2_11[66]}
   );
   gpc615_5 gpc2456 (
      {stage1_11[95], stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99]},
      {stage1_12[54]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[9],stage2_13[38],stage2_12[40],stage2_11[67]}
   );
   gpc615_5 gpc2457 (
      {stage1_11[100], stage1_11[101], stage1_11[102], stage1_11[103], stage1_11[104]},
      {stage1_12[55]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[10],stage2_13[39],stage2_12[41],stage2_11[68]}
   );
   gpc615_5 gpc2458 (
      {stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108], stage1_11[109]},
      {stage1_12[56]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[11],stage2_13[40],stage2_12[42],stage2_11[69]}
   );
   gpc615_5 gpc2459 (
      {stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_12[57]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[12],stage2_13[41],stage2_12[43],stage2_11[70]}
   );
   gpc615_5 gpc2460 (
      {stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119]},
      {stage1_12[58]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[13],stage2_13[42],stage2_12[44],stage2_11[71]}
   );
   gpc615_5 gpc2461 (
      {stage1_11[120], stage1_11[121], stage1_11[122], stage1_11[123], stage1_11[124]},
      {stage1_12[59]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[14],stage2_13[43],stage2_12[45],stage2_11[72]}
   );
   gpc615_5 gpc2462 (
      {stage1_11[125], stage1_11[126], stage1_11[127], stage1_11[128], stage1_11[129]},
      {stage1_12[60]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[15],stage2_13[44],stage2_12[46],stage2_11[73]}
   );
   gpc615_5 gpc2463 (
      {stage1_11[130], stage1_11[131], stage1_11[132], stage1_11[133], stage1_11[134]},
      {stage1_12[61]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[16],stage2_13[45],stage2_12[47],stage2_11[74]}
   );
   gpc615_5 gpc2464 (
      {stage1_11[135], stage1_11[136], stage1_11[137], stage1_11[138], stage1_11[139]},
      {stage1_12[62]},
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage2_15[12],stage2_14[17],stage2_13[46],stage2_12[48],stage2_11[75]}
   );
   gpc615_5 gpc2465 (
      {stage1_11[140], stage1_11[141], stage1_11[142], stage1_11[143], stage1_11[144]},
      {stage1_12[63]},
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage2_15[13],stage2_14[18],stage2_13[47],stage2_12[49],stage2_11[76]}
   );
   gpc615_5 gpc2466 (
      {stage1_11[145], stage1_11[146], stage1_11[147], stage1_11[148], stage1_11[149]},
      {stage1_12[64]},
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage2_15[14],stage2_14[19],stage2_13[48],stage2_12[50],stage2_11[77]}
   );
   gpc615_5 gpc2467 (
      {stage1_11[150], stage1_11[151], stage1_11[152], stage1_11[153], stage1_11[154]},
      {stage1_12[65]},
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage2_15[15],stage2_14[20],stage2_13[49],stage2_12[51],stage2_11[78]}
   );
   gpc615_5 gpc2468 (
      {stage1_11[155], stage1_11[156], stage1_11[157], stage1_11[158], stage1_11[159]},
      {stage1_12[66]},
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage2_15[16],stage2_14[21],stage2_13[50],stage2_12[52],stage2_11[79]}
   );
   gpc615_5 gpc2469 (
      {stage1_11[160], stage1_11[161], stage1_11[162], stage1_11[163], stage1_11[164]},
      {stage1_12[67]},
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage2_15[17],stage2_14[22],stage2_13[51],stage2_12[53],stage2_11[80]}
   );
   gpc615_5 gpc2470 (
      {stage1_11[165], stage1_11[166], stage1_11[167], stage1_11[168], stage1_11[169]},
      {stage1_12[68]},
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage2_15[18],stage2_14[23],stage2_13[52],stage2_12[54],stage2_11[81]}
   );
   gpc615_5 gpc2471 (
      {stage1_11[170], stage1_11[171], stage1_11[172], stage1_11[173], stage1_11[174]},
      {stage1_12[69]},
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage2_15[19],stage2_14[24],stage2_13[53],stage2_12[55],stage2_11[82]}
   );
   gpc615_5 gpc2472 (
      {stage1_11[175], stage1_11[176], stage1_11[177], stage1_11[178], stage1_11[179]},
      {stage1_12[70]},
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage2_15[20],stage2_14[25],stage2_13[54],stage2_12[56],stage2_11[83]}
   );
   gpc615_5 gpc2473 (
      {stage1_11[180], stage1_11[181], stage1_11[182], stage1_11[183], stage1_11[184]},
      {stage1_12[71]},
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage2_15[21],stage2_14[26],stage2_13[55],stage2_12[57],stage2_11[84]}
   );
   gpc615_5 gpc2474 (
      {stage1_11[185], stage1_11[186], stage1_11[187], stage1_11[188], stage1_11[189]},
      {stage1_12[72]},
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136], stage1_13[137]},
      {stage2_15[22],stage2_14[27],stage2_13[56],stage2_12[58],stage2_11[85]}
   );
   gpc615_5 gpc2475 (
      {stage1_11[190], stage1_11[191], stage1_11[192], stage1_11[193], stage1_11[194]},
      {stage1_12[73]},
      {stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141], stage1_13[142], stage1_13[143]},
      {stage2_15[23],stage2_14[28],stage2_13[57],stage2_12[59],stage2_11[86]}
   );
   gpc615_5 gpc2476 (
      {stage1_11[195], stage1_11[196], stage1_11[197], stage1_11[198], stage1_11[199]},
      {stage1_12[74]},
      {stage1_13[144], stage1_13[145], stage1_13[146], stage1_13[147], stage1_13[148], stage1_13[149]},
      {stage2_15[24],stage2_14[29],stage2_13[58],stage2_12[60],stage2_11[87]}
   );
   gpc615_5 gpc2477 (
      {stage1_11[200], stage1_11[201], stage1_11[202], stage1_11[203], stage1_11[204]},
      {stage1_12[75]},
      {stage1_13[150], stage1_13[151], stage1_13[152], stage1_13[153], stage1_13[154], stage1_13[155]},
      {stage2_15[25],stage2_14[30],stage2_13[59],stage2_12[61],stage2_11[88]}
   );
   gpc615_5 gpc2478 (
      {stage1_11[205], stage1_11[206], stage1_11[207], stage1_11[208], stage1_11[209]},
      {stage1_12[76]},
      {stage1_13[156], stage1_13[157], stage1_13[158], stage1_13[159], stage1_13[160], stage1_13[161]},
      {stage2_15[26],stage2_14[31],stage2_13[60],stage2_12[62],stage2_11[89]}
   );
   gpc615_5 gpc2479 (
      {stage1_11[210], stage1_11[211], stage1_11[212], stage1_11[213], stage1_11[214]},
      {stage1_12[77]},
      {stage1_13[162], stage1_13[163], stage1_13[164], stage1_13[165], stage1_13[166], stage1_13[167]},
      {stage2_15[27],stage2_14[32],stage2_13[61],stage2_12[63],stage2_11[90]}
   );
   gpc615_5 gpc2480 (
      {stage1_11[215], stage1_11[216], stage1_11[217], stage1_11[218], stage1_11[219]},
      {stage1_12[78]},
      {stage1_13[168], stage1_13[169], stage1_13[170], stage1_13[171], stage1_13[172], stage1_13[173]},
      {stage2_15[28],stage2_14[33],stage2_13[62],stage2_12[64],stage2_11[91]}
   );
   gpc606_5 gpc2481 (
      {stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83], stage1_12[84]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[29],stage2_14[34],stage2_13[63],stage2_12[65]}
   );
   gpc606_5 gpc2482 (
      {stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89], stage1_12[90]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[30],stage2_14[35],stage2_13[64],stage2_12[66]}
   );
   gpc606_5 gpc2483 (
      {stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95], stage1_12[96]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[31],stage2_14[36],stage2_13[65],stage2_12[67]}
   );
   gpc606_5 gpc2484 (
      {stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101], stage1_12[102]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[32],stage2_14[37],stage2_13[66],stage2_12[68]}
   );
   gpc606_5 gpc2485 (
      {stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107], stage1_12[108]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[33],stage2_14[38],stage2_13[67],stage2_12[69]}
   );
   gpc606_5 gpc2486 (
      {stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113], stage1_12[114]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[34],stage2_14[39],stage2_13[68],stage2_12[70]}
   );
   gpc606_5 gpc2487 (
      {stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119], stage1_12[120]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[35],stage2_14[40],stage2_13[69],stage2_12[71]}
   );
   gpc606_5 gpc2488 (
      {stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125], stage1_12[126]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[36],stage2_14[41],stage2_13[70],stage2_12[72]}
   );
   gpc606_5 gpc2489 (
      {stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131], stage1_12[132]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[37],stage2_14[42],stage2_13[71],stage2_12[73]}
   );
   gpc606_5 gpc2490 (
      {stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136], stage1_12[137], stage1_12[138]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[38],stage2_14[43],stage2_13[72],stage2_12[74]}
   );
   gpc606_5 gpc2491 (
      {stage1_12[139], stage1_12[140], stage1_12[141], stage1_12[142], stage1_12[143], stage1_12[144]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[39],stage2_14[44],stage2_13[73],stage2_12[75]}
   );
   gpc606_5 gpc2492 (
      {stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148], stage1_12[149], stage1_12[150]},
      {stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage2_16[11],stage2_15[40],stage2_14[45],stage2_13[74],stage2_12[76]}
   );
   gpc606_5 gpc2493 (
      {stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154], stage1_12[155], stage1_12[156]},
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage2_16[12],stage2_15[41],stage2_14[46],stage2_13[75],stage2_12[77]}
   );
   gpc606_5 gpc2494 (
      {stage1_12[157], stage1_12[158], stage1_12[159], stage1_12[160], stage1_12[161], stage1_12[162]},
      {stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage2_16[13],stage2_15[42],stage2_14[47],stage2_13[76],stage2_12[78]}
   );
   gpc606_5 gpc2495 (
      {stage1_12[163], stage1_12[164], stage1_12[165], stage1_12[166], stage1_12[167], stage1_12[168]},
      {stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage2_16[14],stage2_15[43],stage2_14[48],stage2_13[77],stage2_12[79]}
   );
   gpc606_5 gpc2496 (
      {stage1_12[169], stage1_12[170], stage1_12[171], stage1_12[172], stage1_12[173], stage1_12[174]},
      {stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage2_16[15],stage2_15[44],stage2_14[49],stage2_13[78],stage2_12[80]}
   );
   gpc606_5 gpc2497 (
      {stage1_12[175], stage1_12[176], stage1_12[177], stage1_12[178], stage1_12[179], stage1_12[180]},
      {stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage2_16[16],stage2_15[45],stage2_14[50],stage2_13[79],stage2_12[81]}
   );
   gpc606_5 gpc2498 (
      {stage1_12[181], stage1_12[182], stage1_12[183], stage1_12[184], stage1_12[185], stage1_12[186]},
      {stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106], stage1_14[107]},
      {stage2_16[17],stage2_15[46],stage2_14[51],stage2_13[80],stage2_12[82]}
   );
   gpc606_5 gpc2499 (
      {stage1_12[187], stage1_12[188], stage1_12[189], stage1_12[190], stage1_12[191], stage1_12[192]},
      {stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111], stage1_14[112], stage1_14[113]},
      {stage2_16[18],stage2_15[47],stage2_14[52],stage2_13[81],stage2_12[83]}
   );
   gpc606_5 gpc2500 (
      {stage1_12[193], stage1_12[194], stage1_12[195], stage1_12[196], stage1_12[197], stage1_12[198]},
      {stage1_14[114], stage1_14[115], stage1_14[116], stage1_14[117], stage1_14[118], stage1_14[119]},
      {stage2_16[19],stage2_15[48],stage2_14[53],stage2_13[82],stage2_12[84]}
   );
   gpc606_5 gpc2501 (
      {stage1_12[199], stage1_12[200], stage1_12[201], stage1_12[202], stage1_12[203], stage1_12[204]},
      {stage1_14[120], stage1_14[121], stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125]},
      {stage2_16[20],stage2_15[49],stage2_14[54],stage2_13[83],stage2_12[85]}
   );
   gpc606_5 gpc2502 (
      {stage1_12[205], stage1_12[206], stage1_12[207], stage1_12[208], stage1_12[209], stage1_12[210]},
      {stage1_14[126], stage1_14[127], stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage2_16[21],stage2_15[50],stage2_14[55],stage2_13[84],stage2_12[86]}
   );
   gpc606_5 gpc2503 (
      {stage1_12[211], stage1_12[212], stage1_12[213], stage1_12[214], stage1_12[215], stage1_12[216]},
      {stage1_14[132], stage1_14[133], stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137]},
      {stage2_16[22],stage2_15[51],stage2_14[56],stage2_13[85],stage2_12[87]}
   );
   gpc606_5 gpc2504 (
      {stage1_12[217], stage1_12[218], stage1_12[219], stage1_12[220], stage1_12[221], stage1_12[222]},
      {stage1_14[138], stage1_14[139], stage1_14[140], stage1_14[141], stage1_14[142], stage1_14[143]},
      {stage2_16[23],stage2_15[52],stage2_14[57],stage2_13[86],stage2_12[88]}
   );
   gpc606_5 gpc2505 (
      {stage1_12[223], stage1_12[224], stage1_12[225], stage1_12[226], stage1_12[227], stage1_12[228]},
      {stage1_14[144], stage1_14[145], stage1_14[146], stage1_14[147], stage1_14[148], stage1_14[149]},
      {stage2_16[24],stage2_15[53],stage2_14[58],stage2_13[87],stage2_12[89]}
   );
   gpc606_5 gpc2506 (
      {stage1_12[229], stage1_12[230], stage1_12[231], stage1_12[232], stage1_12[233], stage1_12[234]},
      {stage1_14[150], stage1_14[151], stage1_14[152], stage1_14[153], stage1_14[154], stage1_14[155]},
      {stage2_16[25],stage2_15[54],stage2_14[59],stage2_13[88],stage2_12[90]}
   );
   gpc606_5 gpc2507 (
      {stage1_12[235], stage1_12[236], stage1_12[237], stage1_12[238], stage1_12[239], stage1_12[240]},
      {stage1_14[156], stage1_14[157], stage1_14[158], stage1_14[159], stage1_14[160], stage1_14[161]},
      {stage2_16[26],stage2_15[55],stage2_14[60],stage2_13[89],stage2_12[91]}
   );
   gpc606_5 gpc2508 (
      {stage1_12[241], stage1_12[242], stage1_12[243], stage1_12[244], stage1_12[245], stage1_12[246]},
      {stage1_14[162], stage1_14[163], stage1_14[164], stage1_14[165], stage1_14[166], stage1_14[167]},
      {stage2_16[27],stage2_15[56],stage2_14[61],stage2_13[90],stage2_12[92]}
   );
   gpc606_5 gpc2509 (
      {stage1_12[247], stage1_12[248], stage1_12[249], stage1_12[250], stage1_12[251], stage1_12[252]},
      {stage1_14[168], stage1_14[169], stage1_14[170], stage1_14[171], stage1_14[172], stage1_14[173]},
      {stage2_16[28],stage2_15[57],stage2_14[62],stage2_13[91],stage2_12[93]}
   );
   gpc606_5 gpc2510 (
      {stage1_12[253], stage1_12[254], stage1_12[255], stage1_12[256], stage1_12[257], stage1_12[258]},
      {stage1_14[174], stage1_14[175], stage1_14[176], stage1_14[177], stage1_14[178], stage1_14[179]},
      {stage2_16[29],stage2_15[58],stage2_14[63],stage2_13[92],stage2_12[94]}
   );
   gpc606_5 gpc2511 (
      {stage1_12[259], stage1_12[260], stage1_12[261], stage1_12[262], stage1_12[263], stage1_12[264]},
      {stage1_14[180], stage1_14[181], stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185]},
      {stage2_16[30],stage2_15[59],stage2_14[64],stage2_13[93],stage2_12[95]}
   );
   gpc606_5 gpc2512 (
      {stage1_12[265], stage1_12[266], stage1_12[267], stage1_12[268], stage1_12[269], stage1_12[270]},
      {stage1_14[186], stage1_14[187], stage1_14[188], stage1_14[189], stage1_14[190], stage1_14[191]},
      {stage2_16[31],stage2_15[60],stage2_14[65],stage2_13[94],stage2_12[96]}
   );
   gpc606_5 gpc2513 (
      {stage1_12[271], stage1_12[272], stage1_12[273], stage1_12[274], stage1_12[275], stage1_12[276]},
      {stage1_14[192], stage1_14[193], stage1_14[194], stage1_14[195], stage1_14[196], stage1_14[197]},
      {stage2_16[32],stage2_15[61],stage2_14[66],stage2_13[95],stage2_12[97]}
   );
   gpc606_5 gpc2514 (
      {stage1_13[174], stage1_13[175], stage1_13[176], stage1_13[177], stage1_13[178], stage1_13[179]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[33],stage2_15[62],stage2_14[67],stage2_13[96]}
   );
   gpc615_5 gpc2515 (
      {stage1_13[180], stage1_13[181], stage1_13[182], stage1_13[183], stage1_13[184]},
      {stage1_14[198]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[34],stage2_15[63],stage2_14[68],stage2_13[97]}
   );
   gpc615_5 gpc2516 (
      {stage1_13[185], stage1_13[186], stage1_13[187], stage1_13[188], stage1_13[189]},
      {stage1_14[199]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[35],stage2_15[64],stage2_14[69],stage2_13[98]}
   );
   gpc615_5 gpc2517 (
      {stage1_13[190], stage1_13[191], stage1_13[192], stage1_13[193], stage1_13[194]},
      {stage1_14[200]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[36],stage2_15[65],stage2_14[70],stage2_13[99]}
   );
   gpc615_5 gpc2518 (
      {stage1_13[195], stage1_13[196], stage1_13[197], stage1_13[198], stage1_13[199]},
      {stage1_14[201]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[37],stage2_15[66],stage2_14[71],stage2_13[100]}
   );
   gpc615_5 gpc2519 (
      {stage1_13[200], stage1_13[201], stage1_13[202], stage1_13[203], stage1_13[204]},
      {stage1_14[202]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[38],stage2_15[67],stage2_14[72],stage2_13[101]}
   );
   gpc615_5 gpc2520 (
      {stage1_14[203], stage1_14[204], stage1_14[205], stage1_14[206], stage1_14[207]},
      {stage1_15[36]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[6],stage2_16[39],stage2_15[68],stage2_14[73]}
   );
   gpc615_5 gpc2521 (
      {stage1_14[208], stage1_14[209], stage1_14[210], stage1_14[211], stage1_14[212]},
      {stage1_15[37]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[7],stage2_16[40],stage2_15[69],stage2_14[74]}
   );
   gpc615_5 gpc2522 (
      {stage1_14[213], stage1_14[214], stage1_14[215], stage1_14[216], stage1_14[217]},
      {stage1_15[38]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[8],stage2_16[41],stage2_15[70],stage2_14[75]}
   );
   gpc615_5 gpc2523 (
      {stage1_14[218], stage1_14[219], stage1_14[220], stage1_14[221], stage1_14[222]},
      {stage1_15[39]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[9],stage2_16[42],stage2_15[71],stage2_14[76]}
   );
   gpc615_5 gpc2524 (
      {stage1_14[223], stage1_14[224], stage1_14[225], stage1_14[226], stage1_14[227]},
      {stage1_15[40]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[10],stage2_16[43],stage2_15[72],stage2_14[77]}
   );
   gpc615_5 gpc2525 (
      {stage1_14[228], stage1_14[229], stage1_14[230], stage1_14[231], stage1_14[232]},
      {stage1_15[41]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[11],stage2_16[44],stage2_15[73],stage2_14[78]}
   );
   gpc615_5 gpc2526 (
      {stage1_14[233], stage1_14[234], stage1_14[235], stage1_14[236], stage1_14[237]},
      {stage1_15[42]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[12],stage2_16[45],stage2_15[74],stage2_14[79]}
   );
   gpc615_5 gpc2527 (
      {stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage1_16[42]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[7],stage2_17[13],stage2_16[46],stage2_15[75]}
   );
   gpc615_5 gpc2528 (
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52]},
      {stage1_16[43]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[8],stage2_17[14],stage2_16[47],stage2_15[76]}
   );
   gpc615_5 gpc2529 (
      {stage1_15[53], stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57]},
      {stage1_16[44]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[9],stage2_17[15],stage2_16[48],stage2_15[77]}
   );
   gpc615_5 gpc2530 (
      {stage1_15[58], stage1_15[59], stage1_15[60], stage1_15[61], stage1_15[62]},
      {stage1_16[45]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[10],stage2_17[16],stage2_16[49],stage2_15[78]}
   );
   gpc615_5 gpc2531 (
      {stage1_15[63], stage1_15[64], stage1_15[65], stage1_15[66], stage1_15[67]},
      {stage1_16[46]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[11],stage2_17[17],stage2_16[50],stage2_15[79]}
   );
   gpc615_5 gpc2532 (
      {stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71], stage1_15[72]},
      {stage1_16[47]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[12],stage2_17[18],stage2_16[51],stage2_15[80]}
   );
   gpc615_5 gpc2533 (
      {stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage1_16[48]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[13],stage2_17[19],stage2_16[52],stage2_15[81]}
   );
   gpc615_5 gpc2534 (
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82]},
      {stage1_16[49]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[14],stage2_17[20],stage2_16[53],stage2_15[82]}
   );
   gpc615_5 gpc2535 (
      {stage1_15[83], stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87]},
      {stage1_16[50]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[15],stage2_17[21],stage2_16[54],stage2_15[83]}
   );
   gpc615_5 gpc2536 (
      {stage1_15[88], stage1_15[89], stage1_15[90], stage1_15[91], stage1_15[92]},
      {stage1_16[51]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[16],stage2_17[22],stage2_16[55],stage2_15[84]}
   );
   gpc615_5 gpc2537 (
      {stage1_15[93], stage1_15[94], stage1_15[95], stage1_15[96], stage1_15[97]},
      {stage1_16[52]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage2_19[10],stage2_18[17],stage2_17[23],stage2_16[56],stage2_15[85]}
   );
   gpc615_5 gpc2538 (
      {stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101], stage1_15[102]},
      {stage1_16[53]},
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage2_19[11],stage2_18[18],stage2_17[24],stage2_16[57],stage2_15[86]}
   );
   gpc615_5 gpc2539 (
      {stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage1_16[54]},
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage2_19[12],stage2_18[19],stage2_17[25],stage2_16[58],stage2_15[87]}
   );
   gpc615_5 gpc2540 (
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112]},
      {stage1_16[55]},
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage2_19[13],stage2_18[20],stage2_17[26],stage2_16[59],stage2_15[88]}
   );
   gpc615_5 gpc2541 (
      {stage1_15[113], stage1_15[114], stage1_15[115], stage1_15[116], stage1_15[117]},
      {stage1_16[56]},
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage2_19[14],stage2_18[21],stage2_17[27],stage2_16[60],stage2_15[89]}
   );
   gpc615_5 gpc2542 (
      {stage1_15[118], stage1_15[119], stage1_15[120], stage1_15[121], stage1_15[122]},
      {stage1_16[57]},
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage2_19[15],stage2_18[22],stage2_17[28],stage2_16[61],stage2_15[90]}
   );
   gpc615_5 gpc2543 (
      {stage1_15[123], stage1_15[124], stage1_15[125], stage1_15[126], stage1_15[127]},
      {stage1_16[58]},
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage2_19[16],stage2_18[23],stage2_17[29],stage2_16[62],stage2_15[91]}
   );
   gpc606_5 gpc2544 (
      {stage1_16[59], stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[17],stage2_18[24],stage2_17[30],stage2_16[63]}
   );
   gpc606_5 gpc2545 (
      {stage1_16[65], stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[18],stage2_18[25],stage2_17[31],stage2_16[64]}
   );
   gpc606_5 gpc2546 (
      {stage1_16[71], stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[19],stage2_18[26],stage2_17[32],stage2_16[65]}
   );
   gpc606_5 gpc2547 (
      {stage1_16[77], stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[20],stage2_18[27],stage2_17[33],stage2_16[66]}
   );
   gpc606_5 gpc2548 (
      {stage1_16[83], stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[21],stage2_18[28],stage2_17[34],stage2_16[67]}
   );
   gpc606_5 gpc2549 (
      {stage1_16[89], stage1_16[90], stage1_16[91], stage1_16[92], stage1_16[93], stage1_16[94]},
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage2_20[5],stage2_19[22],stage2_18[29],stage2_17[35],stage2_16[68]}
   );
   gpc606_5 gpc2550 (
      {stage1_16[95], stage1_16[96], stage1_16[97], stage1_16[98], stage1_16[99], stage1_16[100]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage2_20[6],stage2_19[23],stage2_18[30],stage2_17[36],stage2_16[69]}
   );
   gpc606_5 gpc2551 (
      {stage1_16[101], stage1_16[102], stage1_16[103], stage1_16[104], stage1_16[105], stage1_16[106]},
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage2_20[7],stage2_19[24],stage2_18[31],stage2_17[37],stage2_16[70]}
   );
   gpc606_5 gpc2552 (
      {stage1_16[107], stage1_16[108], stage1_16[109], stage1_16[110], stage1_16[111], stage1_16[112]},
      {stage1_18[48], stage1_18[49], stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53]},
      {stage2_20[8],stage2_19[25],stage2_18[32],stage2_17[38],stage2_16[71]}
   );
   gpc606_5 gpc2553 (
      {stage1_16[113], stage1_16[114], stage1_16[115], stage1_16[116], stage1_16[117], stage1_16[118]},
      {stage1_18[54], stage1_18[55], stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59]},
      {stage2_20[9],stage2_19[26],stage2_18[33],stage2_17[39],stage2_16[72]}
   );
   gpc606_5 gpc2554 (
      {stage1_16[119], stage1_16[120], stage1_16[121], stage1_16[122], stage1_16[123], stage1_16[124]},
      {stage1_18[60], stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage2_20[10],stage2_19[27],stage2_18[34],stage2_17[40],stage2_16[73]}
   );
   gpc606_5 gpc2555 (
      {stage1_16[125], stage1_16[126], stage1_16[127], stage1_16[128], stage1_16[129], stage1_16[130]},
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70], stage1_18[71]},
      {stage2_20[11],stage2_19[28],stage2_18[35],stage2_17[41],stage2_16[74]}
   );
   gpc606_5 gpc2556 (
      {stage1_16[131], stage1_16[132], stage1_16[133], stage1_16[134], stage1_16[135], stage1_16[136]},
      {stage1_18[72], stage1_18[73], stage1_18[74], stage1_18[75], stage1_18[76], stage1_18[77]},
      {stage2_20[12],stage2_19[29],stage2_18[36],stage2_17[42],stage2_16[75]}
   );
   gpc606_5 gpc2557 (
      {stage1_16[137], stage1_16[138], stage1_16[139], stage1_16[140], stage1_16[141], stage1_16[142]},
      {stage1_18[78], stage1_18[79], stage1_18[80], stage1_18[81], stage1_18[82], stage1_18[83]},
      {stage2_20[13],stage2_19[30],stage2_18[37],stage2_17[43],stage2_16[76]}
   );
   gpc606_5 gpc2558 (
      {stage1_16[143], stage1_16[144], stage1_16[145], stage1_16[146], stage1_16[147], stage1_16[148]},
      {stage1_18[84], stage1_18[85], stage1_18[86], stage1_18[87], stage1_18[88], stage1_18[89]},
      {stage2_20[14],stage2_19[31],stage2_18[38],stage2_17[44],stage2_16[77]}
   );
   gpc606_5 gpc2559 (
      {stage1_16[149], stage1_16[150], stage1_16[151], stage1_16[152], stage1_16[153], stage1_16[154]},
      {stage1_18[90], stage1_18[91], stage1_18[92], stage1_18[93], stage1_18[94], stage1_18[95]},
      {stage2_20[15],stage2_19[32],stage2_18[39],stage2_17[45],stage2_16[78]}
   );
   gpc606_5 gpc2560 (
      {stage1_16[155], stage1_16[156], stage1_16[157], stage1_16[158], stage1_16[159], stage1_16[160]},
      {stage1_18[96], stage1_18[97], stage1_18[98], stage1_18[99], stage1_18[100], stage1_18[101]},
      {stage2_20[16],stage2_19[33],stage2_18[40],stage2_17[46],stage2_16[79]}
   );
   gpc606_5 gpc2561 (
      {stage1_16[161], stage1_16[162], stage1_16[163], stage1_16[164], stage1_16[165], stage1_16[166]},
      {stage1_18[102], stage1_18[103], stage1_18[104], stage1_18[105], stage1_18[106], stage1_18[107]},
      {stage2_20[17],stage2_19[34],stage2_18[41],stage2_17[47],stage2_16[80]}
   );
   gpc606_5 gpc2562 (
      {stage1_16[167], stage1_16[168], stage1_16[169], stage1_16[170], stage1_16[171], stage1_16[172]},
      {stage1_18[108], stage1_18[109], stage1_18[110], stage1_18[111], stage1_18[112], stage1_18[113]},
      {stage2_20[18],stage2_19[35],stage2_18[42],stage2_17[48],stage2_16[81]}
   );
   gpc606_5 gpc2563 (
      {stage1_16[173], stage1_16[174], stage1_16[175], stage1_16[176], stage1_16[177], stage1_16[178]},
      {stage1_18[114], stage1_18[115], stage1_18[116], stage1_18[117], stage1_18[118], stage1_18[119]},
      {stage2_20[19],stage2_19[36],stage2_18[43],stage2_17[49],stage2_16[82]}
   );
   gpc606_5 gpc2564 (
      {stage1_16[179], stage1_16[180], stage1_16[181], stage1_16[182], stage1_16[183], stage1_16[184]},
      {stage1_18[120], stage1_18[121], stage1_18[122], stage1_18[123], stage1_18[124], stage1_18[125]},
      {stage2_20[20],stage2_19[37],stage2_18[44],stage2_17[50],stage2_16[83]}
   );
   gpc606_5 gpc2565 (
      {stage1_16[185], stage1_16[186], stage1_16[187], stage1_16[188], stage1_16[189], stage1_16[190]},
      {stage1_18[126], stage1_18[127], stage1_18[128], stage1_18[129], stage1_18[130], stage1_18[131]},
      {stage2_20[21],stage2_19[38],stage2_18[45],stage2_17[51],stage2_16[84]}
   );
   gpc606_5 gpc2566 (
      {stage1_16[191], stage1_16[192], stage1_16[193], stage1_16[194], stage1_16[195], stage1_16[196]},
      {stage1_18[132], stage1_18[133], stage1_18[134], stage1_18[135], stage1_18[136], stage1_18[137]},
      {stage2_20[22],stage2_19[39],stage2_18[46],stage2_17[52],stage2_16[85]}
   );
   gpc606_5 gpc2567 (
      {stage1_16[197], stage1_16[198], stage1_16[199], stage1_16[200], stage1_16[201], stage1_16[202]},
      {stage1_18[138], stage1_18[139], stage1_18[140], stage1_18[141], stage1_18[142], stage1_18[143]},
      {stage2_20[23],stage2_19[40],stage2_18[47],stage2_17[53],stage2_16[86]}
   );
   gpc606_5 gpc2568 (
      {stage1_16[203], stage1_16[204], stage1_16[205], stage1_16[206], stage1_16[207], stage1_16[208]},
      {stage1_18[144], stage1_18[145], stage1_18[146], stage1_18[147], stage1_18[148], stage1_18[149]},
      {stage2_20[24],stage2_19[41],stage2_18[48],stage2_17[54],stage2_16[87]}
   );
   gpc606_5 gpc2569 (
      {stage1_16[209], stage1_16[210], stage1_16[211], stage1_16[212], stage1_16[213], stage1_16[214]},
      {stage1_18[150], stage1_18[151], stage1_18[152], stage1_18[153], stage1_18[154], stage1_18[155]},
      {stage2_20[25],stage2_19[42],stage2_18[49],stage2_17[55],stage2_16[88]}
   );
   gpc606_5 gpc2570 (
      {stage1_16[215], stage1_16[216], stage1_16[217], stage1_16[218], stage1_16[219], stage1_16[220]},
      {stage1_18[156], stage1_18[157], stage1_18[158], stage1_18[159], stage1_18[160], stage1_18[161]},
      {stage2_20[26],stage2_19[43],stage2_18[50],stage2_17[56],stage2_16[89]}
   );
   gpc606_5 gpc2571 (
      {stage1_16[221], stage1_16[222], stage1_16[223], stage1_16[224], stage1_16[225], stage1_16[226]},
      {stage1_18[162], stage1_18[163], stage1_18[164], stage1_18[165], stage1_18[166], stage1_18[167]},
      {stage2_20[27],stage2_19[44],stage2_18[51],stage2_17[57],stage2_16[90]}
   );
   gpc606_5 gpc2572 (
      {stage1_16[227], stage1_16[228], stage1_16[229], stage1_16[230], stage1_16[231], stage1_16[232]},
      {stage1_18[168], stage1_18[169], stage1_18[170], stage1_18[171], stage1_18[172], stage1_18[173]},
      {stage2_20[28],stage2_19[45],stage2_18[52],stage2_17[58],stage2_16[91]}
   );
   gpc606_5 gpc2573 (
      {stage1_16[233], stage1_16[234], stage1_16[235], stage1_16[236], stage1_16[237], stage1_16[238]},
      {stage1_18[174], stage1_18[175], stage1_18[176], stage1_18[177], stage1_18[178], stage1_18[179]},
      {stage2_20[29],stage2_19[46],stage2_18[53],stage2_17[59],stage2_16[92]}
   );
   gpc606_5 gpc2574 (
      {stage1_16[239], stage1_16[240], stage1_16[241], stage1_16[242], stage1_16[243], stage1_16[244]},
      {stage1_18[180], stage1_18[181], stage1_18[182], stage1_18[183], stage1_18[184], stage1_18[185]},
      {stage2_20[30],stage2_19[47],stage2_18[54],stage2_17[60],stage2_16[93]}
   );
   gpc606_5 gpc2575 (
      {stage1_16[245], stage1_16[246], stage1_16[247], stage1_16[248], stage1_16[249], stage1_16[250]},
      {stage1_18[186], stage1_18[187], stage1_18[188], stage1_18[189], stage1_18[190], stage1_18[191]},
      {stage2_20[31],stage2_19[48],stage2_18[55],stage2_17[61],stage2_16[94]}
   );
   gpc606_5 gpc2576 (
      {stage1_16[251], stage1_16[252], stage1_16[253], stage1_16[254], stage1_16[255], stage1_16[256]},
      {stage1_18[192], stage1_18[193], stage1_18[194], stage1_18[195], stage1_18[196], stage1_18[197]},
      {stage2_20[32],stage2_19[49],stage2_18[56],stage2_17[62],stage2_16[95]}
   );
   gpc606_5 gpc2577 (
      {stage1_17[102], stage1_17[103], stage1_17[104], stage1_17[105], stage1_17[106], stage1_17[107]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[33],stage2_19[50],stage2_18[57],stage2_17[63]}
   );
   gpc606_5 gpc2578 (
      {stage1_17[108], stage1_17[109], stage1_17[110], stage1_17[111], stage1_17[112], stage1_17[113]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[34],stage2_19[51],stage2_18[58],stage2_17[64]}
   );
   gpc606_5 gpc2579 (
      {stage1_17[114], stage1_17[115], stage1_17[116], stage1_17[117], stage1_17[118], stage1_17[119]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[35],stage2_19[52],stage2_18[59],stage2_17[65]}
   );
   gpc606_5 gpc2580 (
      {stage1_17[120], stage1_17[121], stage1_17[122], stage1_17[123], stage1_17[124], stage1_17[125]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[36],stage2_19[53],stage2_18[60],stage2_17[66]}
   );
   gpc606_5 gpc2581 (
      {stage1_17[126], stage1_17[127], stage1_17[128], stage1_17[129], stage1_17[130], stage1_17[131]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[37],stage2_19[54],stage2_18[61],stage2_17[67]}
   );
   gpc606_5 gpc2582 (
      {stage1_17[132], stage1_17[133], stage1_17[134], stage1_17[135], stage1_17[136], stage1_17[137]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[38],stage2_19[55],stage2_18[62],stage2_17[68]}
   );
   gpc606_5 gpc2583 (
      {stage1_17[138], stage1_17[139], stage1_17[140], stage1_17[141], stage1_17[142], stage1_17[143]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[39],stage2_19[56],stage2_18[63],stage2_17[69]}
   );
   gpc606_5 gpc2584 (
      {stage1_17[144], stage1_17[145], stage1_17[146], stage1_17[147], stage1_17[148], stage1_17[149]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[40],stage2_19[57],stage2_18[64],stage2_17[70]}
   );
   gpc606_5 gpc2585 (
      {stage1_17[150], stage1_17[151], stage1_17[152], stage1_17[153], stage1_17[154], stage1_17[155]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[41],stage2_19[58],stage2_18[65],stage2_17[71]}
   );
   gpc606_5 gpc2586 (
      {stage1_17[156], stage1_17[157], stage1_17[158], stage1_17[159], stage1_17[160], stage1_17[161]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[42],stage2_19[59],stage2_18[66],stage2_17[72]}
   );
   gpc606_5 gpc2587 (
      {stage1_17[162], stage1_17[163], stage1_17[164], stage1_17[165], stage1_17[166], stage1_17[167]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[43],stage2_19[60],stage2_18[67],stage2_17[73]}
   );
   gpc606_5 gpc2588 (
      {stage1_17[168], stage1_17[169], stage1_17[170], stage1_17[171], stage1_17[172], stage1_17[173]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[44],stage2_19[61],stage2_18[68],stage2_17[74]}
   );
   gpc606_5 gpc2589 (
      {stage1_17[174], stage1_17[175], stage1_17[176], stage1_17[177], stage1_17[178], stage1_17[179]},
      {stage1_19[72], stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage2_21[12],stage2_20[45],stage2_19[62],stage2_18[69],stage2_17[75]}
   );
   gpc606_5 gpc2590 (
      {stage1_17[180], stage1_17[181], stage1_17[182], stage1_17[183], stage1_17[184], stage1_17[185]},
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82], stage1_19[83]},
      {stage2_21[13],stage2_20[46],stage2_19[63],stage2_18[70],stage2_17[76]}
   );
   gpc606_5 gpc2591 (
      {stage1_17[186], stage1_17[187], stage1_17[188], stage1_17[189], stage1_17[190], stage1_17[191]},
      {stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87], stage1_19[88], stage1_19[89]},
      {stage2_21[14],stage2_20[47],stage2_19[64],stage2_18[71],stage2_17[77]}
   );
   gpc606_5 gpc2592 (
      {stage1_17[192], stage1_17[193], stage1_17[194], stage1_17[195], stage1_17[196], stage1_17[197]},
      {stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93], stage1_19[94], stage1_19[95]},
      {stage2_21[15],stage2_20[48],stage2_19[65],stage2_18[72],stage2_17[78]}
   );
   gpc606_5 gpc2593 (
      {stage1_17[198], stage1_17[199], stage1_17[200], stage1_17[201], stage1_17[202], stage1_17[203]},
      {stage1_19[96], stage1_19[97], stage1_19[98], stage1_19[99], stage1_19[100], stage1_19[101]},
      {stage2_21[16],stage2_20[49],stage2_19[66],stage2_18[73],stage2_17[79]}
   );
   gpc606_5 gpc2594 (
      {stage1_17[204], stage1_17[205], stage1_17[206], stage1_17[207], stage1_17[208], stage1_17[209]},
      {stage1_19[102], stage1_19[103], stage1_19[104], stage1_19[105], stage1_19[106], stage1_19[107]},
      {stage2_21[17],stage2_20[50],stage2_19[67],stage2_18[74],stage2_17[80]}
   );
   gpc606_5 gpc2595 (
      {stage1_17[210], stage1_17[211], stage1_17[212], stage1_17[213], stage1_17[214], stage1_17[215]},
      {stage1_19[108], stage1_19[109], stage1_19[110], stage1_19[111], stage1_19[112], stage1_19[113]},
      {stage2_21[18],stage2_20[51],stage2_19[68],stage2_18[75],stage2_17[81]}
   );
   gpc606_5 gpc2596 (
      {stage1_17[216], stage1_17[217], stage1_17[218], stage1_17[219], stage1_17[220], stage1_17[221]},
      {stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117], stage1_19[118], stage1_19[119]},
      {stage2_21[19],stage2_20[52],stage2_19[69],stage2_18[76],stage2_17[82]}
   );
   gpc606_5 gpc2597 (
      {stage1_17[222], stage1_17[223], stage1_17[224], stage1_17[225], stage1_17[226], stage1_17[227]},
      {stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123], stage1_19[124], stage1_19[125]},
      {stage2_21[20],stage2_20[53],stage2_19[70],stage2_18[77],stage2_17[83]}
   );
   gpc606_5 gpc2598 (
      {stage1_17[228], stage1_17[229], stage1_17[230], stage1_17[231], stage1_17[232], stage1_17[233]},
      {stage1_19[126], stage1_19[127], stage1_19[128], stage1_19[129], stage1_19[130], stage1_19[131]},
      {stage2_21[21],stage2_20[54],stage2_19[71],stage2_18[78],stage2_17[84]}
   );
   gpc615_5 gpc2599 (
      {stage1_19[132], stage1_19[133], stage1_19[134], stage1_19[135], stage1_19[136]},
      {stage1_20[0]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[0],stage2_21[22],stage2_20[55],stage2_19[72]}
   );
   gpc615_5 gpc2600 (
      {stage1_19[137], stage1_19[138], stage1_19[139], stage1_19[140], stage1_19[141]},
      {stage1_20[1]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[1],stage2_21[23],stage2_20[56],stage2_19[73]}
   );
   gpc615_5 gpc2601 (
      {stage1_19[142], stage1_19[143], stage1_19[144], stage1_19[145], stage1_19[146]},
      {stage1_20[2]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[2],stage2_21[24],stage2_20[57],stage2_19[74]}
   );
   gpc615_5 gpc2602 (
      {stage1_19[147], stage1_19[148], stage1_19[149], stage1_19[150], stage1_19[151]},
      {stage1_20[3]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[3],stage2_21[25],stage2_20[58],stage2_19[75]}
   );
   gpc615_5 gpc2603 (
      {stage1_19[152], stage1_19[153], stage1_19[154], stage1_19[155], stage1_19[156]},
      {stage1_20[4]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[4],stage2_21[26],stage2_20[59],stage2_19[76]}
   );
   gpc615_5 gpc2604 (
      {stage1_19[157], stage1_19[158], stage1_19[159], stage1_19[160], stage1_19[161]},
      {stage1_20[5]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[5],stage2_21[27],stage2_20[60],stage2_19[77]}
   );
   gpc615_5 gpc2605 (
      {stage1_19[162], stage1_19[163], stage1_19[164], stage1_19[165], stage1_19[166]},
      {stage1_20[6]},
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage2_23[6],stage2_22[6],stage2_21[28],stage2_20[61],stage2_19[78]}
   );
   gpc615_5 gpc2606 (
      {stage1_19[167], stage1_19[168], stage1_19[169], stage1_19[170], stage1_19[171]},
      {stage1_20[7]},
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage2_23[7],stage2_22[7],stage2_21[29],stage2_20[62],stage2_19[79]}
   );
   gpc615_5 gpc2607 (
      {stage1_19[172], stage1_19[173], stage1_19[174], stage1_19[175], stage1_19[176]},
      {stage1_20[8]},
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage2_23[8],stage2_22[8],stage2_21[30],stage2_20[63],stage2_19[80]}
   );
   gpc615_5 gpc2608 (
      {stage1_19[177], stage1_19[178], stage1_19[179], stage1_19[180], stage1_19[181]},
      {stage1_20[9]},
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage2_23[9],stage2_22[9],stage2_21[31],stage2_20[64],stage2_19[81]}
   );
   gpc615_5 gpc2609 (
      {stage1_19[182], stage1_19[183], stage1_19[184], stage1_19[185], stage1_19[186]},
      {stage1_20[10]},
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage2_23[10],stage2_22[10],stage2_21[32],stage2_20[65],stage2_19[82]}
   );
   gpc615_5 gpc2610 (
      {stage1_19[187], stage1_19[188], stage1_19[189], stage1_19[190], stage1_19[191]},
      {stage1_20[11]},
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage2_23[11],stage2_22[11],stage2_21[33],stage2_20[66],stage2_19[83]}
   );
   gpc615_5 gpc2611 (
      {stage1_19[192], stage1_19[193], stage1_19[194], stage1_19[195], stage1_19[196]},
      {stage1_20[12]},
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage2_23[12],stage2_22[12],stage2_21[34],stage2_20[67],stage2_19[84]}
   );
   gpc615_5 gpc2612 (
      {stage1_19[197], stage1_19[198], stage1_19[199], stage1_19[200], stage1_19[201]},
      {stage1_20[13]},
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage2_23[13],stage2_22[13],stage2_21[35],stage2_20[68],stage2_19[85]}
   );
   gpc615_5 gpc2613 (
      {stage1_19[202], stage1_19[203], stage1_19[204], stage1_19[205], stage1_19[206]},
      {stage1_20[14]},
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage2_23[14],stage2_22[14],stage2_21[36],stage2_20[69],stage2_19[86]}
   );
   gpc615_5 gpc2614 (
      {stage1_19[207], stage1_19[208], stage1_19[209], stage1_19[210], stage1_19[211]},
      {stage1_20[15]},
      {stage1_21[90], stage1_21[91], stage1_21[92], stage1_21[93], stage1_21[94], stage1_21[95]},
      {stage2_23[15],stage2_22[15],stage2_21[37],stage2_20[70],stage2_19[87]}
   );
   gpc615_5 gpc2615 (
      {stage1_19[212], stage1_19[213], stage1_19[214], stage1_19[215], stage1_19[216]},
      {stage1_20[16]},
      {stage1_21[96], stage1_21[97], stage1_21[98], stage1_21[99], stage1_21[100], stage1_21[101]},
      {stage2_23[16],stage2_22[16],stage2_21[38],stage2_20[71],stage2_19[88]}
   );
   gpc615_5 gpc2616 (
      {stage1_19[217], stage1_19[218], stage1_19[219], stage1_19[220], stage1_19[221]},
      {stage1_20[17]},
      {stage1_21[102], stage1_21[103], stage1_21[104], stage1_21[105], stage1_21[106], stage1_21[107]},
      {stage2_23[17],stage2_22[17],stage2_21[39],stage2_20[72],stage2_19[89]}
   );
   gpc615_5 gpc2617 (
      {stage1_19[222], stage1_19[223], stage1_19[224], stage1_19[225], stage1_19[226]},
      {stage1_20[18]},
      {stage1_21[108], stage1_21[109], stage1_21[110], stage1_21[111], stage1_21[112], stage1_21[113]},
      {stage2_23[18],stage2_22[18],stage2_21[40],stage2_20[73],stage2_19[90]}
   );
   gpc615_5 gpc2618 (
      {stage1_19[227], stage1_19[228], stage1_19[229], stage1_19[230], stage1_19[231]},
      {stage1_20[19]},
      {stage1_21[114], stage1_21[115], stage1_21[116], stage1_21[117], stage1_21[118], stage1_21[119]},
      {stage2_23[19],stage2_22[19],stage2_21[41],stage2_20[74],stage2_19[91]}
   );
   gpc615_5 gpc2619 (
      {stage1_19[232], stage1_19[233], stage1_19[234], stage1_19[235], stage1_19[236]},
      {stage1_20[20]},
      {stage1_21[120], stage1_21[121], stage1_21[122], stage1_21[123], stage1_21[124], stage1_21[125]},
      {stage2_23[20],stage2_22[20],stage2_21[42],stage2_20[75],stage2_19[92]}
   );
   gpc615_5 gpc2620 (
      {stage1_19[237], stage1_19[238], stage1_19[239], stage1_19[240], stage1_19[241]},
      {stage1_20[21]},
      {stage1_21[126], stage1_21[127], stage1_21[128], stage1_21[129], stage1_21[130], stage1_21[131]},
      {stage2_23[21],stage2_22[21],stage2_21[43],stage2_20[76],stage2_19[93]}
   );
   gpc615_5 gpc2621 (
      {stage1_19[242], stage1_19[243], stage1_19[244], stage1_19[245], stage1_19[246]},
      {stage1_20[22]},
      {stage1_21[132], stage1_21[133], stage1_21[134], stage1_21[135], stage1_21[136], stage1_21[137]},
      {stage2_23[22],stage2_22[22],stage2_21[44],stage2_20[77],stage2_19[94]}
   );
   gpc615_5 gpc2622 (
      {stage1_19[247], stage1_19[248], stage1_19[249], stage1_19[250], stage1_19[251]},
      {stage1_20[23]},
      {stage1_21[138], stage1_21[139], stage1_21[140], stage1_21[141], stage1_21[142], stage1_21[143]},
      {stage2_23[23],stage2_22[23],stage2_21[45],stage2_20[78],stage2_19[95]}
   );
   gpc615_5 gpc2623 (
      {stage1_19[252], stage1_19[253], stage1_19[254], stage1_19[255], stage1_19[256]},
      {stage1_20[24]},
      {stage1_21[144], stage1_21[145], stage1_21[146], stage1_21[147], stage1_21[148], stage1_21[149]},
      {stage2_23[24],stage2_22[24],stage2_21[46],stage2_20[79],stage2_19[96]}
   );
   gpc615_5 gpc2624 (
      {stage1_19[257], stage1_19[258], stage1_19[259], stage1_19[260], stage1_19[261]},
      {stage1_20[25]},
      {stage1_21[150], stage1_21[151], stage1_21[152], stage1_21[153], stage1_21[154], stage1_21[155]},
      {stage2_23[25],stage2_22[25],stage2_21[47],stage2_20[80],stage2_19[97]}
   );
   gpc615_5 gpc2625 (
      {stage1_19[262], stage1_19[263], stage1_19[264], stage1_19[265], stage1_19[266]},
      {stage1_20[26]},
      {stage1_21[156], stage1_21[157], stage1_21[158], stage1_21[159], stage1_21[160], stage1_21[161]},
      {stage2_23[26],stage2_22[26],stage2_21[48],stage2_20[81],stage2_19[98]}
   );
   gpc615_5 gpc2626 (
      {stage1_19[267], stage1_19[268], stage1_19[269], stage1_19[270], stage1_19[271]},
      {stage1_20[27]},
      {stage1_21[162], stage1_21[163], stage1_21[164], stage1_21[165], stage1_21[166], stage1_21[167]},
      {stage2_23[27],stage2_22[27],stage2_21[49],stage2_20[82],stage2_19[99]}
   );
   gpc615_5 gpc2627 (
      {stage1_19[272], stage1_19[273], stage1_19[274], stage1_19[275], stage1_19[276]},
      {stage1_20[28]},
      {stage1_21[168], stage1_21[169], stage1_21[170], stage1_21[171], stage1_21[172], stage1_21[173]},
      {stage2_23[28],stage2_22[28],stage2_21[50],stage2_20[83],stage2_19[100]}
   );
   gpc615_5 gpc2628 (
      {stage1_19[277], stage1_19[278], stage1_19[279], stage1_19[280], stage1_19[281]},
      {stage1_20[29]},
      {stage1_21[174], stage1_21[175], stage1_21[176], stage1_21[177], stage1_21[178], stage1_21[179]},
      {stage2_23[29],stage2_22[29],stage2_21[51],stage2_20[84],stage2_19[101]}
   );
   gpc615_5 gpc2629 (
      {stage1_19[282], stage1_19[283], stage1_19[284], stage1_19[285], stage1_19[286]},
      {stage1_20[30]},
      {stage1_21[180], stage1_21[181], stage1_21[182], stage1_21[183], stage1_21[184], stage1_21[185]},
      {stage2_23[30],stage2_22[30],stage2_21[52],stage2_20[85],stage2_19[102]}
   );
   gpc615_5 gpc2630 (
      {stage1_19[287], stage1_19[288], stage1_19[289], stage1_19[290], stage1_19[291]},
      {stage1_20[31]},
      {stage1_21[186], stage1_21[187], stage1_21[188], stage1_21[189], stage1_21[190], stage1_21[191]},
      {stage2_23[31],stage2_22[31],stage2_21[53],stage2_20[86],stage2_19[103]}
   );
   gpc623_5 gpc2631 (
      {stage1_19[292], stage1_19[293], stage1_19[294]},
      {stage1_20[32], stage1_20[33]},
      {stage1_21[192], stage1_21[193], stage1_21[194], stage1_21[195], stage1_21[196], stage1_21[197]},
      {stage2_23[32],stage2_22[32],stage2_21[54],stage2_20[87],stage2_19[104]}
   );
   gpc606_5 gpc2632 (
      {stage1_20[34], stage1_20[35], stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[33],stage2_22[33],stage2_21[55],stage2_20[88]}
   );
   gpc606_5 gpc2633 (
      {stage1_20[40], stage1_20[41], stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[34],stage2_22[34],stage2_21[56],stage2_20[89]}
   );
   gpc606_5 gpc2634 (
      {stage1_20[46], stage1_20[47], stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[35],stage2_22[35],stage2_21[57],stage2_20[90]}
   );
   gpc606_5 gpc2635 (
      {stage1_20[52], stage1_20[53], stage1_20[54], stage1_20[55], stage1_20[56], stage1_20[57]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[36],stage2_22[36],stage2_21[58],stage2_20[91]}
   );
   gpc606_5 gpc2636 (
      {stage1_20[58], stage1_20[59], stage1_20[60], stage1_20[61], stage1_20[62], stage1_20[63]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[37],stage2_22[37],stage2_21[59],stage2_20[92]}
   );
   gpc606_5 gpc2637 (
      {stage1_20[64], stage1_20[65], stage1_20[66], stage1_20[67], stage1_20[68], stage1_20[69]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[38],stage2_22[38],stage2_21[60],stage2_20[93]}
   );
   gpc606_5 gpc2638 (
      {stage1_20[70], stage1_20[71], stage1_20[72], stage1_20[73], stage1_20[74], stage1_20[75]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[39],stage2_22[39],stage2_21[61],stage2_20[94]}
   );
   gpc606_5 gpc2639 (
      {stage1_20[76], stage1_20[77], stage1_20[78], stage1_20[79], stage1_20[80], stage1_20[81]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[40],stage2_22[40],stage2_21[62],stage2_20[95]}
   );
   gpc606_5 gpc2640 (
      {stage1_20[82], stage1_20[83], stage1_20[84], stage1_20[85], stage1_20[86], stage1_20[87]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[41],stage2_22[41],stage2_21[63],stage2_20[96]}
   );
   gpc606_5 gpc2641 (
      {stage1_20[88], stage1_20[89], stage1_20[90], stage1_20[91], stage1_20[92], stage1_20[93]},
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage2_24[9],stage2_23[42],stage2_22[42],stage2_21[64],stage2_20[97]}
   );
   gpc606_5 gpc2642 (
      {stage1_20[94], stage1_20[95], stage1_20[96], stage1_20[97], stage1_20[98], stage1_20[99]},
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage2_24[10],stage2_23[43],stage2_22[43],stage2_21[65],stage2_20[98]}
   );
   gpc606_5 gpc2643 (
      {stage1_20[100], stage1_20[101], stage1_20[102], stage1_20[103], stage1_20[104], stage1_20[105]},
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage2_24[11],stage2_23[44],stage2_22[44],stage2_21[66],stage2_20[99]}
   );
   gpc606_5 gpc2644 (
      {stage1_20[106], stage1_20[107], stage1_20[108], stage1_20[109], stage1_20[110], stage1_20[111]},
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76], stage1_22[77]},
      {stage2_24[12],stage2_23[45],stage2_22[45],stage2_21[67],stage2_20[100]}
   );
   gpc606_5 gpc2645 (
      {stage1_20[112], stage1_20[113], stage1_20[114], stage1_20[115], stage1_20[116], stage1_20[117]},
      {stage1_22[78], stage1_22[79], stage1_22[80], stage1_22[81], stage1_22[82], stage1_22[83]},
      {stage2_24[13],stage2_23[46],stage2_22[46],stage2_21[68],stage2_20[101]}
   );
   gpc606_5 gpc2646 (
      {stage1_20[118], stage1_20[119], stage1_20[120], stage1_20[121], stage1_20[122], stage1_20[123]},
      {stage1_22[84], stage1_22[85], stage1_22[86], stage1_22[87], stage1_22[88], stage1_22[89]},
      {stage2_24[14],stage2_23[47],stage2_22[47],stage2_21[69],stage2_20[102]}
   );
   gpc606_5 gpc2647 (
      {stage1_20[124], stage1_20[125], stage1_20[126], stage1_20[127], stage1_20[128], stage1_20[129]},
      {stage1_22[90], stage1_22[91], stage1_22[92], stage1_22[93], stage1_22[94], stage1_22[95]},
      {stage2_24[15],stage2_23[48],stage2_22[48],stage2_21[70],stage2_20[103]}
   );
   gpc606_5 gpc2648 (
      {stage1_20[130], stage1_20[131], stage1_20[132], stage1_20[133], stage1_20[134], stage1_20[135]},
      {stage1_22[96], stage1_22[97], stage1_22[98], stage1_22[99], stage1_22[100], stage1_22[101]},
      {stage2_24[16],stage2_23[49],stage2_22[49],stage2_21[71],stage2_20[104]}
   );
   gpc606_5 gpc2649 (
      {stage1_20[136], stage1_20[137], stage1_20[138], stage1_20[139], stage1_20[140], stage1_20[141]},
      {stage1_22[102], stage1_22[103], stage1_22[104], stage1_22[105], stage1_22[106], stage1_22[107]},
      {stage2_24[17],stage2_23[50],stage2_22[50],stage2_21[72],stage2_20[105]}
   );
   gpc606_5 gpc2650 (
      {stage1_20[142], stage1_20[143], stage1_20[144], stage1_20[145], stage1_20[146], stage1_20[147]},
      {stage1_22[108], stage1_22[109], stage1_22[110], stage1_22[111], stage1_22[112], stage1_22[113]},
      {stage2_24[18],stage2_23[51],stage2_22[51],stage2_21[73],stage2_20[106]}
   );
   gpc606_5 gpc2651 (
      {stage1_20[148], stage1_20[149], stage1_20[150], stage1_20[151], stage1_20[152], stage1_20[153]},
      {stage1_22[114], stage1_22[115], stage1_22[116], stage1_22[117], stage1_22[118], stage1_22[119]},
      {stage2_24[19],stage2_23[52],stage2_22[52],stage2_21[74],stage2_20[107]}
   );
   gpc606_5 gpc2652 (
      {stage1_20[154], stage1_20[155], stage1_20[156], stage1_20[157], stage1_20[158], stage1_20[159]},
      {stage1_22[120], stage1_22[121], stage1_22[122], stage1_22[123], stage1_22[124], stage1_22[125]},
      {stage2_24[20],stage2_23[53],stage2_22[53],stage2_21[75],stage2_20[108]}
   );
   gpc606_5 gpc2653 (
      {stage1_20[160], stage1_20[161], stage1_20[162], stage1_20[163], stage1_20[164], stage1_20[165]},
      {stage1_22[126], stage1_22[127], stage1_22[128], stage1_22[129], stage1_22[130], stage1_22[131]},
      {stage2_24[21],stage2_23[54],stage2_22[54],stage2_21[76],stage2_20[109]}
   );
   gpc606_5 gpc2654 (
      {stage1_20[166], stage1_20[167], stage1_20[168], stage1_20[169], stage1_20[170], stage1_20[171]},
      {stage1_22[132], stage1_22[133], stage1_22[134], stage1_22[135], stage1_22[136], stage1_22[137]},
      {stage2_24[22],stage2_23[55],stage2_22[55],stage2_21[77],stage2_20[110]}
   );
   gpc615_5 gpc2655 (
      {stage1_22[138], stage1_22[139], stage1_22[140], stage1_22[141], stage1_22[142]},
      {stage1_23[0]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[0],stage2_24[23],stage2_23[56],stage2_22[56]}
   );
   gpc615_5 gpc2656 (
      {stage1_22[143], stage1_22[144], stage1_22[145], stage1_22[146], stage1_22[147]},
      {stage1_23[1]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[1],stage2_24[24],stage2_23[57],stage2_22[57]}
   );
   gpc615_5 gpc2657 (
      {stage1_22[148], stage1_22[149], stage1_22[150], stage1_22[151], stage1_22[152]},
      {stage1_23[2]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[2],stage2_24[25],stage2_23[58],stage2_22[58]}
   );
   gpc615_5 gpc2658 (
      {stage1_22[153], stage1_22[154], stage1_22[155], stage1_22[156], stage1_22[157]},
      {stage1_23[3]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[3],stage2_24[26],stage2_23[59],stage2_22[59]}
   );
   gpc615_5 gpc2659 (
      {stage1_22[158], stage1_22[159], stage1_22[160], stage1_22[161], stage1_22[162]},
      {stage1_23[4]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[4],stage2_24[27],stage2_23[60],stage2_22[60]}
   );
   gpc615_5 gpc2660 (
      {stage1_22[163], stage1_22[164], stage1_22[165], stage1_22[166], stage1_22[167]},
      {stage1_23[5]},
      {stage1_24[30], stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35]},
      {stage2_26[5],stage2_25[5],stage2_24[28],stage2_23[61],stage2_22[61]}
   );
   gpc615_5 gpc2661 (
      {stage1_22[168], stage1_22[169], stage1_22[170], stage1_22[171], stage1_22[172]},
      {stage1_23[6]},
      {stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41]},
      {stage2_26[6],stage2_25[6],stage2_24[29],stage2_23[62],stage2_22[62]}
   );
   gpc615_5 gpc2662 (
      {stage1_22[173], stage1_22[174], stage1_22[175], stage1_22[176], stage1_22[177]},
      {stage1_23[7]},
      {stage1_24[42], stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47]},
      {stage2_26[7],stage2_25[7],stage2_24[30],stage2_23[63],stage2_22[63]}
   );
   gpc615_5 gpc2663 (
      {stage1_22[178], stage1_22[179], stage1_22[180], stage1_22[181], stage1_22[182]},
      {stage1_23[8]},
      {stage1_24[48], stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage2_26[8],stage2_25[8],stage2_24[31],stage2_23[64],stage2_22[64]}
   );
   gpc615_5 gpc2664 (
      {stage1_22[183], stage1_22[184], stage1_22[185], stage1_22[186], stage1_22[187]},
      {stage1_23[9]},
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage2_26[9],stage2_25[9],stage2_24[32],stage2_23[65],stage2_22[65]}
   );
   gpc615_5 gpc2665 (
      {stage1_22[188], stage1_22[189], stage1_22[190], stage1_22[191], stage1_22[192]},
      {stage1_23[10]},
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65]},
      {stage2_26[10],stage2_25[10],stage2_24[33],stage2_23[66],stage2_22[66]}
   );
   gpc615_5 gpc2666 (
      {stage1_22[193], stage1_22[194], stage1_22[195], stage1_22[196], stage1_22[197]},
      {stage1_23[11]},
      {stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71]},
      {stage2_26[11],stage2_25[11],stage2_24[34],stage2_23[67],stage2_22[67]}
   );
   gpc615_5 gpc2667 (
      {stage1_22[198], stage1_22[199], stage1_22[200], stage1_22[201], stage1_22[202]},
      {stage1_23[12]},
      {stage1_24[72], stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77]},
      {stage2_26[12],stage2_25[12],stage2_24[35],stage2_23[68],stage2_22[68]}
   );
   gpc615_5 gpc2668 (
      {stage1_22[203], stage1_22[204], stage1_22[205], stage1_22[206], stage1_22[207]},
      {stage1_23[13]},
      {stage1_24[78], stage1_24[79], stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83]},
      {stage2_26[13],stage2_25[13],stage2_24[36],stage2_23[69],stage2_22[69]}
   );
   gpc615_5 gpc2669 (
      {stage1_22[208], stage1_22[209], stage1_22[210], stage1_22[211], stage1_22[212]},
      {stage1_23[14]},
      {stage1_24[84], stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage2_26[14],stage2_25[14],stage2_24[37],stage2_23[70],stage2_22[70]}
   );
   gpc615_5 gpc2670 (
      {stage1_22[213], stage1_22[214], stage1_22[215], stage1_22[216], stage1_22[217]},
      {stage1_23[15]},
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94], stage1_24[95]},
      {stage2_26[15],stage2_25[15],stage2_24[38],stage2_23[71],stage2_22[71]}
   );
   gpc615_5 gpc2671 (
      {stage1_22[218], stage1_22[219], stage1_22[220], stage1_22[221], stage1_22[222]},
      {stage1_23[16]},
      {stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99], stage1_24[100], stage1_24[101]},
      {stage2_26[16],stage2_25[16],stage2_24[39],stage2_23[72],stage2_22[72]}
   );
   gpc615_5 gpc2672 (
      {stage1_22[223], stage1_22[224], stage1_22[225], stage1_22[226], stage1_22[227]},
      {stage1_23[17]},
      {stage1_24[102], stage1_24[103], stage1_24[104], stage1_24[105], stage1_24[106], stage1_24[107]},
      {stage2_26[17],stage2_25[17],stage2_24[40],stage2_23[73],stage2_22[73]}
   );
   gpc615_5 gpc2673 (
      {stage1_22[228], stage1_22[229], stage1_22[230], stage1_22[231], stage1_22[232]},
      {stage1_23[18]},
      {stage1_24[108], stage1_24[109], stage1_24[110], stage1_24[111], stage1_24[112], stage1_24[113]},
      {stage2_26[18],stage2_25[18],stage2_24[41],stage2_23[74],stage2_22[74]}
   );
   gpc615_5 gpc2674 (
      {stage1_22[233], stage1_22[234], stage1_22[235], stage1_22[236], stage1_22[237]},
      {stage1_23[19]},
      {stage1_24[114], stage1_24[115], stage1_24[116], stage1_24[117], stage1_24[118], stage1_24[119]},
      {stage2_26[19],stage2_25[19],stage2_24[42],stage2_23[75],stage2_22[75]}
   );
   gpc615_5 gpc2675 (
      {stage1_22[238], stage1_22[239], stage1_22[240], stage1_22[241], stage1_22[242]},
      {stage1_23[20]},
      {stage1_24[120], stage1_24[121], stage1_24[122], stage1_24[123], stage1_24[124], stage1_24[125]},
      {stage2_26[20],stage2_25[20],stage2_24[43],stage2_23[76],stage2_22[76]}
   );
   gpc615_5 gpc2676 (
      {stage1_22[243], stage1_22[244], stage1_22[245], stage1_22[246], stage1_22[247]},
      {stage1_23[21]},
      {stage1_24[126], stage1_24[127], stage1_24[128], stage1_24[129], stage1_24[130], stage1_24[131]},
      {stage2_26[21],stage2_25[21],stage2_24[44],stage2_23[77],stage2_22[77]}
   );
   gpc615_5 gpc2677 (
      {stage1_22[248], stage1_22[249], stage1_22[250], 1'b0, 1'b0},
      {stage1_23[22]},
      {stage1_24[132], stage1_24[133], stage1_24[134], stage1_24[135], stage1_24[136], stage1_24[137]},
      {stage2_26[22],stage2_25[22],stage2_24[45],stage2_23[78],stage2_22[78]}
   );
   gpc615_5 gpc2678 (
      {stage1_23[23], stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27]},
      {stage1_24[138]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[23],stage2_25[23],stage2_24[46],stage2_23[79]}
   );
   gpc615_5 gpc2679 (
      {stage1_23[28], stage1_23[29], stage1_23[30], stage1_23[31], stage1_23[32]},
      {stage1_24[139]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[24],stage2_25[24],stage2_24[47],stage2_23[80]}
   );
   gpc615_5 gpc2680 (
      {stage1_23[33], stage1_23[34], stage1_23[35], stage1_23[36], stage1_23[37]},
      {stage1_24[140]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[25],stage2_25[25],stage2_24[48],stage2_23[81]}
   );
   gpc615_5 gpc2681 (
      {stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41], stage1_23[42]},
      {stage1_24[141]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[26],stage2_25[26],stage2_24[49],stage2_23[82]}
   );
   gpc615_5 gpc2682 (
      {stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage1_24[142]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[27],stage2_25[27],stage2_24[50],stage2_23[83]}
   );
   gpc615_5 gpc2683 (
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52]},
      {stage1_24[143]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[28],stage2_25[28],stage2_24[51],stage2_23[84]}
   );
   gpc615_5 gpc2684 (
      {stage1_23[53], stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57]},
      {stage1_24[144]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[29],stage2_25[29],stage2_24[52],stage2_23[85]}
   );
   gpc615_5 gpc2685 (
      {stage1_23[58], stage1_23[59], stage1_23[60], stage1_23[61], stage1_23[62]},
      {stage1_24[145]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[30],stage2_25[30],stage2_24[53],stage2_23[86]}
   );
   gpc615_5 gpc2686 (
      {stage1_23[63], stage1_23[64], stage1_23[65], stage1_23[66], stage1_23[67]},
      {stage1_24[146]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage2_27[8],stage2_26[31],stage2_25[31],stage2_24[54],stage2_23[87]}
   );
   gpc615_5 gpc2687 (
      {stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71], stage1_23[72]},
      {stage1_24[147]},
      {stage1_25[54], stage1_25[55], stage1_25[56], stage1_25[57], stage1_25[58], stage1_25[59]},
      {stage2_27[9],stage2_26[32],stage2_25[32],stage2_24[55],stage2_23[88]}
   );
   gpc615_5 gpc2688 (
      {stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage1_24[148]},
      {stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64], stage1_25[65]},
      {stage2_27[10],stage2_26[33],stage2_25[33],stage2_24[56],stage2_23[89]}
   );
   gpc615_5 gpc2689 (
      {stage1_23[78], stage1_23[79], stage1_23[80], stage1_23[81], stage1_23[82]},
      {stage1_24[149]},
      {stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70], stage1_25[71]},
      {stage2_27[11],stage2_26[34],stage2_25[34],stage2_24[57],stage2_23[90]}
   );
   gpc615_5 gpc2690 (
      {stage1_23[83], stage1_23[84], stage1_23[85], stage1_23[86], stage1_23[87]},
      {stage1_24[150]},
      {stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76], stage1_25[77]},
      {stage2_27[12],stage2_26[35],stage2_25[35],stage2_24[58],stage2_23[91]}
   );
   gpc615_5 gpc2691 (
      {stage1_23[88], stage1_23[89], stage1_23[90], stage1_23[91], stage1_23[92]},
      {stage1_24[151]},
      {stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82], stage1_25[83]},
      {stage2_27[13],stage2_26[36],stage2_25[36],stage2_24[59],stage2_23[92]}
   );
   gpc615_5 gpc2692 (
      {stage1_23[93], stage1_23[94], stage1_23[95], stage1_23[96], stage1_23[97]},
      {stage1_24[152]},
      {stage1_25[84], stage1_25[85], stage1_25[86], stage1_25[87], stage1_25[88], stage1_25[89]},
      {stage2_27[14],stage2_26[37],stage2_25[37],stage2_24[60],stage2_23[93]}
   );
   gpc615_5 gpc2693 (
      {stage1_23[98], stage1_23[99], stage1_23[100], stage1_23[101], stage1_23[102]},
      {stage1_24[153]},
      {stage1_25[90], stage1_25[91], stage1_25[92], stage1_25[93], stage1_25[94], stage1_25[95]},
      {stage2_27[15],stage2_26[38],stage2_25[38],stage2_24[61],stage2_23[94]}
   );
   gpc615_5 gpc2694 (
      {stage1_23[103], stage1_23[104], stage1_23[105], stage1_23[106], stage1_23[107]},
      {stage1_24[154]},
      {stage1_25[96], stage1_25[97], stage1_25[98], stage1_25[99], stage1_25[100], stage1_25[101]},
      {stage2_27[16],stage2_26[39],stage2_25[39],stage2_24[62],stage2_23[95]}
   );
   gpc615_5 gpc2695 (
      {stage1_23[108], stage1_23[109], stage1_23[110], stage1_23[111], stage1_23[112]},
      {stage1_24[155]},
      {stage1_25[102], stage1_25[103], stage1_25[104], stage1_25[105], stage1_25[106], stage1_25[107]},
      {stage2_27[17],stage2_26[40],stage2_25[40],stage2_24[63],stage2_23[96]}
   );
   gpc615_5 gpc2696 (
      {stage1_23[113], stage1_23[114], stage1_23[115], stage1_23[116], stage1_23[117]},
      {stage1_24[156]},
      {stage1_25[108], stage1_25[109], stage1_25[110], stage1_25[111], stage1_25[112], stage1_25[113]},
      {stage2_27[18],stage2_26[41],stage2_25[41],stage2_24[64],stage2_23[97]}
   );
   gpc615_5 gpc2697 (
      {stage1_23[118], stage1_23[119], stage1_23[120], stage1_23[121], stage1_23[122]},
      {stage1_24[157]},
      {stage1_25[114], stage1_25[115], stage1_25[116], stage1_25[117], stage1_25[118], stage1_25[119]},
      {stage2_27[19],stage2_26[42],stage2_25[42],stage2_24[65],stage2_23[98]}
   );
   gpc615_5 gpc2698 (
      {stage1_23[123], stage1_23[124], stage1_23[125], stage1_23[126], stage1_23[127]},
      {stage1_24[158]},
      {stage1_25[120], stage1_25[121], stage1_25[122], stage1_25[123], stage1_25[124], stage1_25[125]},
      {stage2_27[20],stage2_26[43],stage2_25[43],stage2_24[66],stage2_23[99]}
   );
   gpc615_5 gpc2699 (
      {stage1_23[128], stage1_23[129], stage1_23[130], stage1_23[131], stage1_23[132]},
      {stage1_24[159]},
      {stage1_25[126], stage1_25[127], stage1_25[128], stage1_25[129], stage1_25[130], stage1_25[131]},
      {stage2_27[21],stage2_26[44],stage2_25[44],stage2_24[67],stage2_23[100]}
   );
   gpc615_5 gpc2700 (
      {stage1_23[133], stage1_23[134], stage1_23[135], stage1_23[136], stage1_23[137]},
      {stage1_24[160]},
      {stage1_25[132], stage1_25[133], stage1_25[134], stage1_25[135], stage1_25[136], stage1_25[137]},
      {stage2_27[22],stage2_26[45],stage2_25[45],stage2_24[68],stage2_23[101]}
   );
   gpc615_5 gpc2701 (
      {stage1_23[138], stage1_23[139], stage1_23[140], stage1_23[141], stage1_23[142]},
      {stage1_24[161]},
      {stage1_25[138], stage1_25[139], stage1_25[140], stage1_25[141], stage1_25[142], stage1_25[143]},
      {stage2_27[23],stage2_26[46],stage2_25[46],stage2_24[69],stage2_23[102]}
   );
   gpc615_5 gpc2702 (
      {stage1_23[143], stage1_23[144], stage1_23[145], stage1_23[146], stage1_23[147]},
      {stage1_24[162]},
      {stage1_25[144], stage1_25[145], stage1_25[146], stage1_25[147], stage1_25[148], stage1_25[149]},
      {stage2_27[24],stage2_26[47],stage2_25[47],stage2_24[70],stage2_23[103]}
   );
   gpc615_5 gpc2703 (
      {stage1_23[148], stage1_23[149], stage1_23[150], stage1_23[151], stage1_23[152]},
      {stage1_24[163]},
      {stage1_25[150], stage1_25[151], stage1_25[152], stage1_25[153], stage1_25[154], stage1_25[155]},
      {stage2_27[25],stage2_26[48],stage2_25[48],stage2_24[71],stage2_23[104]}
   );
   gpc615_5 gpc2704 (
      {stage1_23[153], stage1_23[154], stage1_23[155], stage1_23[156], stage1_23[157]},
      {stage1_24[164]},
      {stage1_25[156], stage1_25[157], stage1_25[158], stage1_25[159], stage1_25[160], stage1_25[161]},
      {stage2_27[26],stage2_26[49],stage2_25[49],stage2_24[72],stage2_23[105]}
   );
   gpc615_5 gpc2705 (
      {stage1_23[158], stage1_23[159], stage1_23[160], stage1_23[161], stage1_23[162]},
      {stage1_24[165]},
      {stage1_25[162], stage1_25[163], stage1_25[164], stage1_25[165], stage1_25[166], stage1_25[167]},
      {stage2_27[27],stage2_26[50],stage2_25[50],stage2_24[73],stage2_23[106]}
   );
   gpc615_5 gpc2706 (
      {stage1_23[163], stage1_23[164], stage1_23[165], stage1_23[166], stage1_23[167]},
      {stage1_24[166]},
      {stage1_25[168], stage1_25[169], stage1_25[170], stage1_25[171], stage1_25[172], stage1_25[173]},
      {stage2_27[28],stage2_26[51],stage2_25[51],stage2_24[74],stage2_23[107]}
   );
   gpc615_5 gpc2707 (
      {stage1_23[168], stage1_23[169], stage1_23[170], stage1_23[171], stage1_23[172]},
      {stage1_24[167]},
      {stage1_25[174], stage1_25[175], stage1_25[176], stage1_25[177], stage1_25[178], stage1_25[179]},
      {stage2_27[29],stage2_26[52],stage2_25[52],stage2_24[75],stage2_23[108]}
   );
   gpc615_5 gpc2708 (
      {stage1_23[173], stage1_23[174], stage1_23[175], stage1_23[176], stage1_23[177]},
      {stage1_24[168]},
      {stage1_25[180], stage1_25[181], stage1_25[182], stage1_25[183], stage1_25[184], stage1_25[185]},
      {stage2_27[30],stage2_26[53],stage2_25[53],stage2_24[76],stage2_23[109]}
   );
   gpc615_5 gpc2709 (
      {stage1_24[169], stage1_24[170], stage1_24[171], stage1_24[172], stage1_24[173]},
      {stage1_25[186]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[31],stage2_26[54],stage2_25[54],stage2_24[77]}
   );
   gpc615_5 gpc2710 (
      {stage1_24[174], stage1_24[175], stage1_24[176], stage1_24[177], stage1_24[178]},
      {stage1_25[187]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[32],stage2_26[55],stage2_25[55],stage2_24[78]}
   );
   gpc615_5 gpc2711 (
      {stage1_24[179], stage1_24[180], stage1_24[181], stage1_24[182], stage1_24[183]},
      {stage1_25[188]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[33],stage2_26[56],stage2_25[56],stage2_24[79]}
   );
   gpc615_5 gpc2712 (
      {stage1_24[184], stage1_24[185], stage1_24[186], stage1_24[187], stage1_24[188]},
      {stage1_25[189]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[34],stage2_26[57],stage2_25[57],stage2_24[80]}
   );
   gpc615_5 gpc2713 (
      {stage1_24[189], stage1_24[190], stage1_24[191], stage1_24[192], stage1_24[193]},
      {stage1_25[190]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[35],stage2_26[58],stage2_25[58],stage2_24[81]}
   );
   gpc606_5 gpc2714 (
      {stage1_25[191], stage1_25[192], stage1_25[193], stage1_25[194], stage1_25[195], stage1_25[196]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[5],stage2_27[36],stage2_26[59],stage2_25[59]}
   );
   gpc606_5 gpc2715 (
      {stage1_25[197], stage1_25[198], stage1_25[199], stage1_25[200], stage1_25[201], stage1_25[202]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[6],stage2_27[37],stage2_26[60],stage2_25[60]}
   );
   gpc606_5 gpc2716 (
      {stage1_25[203], stage1_25[204], stage1_25[205], stage1_25[206], stage1_25[207], stage1_25[208]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[7],stage2_27[38],stage2_26[61],stage2_25[61]}
   );
   gpc615_5 gpc2717 (
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34]},
      {stage1_27[18]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[3],stage2_28[8],stage2_27[39],stage2_26[62]}
   );
   gpc615_5 gpc2718 (
      {stage1_26[35], stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39]},
      {stage1_27[19]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[4],stage2_28[9],stage2_27[40],stage2_26[63]}
   );
   gpc615_5 gpc2719 (
      {stage1_26[40], stage1_26[41], stage1_26[42], stage1_26[43], stage1_26[44]},
      {stage1_27[20]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[5],stage2_28[10],stage2_27[41],stage2_26[64]}
   );
   gpc615_5 gpc2720 (
      {stage1_26[45], stage1_26[46], stage1_26[47], stage1_26[48], stage1_26[49]},
      {stage1_27[21]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[6],stage2_28[11],stage2_27[42],stage2_26[65]}
   );
   gpc615_5 gpc2721 (
      {stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53], stage1_26[54]},
      {stage1_27[22]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[7],stage2_28[12],stage2_27[43],stage2_26[66]}
   );
   gpc615_5 gpc2722 (
      {stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58], stage1_26[59]},
      {stage1_27[23]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[8],stage2_28[13],stage2_27[44],stage2_26[67]}
   );
   gpc615_5 gpc2723 (
      {stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63], stage1_26[64]},
      {stage1_27[24]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[9],stage2_28[14],stage2_27[45],stage2_26[68]}
   );
   gpc615_5 gpc2724 (
      {stage1_26[65], stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69]},
      {stage1_27[25]},
      {stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45], stage1_28[46], stage1_28[47]},
      {stage2_30[7],stage2_29[10],stage2_28[15],stage2_27[46],stage2_26[69]}
   );
   gpc615_5 gpc2725 (
      {stage1_26[70], stage1_26[71], stage1_26[72], stage1_26[73], stage1_26[74]},
      {stage1_27[26]},
      {stage1_28[48], stage1_28[49], stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53]},
      {stage2_30[8],stage2_29[11],stage2_28[16],stage2_27[47],stage2_26[70]}
   );
   gpc615_5 gpc2726 (
      {stage1_26[75], stage1_26[76], stage1_26[77], stage1_26[78], stage1_26[79]},
      {stage1_27[27]},
      {stage1_28[54], stage1_28[55], stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59]},
      {stage2_30[9],stage2_29[12],stage2_28[17],stage2_27[48],stage2_26[71]}
   );
   gpc615_5 gpc2727 (
      {stage1_26[80], stage1_26[81], stage1_26[82], stage1_26[83], stage1_26[84]},
      {stage1_27[28]},
      {stage1_28[60], stage1_28[61], stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65]},
      {stage2_30[10],stage2_29[13],stage2_28[18],stage2_27[49],stage2_26[72]}
   );
   gpc615_5 gpc2728 (
      {stage1_26[85], stage1_26[86], stage1_26[87], stage1_26[88], stage1_26[89]},
      {stage1_27[29]},
      {stage1_28[66], stage1_28[67], stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71]},
      {stage2_30[11],stage2_29[14],stage2_28[19],stage2_27[50],stage2_26[73]}
   );
   gpc615_5 gpc2729 (
      {stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93], stage1_26[94]},
      {stage1_27[30]},
      {stage1_28[72], stage1_28[73], stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77]},
      {stage2_30[12],stage2_29[15],stage2_28[20],stage2_27[51],stage2_26[74]}
   );
   gpc615_5 gpc2730 (
      {stage1_26[95], stage1_26[96], stage1_26[97], stage1_26[98], stage1_26[99]},
      {stage1_27[31]},
      {stage1_28[78], stage1_28[79], stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83]},
      {stage2_30[13],stage2_29[16],stage2_28[21],stage2_27[52],stage2_26[75]}
   );
   gpc615_5 gpc2731 (
      {stage1_26[100], stage1_26[101], stage1_26[102], stage1_26[103], stage1_26[104]},
      {stage1_27[32]},
      {stage1_28[84], stage1_28[85], stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89]},
      {stage2_30[14],stage2_29[17],stage2_28[22],stage2_27[53],stage2_26[76]}
   );
   gpc615_5 gpc2732 (
      {stage1_26[105], stage1_26[106], stage1_26[107], stage1_26[108], stage1_26[109]},
      {stage1_27[33]},
      {stage1_28[90], stage1_28[91], stage1_28[92], stage1_28[93], stage1_28[94], stage1_28[95]},
      {stage2_30[15],stage2_29[18],stage2_28[23],stage2_27[54],stage2_26[77]}
   );
   gpc615_5 gpc2733 (
      {stage1_26[110], stage1_26[111], stage1_26[112], stage1_26[113], stage1_26[114]},
      {stage1_27[34]},
      {stage1_28[96], stage1_28[97], stage1_28[98], stage1_28[99], stage1_28[100], stage1_28[101]},
      {stage2_30[16],stage2_29[19],stage2_28[24],stage2_27[55],stage2_26[78]}
   );
   gpc615_5 gpc2734 (
      {stage1_26[115], stage1_26[116], stage1_26[117], stage1_26[118], stage1_26[119]},
      {stage1_27[35]},
      {stage1_28[102], stage1_28[103], stage1_28[104], stage1_28[105], stage1_28[106], stage1_28[107]},
      {stage2_30[17],stage2_29[20],stage2_28[25],stage2_27[56],stage2_26[79]}
   );
   gpc615_5 gpc2735 (
      {stage1_26[120], stage1_26[121], stage1_26[122], stage1_26[123], stage1_26[124]},
      {stage1_27[36]},
      {stage1_28[108], stage1_28[109], stage1_28[110], stage1_28[111], stage1_28[112], stage1_28[113]},
      {stage2_30[18],stage2_29[21],stage2_28[26],stage2_27[57],stage2_26[80]}
   );
   gpc615_5 gpc2736 (
      {stage1_26[125], stage1_26[126], stage1_26[127], stage1_26[128], stage1_26[129]},
      {stage1_27[37]},
      {stage1_28[114], stage1_28[115], stage1_28[116], stage1_28[117], stage1_28[118], stage1_28[119]},
      {stage2_30[19],stage2_29[22],stage2_28[27],stage2_27[58],stage2_26[81]}
   );
   gpc615_5 gpc2737 (
      {stage1_26[130], stage1_26[131], stage1_26[132], stage1_26[133], stage1_26[134]},
      {stage1_27[38]},
      {stage1_28[120], stage1_28[121], stage1_28[122], stage1_28[123], stage1_28[124], stage1_28[125]},
      {stage2_30[20],stage2_29[23],stage2_28[28],stage2_27[59],stage2_26[82]}
   );
   gpc615_5 gpc2738 (
      {stage1_26[135], stage1_26[136], stage1_26[137], stage1_26[138], stage1_26[139]},
      {stage1_27[39]},
      {stage1_28[126], stage1_28[127], stage1_28[128], stage1_28[129], stage1_28[130], stage1_28[131]},
      {stage2_30[21],stage2_29[24],stage2_28[29],stage2_27[60],stage2_26[83]}
   );
   gpc615_5 gpc2739 (
      {stage1_26[140], stage1_26[141], stage1_26[142], stage1_26[143], stage1_26[144]},
      {stage1_27[40]},
      {stage1_28[132], stage1_28[133], stage1_28[134], stage1_28[135], stage1_28[136], stage1_28[137]},
      {stage2_30[22],stage2_29[25],stage2_28[30],stage2_27[61],stage2_26[84]}
   );
   gpc615_5 gpc2740 (
      {stage1_26[145], stage1_26[146], stage1_26[147], stage1_26[148], stage1_26[149]},
      {stage1_27[41]},
      {stage1_28[138], stage1_28[139], stage1_28[140], stage1_28[141], stage1_28[142], stage1_28[143]},
      {stage2_30[23],stage2_29[26],stage2_28[31],stage2_27[62],stage2_26[85]}
   );
   gpc615_5 gpc2741 (
      {stage1_26[150], stage1_26[151], stage1_26[152], stage1_26[153], stage1_26[154]},
      {stage1_27[42]},
      {stage1_28[144], stage1_28[145], stage1_28[146], stage1_28[147], stage1_28[148], stage1_28[149]},
      {stage2_30[24],stage2_29[27],stage2_28[32],stage2_27[63],stage2_26[86]}
   );
   gpc615_5 gpc2742 (
      {stage1_26[155], stage1_26[156], stage1_26[157], stage1_26[158], stage1_26[159]},
      {stage1_27[43]},
      {stage1_28[150], stage1_28[151], stage1_28[152], stage1_28[153], stage1_28[154], stage1_28[155]},
      {stage2_30[25],stage2_29[28],stage2_28[33],stage2_27[64],stage2_26[87]}
   );
   gpc615_5 gpc2743 (
      {stage1_26[160], stage1_26[161], stage1_26[162], stage1_26[163], stage1_26[164]},
      {stage1_27[44]},
      {stage1_28[156], stage1_28[157], stage1_28[158], stage1_28[159], stage1_28[160], stage1_28[161]},
      {stage2_30[26],stage2_29[29],stage2_28[34],stage2_27[65],stage2_26[88]}
   );
   gpc615_5 gpc2744 (
      {stage1_26[165], stage1_26[166], stage1_26[167], stage1_26[168], stage1_26[169]},
      {stage1_27[45]},
      {stage1_28[162], stage1_28[163], stage1_28[164], stage1_28[165], stage1_28[166], stage1_28[167]},
      {stage2_30[27],stage2_29[30],stage2_28[35],stage2_27[66],stage2_26[89]}
   );
   gpc615_5 gpc2745 (
      {stage1_26[170], stage1_26[171], stage1_26[172], stage1_26[173], stage1_26[174]},
      {stage1_27[46]},
      {stage1_28[168], stage1_28[169], stage1_28[170], stage1_28[171], stage1_28[172], stage1_28[173]},
      {stage2_30[28],stage2_29[31],stage2_28[36],stage2_27[67],stage2_26[90]}
   );
   gpc615_5 gpc2746 (
      {stage1_26[175], stage1_26[176], stage1_26[177], stage1_26[178], stage1_26[179]},
      {stage1_27[47]},
      {stage1_28[174], stage1_28[175], stage1_28[176], stage1_28[177], stage1_28[178], stage1_28[179]},
      {stage2_30[29],stage2_29[32],stage2_28[37],stage2_27[68],stage2_26[91]}
   );
   gpc615_5 gpc2747 (
      {stage1_26[180], stage1_26[181], stage1_26[182], stage1_26[183], stage1_26[184]},
      {stage1_27[48]},
      {stage1_28[180], stage1_28[181], stage1_28[182], stage1_28[183], stage1_28[184], stage1_28[185]},
      {stage2_30[30],stage2_29[33],stage2_28[38],stage2_27[69],stage2_26[92]}
   );
   gpc615_5 gpc2748 (
      {stage1_26[185], stage1_26[186], stage1_26[187], stage1_26[188], stage1_26[189]},
      {stage1_27[49]},
      {stage1_28[186], stage1_28[187], stage1_28[188], stage1_28[189], stage1_28[190], stage1_28[191]},
      {stage2_30[31],stage2_29[34],stage2_28[39],stage2_27[70],stage2_26[93]}
   );
   gpc615_5 gpc2749 (
      {stage1_26[190], stage1_26[191], stage1_26[192], stage1_26[193], stage1_26[194]},
      {stage1_27[50]},
      {stage1_28[192], stage1_28[193], stage1_28[194], stage1_28[195], stage1_28[196], stage1_28[197]},
      {stage2_30[32],stage2_29[35],stage2_28[40],stage2_27[71],stage2_26[94]}
   );
   gpc615_5 gpc2750 (
      {stage1_26[195], stage1_26[196], stage1_26[197], stage1_26[198], stage1_26[199]},
      {stage1_27[51]},
      {stage1_28[198], stage1_28[199], stage1_28[200], stage1_28[201], stage1_28[202], stage1_28[203]},
      {stage2_30[33],stage2_29[36],stage2_28[41],stage2_27[72],stage2_26[95]}
   );
   gpc615_5 gpc2751 (
      {stage1_26[200], stage1_26[201], stage1_26[202], stage1_26[203], stage1_26[204]},
      {stage1_27[52]},
      {stage1_28[204], stage1_28[205], stage1_28[206], stage1_28[207], stage1_28[208], stage1_28[209]},
      {stage2_30[34],stage2_29[37],stage2_28[42],stage2_27[73],stage2_26[96]}
   );
   gpc615_5 gpc2752 (
      {stage1_26[205], stage1_26[206], stage1_26[207], stage1_26[208], stage1_26[209]},
      {stage1_27[53]},
      {stage1_28[210], stage1_28[211], stage1_28[212], stage1_28[213], stage1_28[214], stage1_28[215]},
      {stage2_30[35],stage2_29[38],stage2_28[43],stage2_27[74],stage2_26[97]}
   );
   gpc615_5 gpc2753 (
      {stage1_26[210], stage1_26[211], stage1_26[212], stage1_26[213], stage1_26[214]},
      {stage1_27[54]},
      {stage1_28[216], stage1_28[217], stage1_28[218], stage1_28[219], stage1_28[220], stage1_28[221]},
      {stage2_30[36],stage2_29[39],stage2_28[44],stage2_27[75],stage2_26[98]}
   );
   gpc615_5 gpc2754 (
      {stage1_27[55], stage1_27[56], stage1_27[57], stage1_27[58], stage1_27[59]},
      {stage1_28[222]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[37],stage2_29[40],stage2_28[45],stage2_27[76]}
   );
   gpc615_5 gpc2755 (
      {stage1_27[60], stage1_27[61], stage1_27[62], stage1_27[63], stage1_27[64]},
      {stage1_28[223]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[38],stage2_29[41],stage2_28[46],stage2_27[77]}
   );
   gpc615_5 gpc2756 (
      {stage1_27[65], stage1_27[66], stage1_27[67], stage1_27[68], stage1_27[69]},
      {stage1_28[224]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[39],stage2_29[42],stage2_28[47],stage2_27[78]}
   );
   gpc615_5 gpc2757 (
      {stage1_27[70], stage1_27[71], stage1_27[72], stage1_27[73], stage1_27[74]},
      {stage1_28[225]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[40],stage2_29[43],stage2_28[48],stage2_27[79]}
   );
   gpc615_5 gpc2758 (
      {stage1_27[75], stage1_27[76], stage1_27[77], stage1_27[78], stage1_27[79]},
      {stage1_28[226]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[41],stage2_29[44],stage2_28[49],stage2_27[80]}
   );
   gpc615_5 gpc2759 (
      {stage1_27[80], stage1_27[81], stage1_27[82], stage1_27[83], stage1_27[84]},
      {stage1_28[227]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[42],stage2_29[45],stage2_28[50],stage2_27[81]}
   );
   gpc615_5 gpc2760 (
      {stage1_27[85], stage1_27[86], stage1_27[87], stage1_27[88], stage1_27[89]},
      {stage1_28[228]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[43],stage2_29[46],stage2_28[51],stage2_27[82]}
   );
   gpc615_5 gpc2761 (
      {stage1_27[90], stage1_27[91], stage1_27[92], stage1_27[93], stage1_27[94]},
      {stage1_28[229]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[44],stage2_29[47],stage2_28[52],stage2_27[83]}
   );
   gpc615_5 gpc2762 (
      {stage1_27[95], stage1_27[96], stage1_27[97], stage1_27[98], stage1_27[99]},
      {stage1_28[230]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[45],stage2_29[48],stage2_28[53],stage2_27[84]}
   );
   gpc615_5 gpc2763 (
      {stage1_27[100], stage1_27[101], stage1_27[102], stage1_27[103], stage1_27[104]},
      {stage1_28[231]},
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage2_31[9],stage2_30[46],stage2_29[49],stage2_28[54],stage2_27[85]}
   );
   gpc615_5 gpc2764 (
      {stage1_27[105], stage1_27[106], stage1_27[107], stage1_27[108], stage1_27[109]},
      {stage1_28[232]},
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage2_31[10],stage2_30[47],stage2_29[50],stage2_28[55],stage2_27[86]}
   );
   gpc615_5 gpc2765 (
      {stage1_27[110], stage1_27[111], stage1_27[112], stage1_27[113], stage1_27[114]},
      {stage1_28[233]},
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage2_31[11],stage2_30[48],stage2_29[51],stage2_28[56],stage2_27[87]}
   );
   gpc615_5 gpc2766 (
      {stage1_27[115], stage1_27[116], stage1_27[117], stage1_27[118], stage1_27[119]},
      {stage1_28[234]},
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage2_31[12],stage2_30[49],stage2_29[52],stage2_28[57],stage2_27[88]}
   );
   gpc615_5 gpc2767 (
      {stage1_27[120], stage1_27[121], stage1_27[122], stage1_27[123], stage1_27[124]},
      {stage1_28[235]},
      {stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82], stage1_29[83]},
      {stage2_31[13],stage2_30[50],stage2_29[53],stage2_28[58],stage2_27[89]}
   );
   gpc615_5 gpc2768 (
      {stage1_27[125], stage1_27[126], stage1_27[127], stage1_27[128], stage1_27[129]},
      {stage1_28[236]},
      {stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88], stage1_29[89]},
      {stage2_31[14],stage2_30[51],stage2_29[54],stage2_28[59],stage2_27[90]}
   );
   gpc615_5 gpc2769 (
      {stage1_27[130], stage1_27[131], stage1_27[132], stage1_27[133], stage1_27[134]},
      {stage1_28[237]},
      {stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93], stage1_29[94], stage1_29[95]},
      {stage2_31[15],stage2_30[52],stage2_29[55],stage2_28[60],stage2_27[91]}
   );
   gpc615_5 gpc2770 (
      {stage1_27[135], stage1_27[136], stage1_27[137], stage1_27[138], stage1_27[139]},
      {stage1_28[238]},
      {stage1_29[96], stage1_29[97], stage1_29[98], stage1_29[99], stage1_29[100], stage1_29[101]},
      {stage2_31[16],stage2_30[53],stage2_29[56],stage2_28[61],stage2_27[92]}
   );
   gpc615_5 gpc2771 (
      {stage1_27[140], stage1_27[141], stage1_27[142], stage1_27[143], stage1_27[144]},
      {stage1_28[239]},
      {stage1_29[102], stage1_29[103], stage1_29[104], stage1_29[105], stage1_29[106], stage1_29[107]},
      {stage2_31[17],stage2_30[54],stage2_29[57],stage2_28[62],stage2_27[93]}
   );
   gpc615_5 gpc2772 (
      {stage1_27[145], stage1_27[146], stage1_27[147], stage1_27[148], stage1_27[149]},
      {stage1_28[240]},
      {stage1_29[108], stage1_29[109], stage1_29[110], stage1_29[111], stage1_29[112], stage1_29[113]},
      {stage2_31[18],stage2_30[55],stage2_29[58],stage2_28[63],stage2_27[94]}
   );
   gpc615_5 gpc2773 (
      {stage1_27[150], stage1_27[151], stage1_27[152], stage1_27[153], stage1_27[154]},
      {stage1_28[241]},
      {stage1_29[114], stage1_29[115], stage1_29[116], stage1_29[117], stage1_29[118], stage1_29[119]},
      {stage2_31[19],stage2_30[56],stage2_29[59],stage2_28[64],stage2_27[95]}
   );
   gpc615_5 gpc2774 (
      {stage1_27[155], stage1_27[156], stage1_27[157], stage1_27[158], 1'b0},
      {stage1_28[242]},
      {stage1_29[120], stage1_29[121], stage1_29[122], stage1_29[123], stage1_29[124], stage1_29[125]},
      {stage2_31[20],stage2_30[57],stage2_29[60],stage2_28[65],stage2_27[96]}
   );
   gpc606_5 gpc2775 (
      {stage1_29[126], stage1_29[127], stage1_29[128], stage1_29[129], stage1_29[130], stage1_29[131]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[0],stage2_31[21],stage2_30[58],stage2_29[61]}
   );
   gpc606_5 gpc2776 (
      {stage1_29[132], stage1_29[133], stage1_29[134], stage1_29[135], stage1_29[136], stage1_29[137]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[1],stage2_31[22],stage2_30[59],stage2_29[62]}
   );
   gpc606_5 gpc2777 (
      {stage1_29[138], stage1_29[139], stage1_29[140], stage1_29[141], stage1_29[142], stage1_29[143]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[2],stage2_31[23],stage2_30[60],stage2_29[63]}
   );
   gpc606_5 gpc2778 (
      {stage1_29[144], stage1_29[145], stage1_29[146], stage1_29[147], stage1_29[148], stage1_29[149]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[3],stage2_31[24],stage2_30[61],stage2_29[64]}
   );
   gpc606_5 gpc2779 (
      {stage1_29[150], stage1_29[151], stage1_29[152], stage1_29[153], stage1_29[154], stage1_29[155]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[4],stage2_31[25],stage2_30[62],stage2_29[65]}
   );
   gpc606_5 gpc2780 (
      {stage1_29[156], stage1_29[157], stage1_29[158], stage1_29[159], stage1_29[160], stage1_29[161]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[5],stage2_31[26],stage2_30[63],stage2_29[66]}
   );
   gpc606_5 gpc2781 (
      {stage1_29[162], stage1_29[163], stage1_29[164], stage1_29[165], stage1_29[166], stage1_29[167]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[6],stage2_31[27],stage2_30[64],stage2_29[67]}
   );
   gpc606_5 gpc2782 (
      {stage1_29[168], stage1_29[169], stage1_29[170], stage1_29[171], stage1_29[172], stage1_29[173]},
      {stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47]},
      {stage2_33[7],stage2_32[7],stage2_31[28],stage2_30[65],stage2_29[68]}
   );
   gpc606_5 gpc2783 (
      {stage1_29[174], stage1_29[175], stage1_29[176], stage1_29[177], stage1_29[178], stage1_29[179]},
      {stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage2_33[8],stage2_32[8],stage2_31[29],stage2_30[66],stage2_29[69]}
   );
   gpc606_5 gpc2784 (
      {stage1_29[180], stage1_29[181], stage1_29[182], stage1_29[183], stage1_29[184], stage1_29[185]},
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59]},
      {stage2_33[9],stage2_32[9],stage2_31[30],stage2_30[67],stage2_29[70]}
   );
   gpc606_5 gpc2785 (
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[10],stage2_32[10],stage2_31[31],stage2_30[68]}
   );
   gpc606_5 gpc2786 (
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[11],stage2_32[11],stage2_31[32],stage2_30[69]}
   );
   gpc606_5 gpc2787 (
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[12],stage2_32[12],stage2_31[33],stage2_30[70]}
   );
   gpc606_5 gpc2788 (
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[13],stage2_32[13],stage2_31[34],stage2_30[71]}
   );
   gpc606_5 gpc2789 (
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27], stage1_32[28], stage1_32[29]},
      {stage2_34[4],stage2_33[14],stage2_32[14],stage2_31[35],stage2_30[72]}
   );
   gpc606_5 gpc2790 (
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33], stage1_32[34], stage1_32[35]},
      {stage2_34[5],stage2_33[15],stage2_32[15],stage2_31[36],stage2_30[73]}
   );
   gpc606_5 gpc2791 (
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39], stage1_32[40], stage1_32[41]},
      {stage2_34[6],stage2_33[16],stage2_32[16],stage2_31[37],stage2_30[74]}
   );
   gpc606_5 gpc2792 (
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45], stage1_32[46], stage1_32[47]},
      {stage2_34[7],stage2_33[17],stage2_32[17],stage2_31[38],stage2_30[75]}
   );
   gpc606_5 gpc2793 (
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51], stage1_32[52], stage1_32[53]},
      {stage2_34[8],stage2_33[18],stage2_32[18],stage2_31[39],stage2_30[76]}
   );
   gpc606_5 gpc2794 (
      {stage1_30[54], stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59]},
      {stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57], stage1_32[58], stage1_32[59]},
      {stage2_34[9],stage2_33[19],stage2_32[19],stage2_31[40],stage2_30[77]}
   );
   gpc606_5 gpc2795 (
      {stage1_30[60], stage1_30[61], stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65]},
      {stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63], stage1_32[64], stage1_32[65]},
      {stage2_34[10],stage2_33[20],stage2_32[20],stage2_31[41],stage2_30[78]}
   );
   gpc606_5 gpc2796 (
      {stage1_30[66], stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69], stage1_32[70], stage1_32[71]},
      {stage2_34[11],stage2_33[21],stage2_32[21],stage2_31[42],stage2_30[79]}
   );
   gpc606_5 gpc2797 (
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76], stage1_30[77]},
      {stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75], stage1_32[76], stage1_32[77]},
      {stage2_34[12],stage2_33[22],stage2_32[22],stage2_31[43],stage2_30[80]}
   );
   gpc606_5 gpc2798 (
      {stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81], stage1_30[82], stage1_30[83]},
      {stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81], stage1_32[82], stage1_32[83]},
      {stage2_34[13],stage2_33[23],stage2_32[23],stage2_31[44],stage2_30[81]}
   );
   gpc606_5 gpc2799 (
      {stage1_30[84], stage1_30[85], stage1_30[86], stage1_30[87], stage1_30[88], stage1_30[89]},
      {stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87], stage1_32[88], stage1_32[89]},
      {stage2_34[14],stage2_33[24],stage2_32[24],stage2_31[45],stage2_30[82]}
   );
   gpc606_5 gpc2800 (
      {stage1_30[90], stage1_30[91], stage1_30[92], stage1_30[93], stage1_30[94], stage1_30[95]},
      {stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93], stage1_32[94], stage1_32[95]},
      {stage2_34[15],stage2_33[25],stage2_32[25],stage2_31[46],stage2_30[83]}
   );
   gpc606_5 gpc2801 (
      {stage1_30[96], stage1_30[97], stage1_30[98], stage1_30[99], stage1_30[100], stage1_30[101]},
      {stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99], stage1_32[100], stage1_32[101]},
      {stage2_34[16],stage2_33[26],stage2_32[26],stage2_31[47],stage2_30[84]}
   );
   gpc606_5 gpc2802 (
      {stage1_30[102], stage1_30[103], stage1_30[104], stage1_30[105], stage1_30[106], stage1_30[107]},
      {stage1_32[102], stage1_32[103], stage1_32[104], stage1_32[105], stage1_32[106], stage1_32[107]},
      {stage2_34[17],stage2_33[27],stage2_32[27],stage2_31[48],stage2_30[85]}
   );
   gpc606_5 gpc2803 (
      {stage1_30[108], stage1_30[109], stage1_30[110], stage1_30[111], stage1_30[112], stage1_30[113]},
      {stage1_32[108], stage1_32[109], stage1_32[110], stage1_32[111], stage1_32[112], stage1_32[113]},
      {stage2_34[18],stage2_33[28],stage2_32[28],stage2_31[49],stage2_30[86]}
   );
   gpc606_5 gpc2804 (
      {stage1_30[114], stage1_30[115], stage1_30[116], stage1_30[117], stage1_30[118], stage1_30[119]},
      {stage1_32[114], stage1_32[115], stage1_32[116], stage1_32[117], stage1_32[118], stage1_32[119]},
      {stage2_34[19],stage2_33[29],stage2_32[29],stage2_31[50],stage2_30[87]}
   );
   gpc606_5 gpc2805 (
      {stage1_30[120], stage1_30[121], stage1_30[122], stage1_30[123], stage1_30[124], stage1_30[125]},
      {stage1_32[120], stage1_32[121], stage1_32[122], stage1_32[123], stage1_32[124], stage1_32[125]},
      {stage2_34[20],stage2_33[30],stage2_32[30],stage2_31[51],stage2_30[88]}
   );
   gpc606_5 gpc2806 (
      {stage1_30[126], stage1_30[127], stage1_30[128], stage1_30[129], stage1_30[130], stage1_30[131]},
      {stage1_32[126], stage1_32[127], stage1_32[128], stage1_32[129], stage1_32[130], stage1_32[131]},
      {stage2_34[21],stage2_33[31],stage2_32[31],stage2_31[52],stage2_30[89]}
   );
   gpc606_5 gpc2807 (
      {stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63], stage1_31[64], stage1_31[65]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[22],stage2_33[32],stage2_32[32],stage2_31[53]}
   );
   gpc606_5 gpc2808 (
      {stage1_31[66], stage1_31[67], stage1_31[68], stage1_31[69], stage1_31[70], stage1_31[71]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[23],stage2_33[33],stage2_32[33],stage2_31[54]}
   );
   gpc606_5 gpc2809 (
      {stage1_31[72], stage1_31[73], stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[24],stage2_33[34],stage2_32[34],stage2_31[55]}
   );
   gpc606_5 gpc2810 (
      {stage1_31[78], stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[25],stage2_33[35],stage2_32[35],stage2_31[56]}
   );
   gpc606_5 gpc2811 (
      {stage1_31[84], stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88], stage1_31[89]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[26],stage2_33[36],stage2_32[36],stage2_31[57]}
   );
   gpc606_5 gpc2812 (
      {stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93], stage1_31[94], stage1_31[95]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage2_35[5],stage2_34[27],stage2_33[37],stage2_32[37],stage2_31[58]}
   );
   gpc606_5 gpc2813 (
      {stage1_31[96], stage1_31[97], stage1_31[98], stage1_31[99], stage1_31[100], stage1_31[101]},
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41]},
      {stage2_35[6],stage2_34[28],stage2_33[38],stage2_32[38],stage2_31[59]}
   );
   gpc606_5 gpc2814 (
      {stage1_31[102], stage1_31[103], stage1_31[104], stage1_31[105], stage1_31[106], stage1_31[107]},
      {stage1_33[42], stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47]},
      {stage2_35[7],stage2_34[29],stage2_33[39],stage2_32[39],stage2_31[60]}
   );
   gpc606_5 gpc2815 (
      {stage1_31[108], stage1_31[109], stage1_31[110], stage1_31[111], stage1_31[112], stage1_31[113]},
      {stage1_33[48], stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53]},
      {stage2_35[8],stage2_34[30],stage2_33[40],stage2_32[40],stage2_31[61]}
   );
   gpc606_5 gpc2816 (
      {stage1_31[114], stage1_31[115], stage1_31[116], stage1_31[117], stage1_31[118], stage1_31[119]},
      {stage1_33[54], stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59]},
      {stage2_35[9],stage2_34[31],stage2_33[41],stage2_32[41],stage2_31[62]}
   );
   gpc606_5 gpc2817 (
      {stage1_31[120], stage1_31[121], stage1_31[122], stage1_31[123], stage1_31[124], stage1_31[125]},
      {stage1_33[60], stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65]},
      {stage2_35[10],stage2_34[32],stage2_33[42],stage2_32[42],stage2_31[63]}
   );
   gpc606_5 gpc2818 (
      {stage1_31[126], stage1_31[127], stage1_31[128], stage1_31[129], stage1_31[130], stage1_31[131]},
      {stage1_33[66], stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71]},
      {stage2_35[11],stage2_34[33],stage2_33[43],stage2_32[43],stage2_31[64]}
   );
   gpc606_5 gpc2819 (
      {stage1_31[132], stage1_31[133], stage1_31[134], stage1_31[135], stage1_31[136], stage1_31[137]},
      {stage1_33[72], stage1_33[73], stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77]},
      {stage2_35[12],stage2_34[34],stage2_33[44],stage2_32[44],stage2_31[65]}
   );
   gpc606_5 gpc2820 (
      {stage1_31[138], stage1_31[139], stage1_31[140], stage1_31[141], stage1_31[142], stage1_31[143]},
      {stage1_33[78], stage1_33[79], stage1_33[80], 1'b0, 1'b0, 1'b0},
      {stage2_35[13],stage2_34[35],stage2_33[45],stage2_32[45],stage2_31[66]}
   );
   gpc1_1 gpc2821 (
      {stage1_1[62]},
      {stage2_1[31]}
   );
   gpc1_1 gpc2822 (
      {stage1_1[63]},
      {stage2_1[32]}
   );
   gpc1_1 gpc2823 (
      {stage1_1[64]},
      {stage2_1[33]}
   );
   gpc1_1 gpc2824 (
      {stage1_1[65]},
      {stage2_1[34]}
   );
   gpc1_1 gpc2825 (
      {stage1_1[66]},
      {stage2_1[35]}
   );
   gpc1_1 gpc2826 (
      {stage1_1[67]},
      {stage2_1[36]}
   );
   gpc1_1 gpc2827 (
      {stage1_1[68]},
      {stage2_1[37]}
   );
   gpc1_1 gpc2828 (
      {stage1_1[69]},
      {stage2_1[38]}
   );
   gpc1_1 gpc2829 (
      {stage1_1[70]},
      {stage2_1[39]}
   );
   gpc1_1 gpc2830 (
      {stage1_1[71]},
      {stage2_1[40]}
   );
   gpc1_1 gpc2831 (
      {stage1_1[72]},
      {stage2_1[41]}
   );
   gpc1_1 gpc2832 (
      {stage1_1[73]},
      {stage2_1[42]}
   );
   gpc1_1 gpc2833 (
      {stage1_1[74]},
      {stage2_1[43]}
   );
   gpc1_1 gpc2834 (
      {stage1_1[75]},
      {stage2_1[44]}
   );
   gpc1_1 gpc2835 (
      {stage1_1[76]},
      {stage2_1[45]}
   );
   gpc1_1 gpc2836 (
      {stage1_1[77]},
      {stage2_1[46]}
   );
   gpc1_1 gpc2837 (
      {stage1_1[78]},
      {stage2_1[47]}
   );
   gpc1_1 gpc2838 (
      {stage1_1[79]},
      {stage2_1[48]}
   );
   gpc1_1 gpc2839 (
      {stage1_1[80]},
      {stage2_1[49]}
   );
   gpc1_1 gpc2840 (
      {stage1_1[81]},
      {stage2_1[50]}
   );
   gpc1_1 gpc2841 (
      {stage1_1[82]},
      {stage2_1[51]}
   );
   gpc1_1 gpc2842 (
      {stage1_1[83]},
      {stage2_1[52]}
   );
   gpc1_1 gpc2843 (
      {stage1_1[84]},
      {stage2_1[53]}
   );
   gpc1_1 gpc2844 (
      {stage1_1[85]},
      {stage2_1[54]}
   );
   gpc1_1 gpc2845 (
      {stage1_1[86]},
      {stage2_1[55]}
   );
   gpc1_1 gpc2846 (
      {stage1_1[87]},
      {stage2_1[56]}
   );
   gpc1_1 gpc2847 (
      {stage1_1[88]},
      {stage2_1[57]}
   );
   gpc1_1 gpc2848 (
      {stage1_1[89]},
      {stage2_1[58]}
   );
   gpc1_1 gpc2849 (
      {stage1_1[90]},
      {stage2_1[59]}
   );
   gpc1_1 gpc2850 (
      {stage1_1[91]},
      {stage2_1[60]}
   );
   gpc1_1 gpc2851 (
      {stage1_1[92]},
      {stage2_1[61]}
   );
   gpc1_1 gpc2852 (
      {stage1_1[93]},
      {stage2_1[62]}
   );
   gpc1_1 gpc2853 (
      {stage1_1[94]},
      {stage2_1[63]}
   );
   gpc1_1 gpc2854 (
      {stage1_1[95]},
      {stage2_1[64]}
   );
   gpc1_1 gpc2855 (
      {stage1_1[96]},
      {stage2_1[65]}
   );
   gpc1_1 gpc2856 (
      {stage1_1[97]},
      {stage2_1[66]}
   );
   gpc1_1 gpc2857 (
      {stage1_1[98]},
      {stage2_1[67]}
   );
   gpc1_1 gpc2858 (
      {stage1_1[99]},
      {stage2_1[68]}
   );
   gpc1_1 gpc2859 (
      {stage1_1[100]},
      {stage2_1[69]}
   );
   gpc1_1 gpc2860 (
      {stage1_1[101]},
      {stage2_1[70]}
   );
   gpc1_1 gpc2861 (
      {stage1_1[102]},
      {stage2_1[71]}
   );
   gpc1_1 gpc2862 (
      {stage1_1[103]},
      {stage2_1[72]}
   );
   gpc1_1 gpc2863 (
      {stage1_1[104]},
      {stage2_1[73]}
   );
   gpc1_1 gpc2864 (
      {stage1_1[105]},
      {stage2_1[74]}
   );
   gpc1_1 gpc2865 (
      {stage1_1[106]},
      {stage2_1[75]}
   );
   gpc1_1 gpc2866 (
      {stage1_1[107]},
      {stage2_1[76]}
   );
   gpc1_1 gpc2867 (
      {stage1_1[108]},
      {stage2_1[77]}
   );
   gpc1_1 gpc2868 (
      {stage1_1[109]},
      {stage2_1[78]}
   );
   gpc1_1 gpc2869 (
      {stage1_1[110]},
      {stage2_1[79]}
   );
   gpc1_1 gpc2870 (
      {stage1_1[111]},
      {stage2_1[80]}
   );
   gpc1_1 gpc2871 (
      {stage1_1[112]},
      {stage2_1[81]}
   );
   gpc1_1 gpc2872 (
      {stage1_1[113]},
      {stage2_1[82]}
   );
   gpc1_1 gpc2873 (
      {stage1_1[114]},
      {stage2_1[83]}
   );
   gpc1_1 gpc2874 (
      {stage1_1[115]},
      {stage2_1[84]}
   );
   gpc1_1 gpc2875 (
      {stage1_1[116]},
      {stage2_1[85]}
   );
   gpc1_1 gpc2876 (
      {stage1_1[117]},
      {stage2_1[86]}
   );
   gpc1_1 gpc2877 (
      {stage1_1[118]},
      {stage2_1[87]}
   );
   gpc1_1 gpc2878 (
      {stage1_1[119]},
      {stage2_1[88]}
   );
   gpc1_1 gpc2879 (
      {stage1_1[120]},
      {stage2_1[89]}
   );
   gpc1_1 gpc2880 (
      {stage1_1[121]},
      {stage2_1[90]}
   );
   gpc1_1 gpc2881 (
      {stage1_1[122]},
      {stage2_1[91]}
   );
   gpc1_1 gpc2882 (
      {stage1_1[123]},
      {stage2_1[92]}
   );
   gpc1_1 gpc2883 (
      {stage1_1[124]},
      {stage2_1[93]}
   );
   gpc1_1 gpc2884 (
      {stage1_1[125]},
      {stage2_1[94]}
   );
   gpc1_1 gpc2885 (
      {stage1_1[126]},
      {stage2_1[95]}
   );
   gpc1_1 gpc2886 (
      {stage1_1[127]},
      {stage2_1[96]}
   );
   gpc1_1 gpc2887 (
      {stage1_1[128]},
      {stage2_1[97]}
   );
   gpc1_1 gpc2888 (
      {stage1_1[129]},
      {stage2_1[98]}
   );
   gpc1_1 gpc2889 (
      {stage1_1[130]},
      {stage2_1[99]}
   );
   gpc1_1 gpc2890 (
      {stage1_1[131]},
      {stage2_1[100]}
   );
   gpc1_1 gpc2891 (
      {stage1_1[132]},
      {stage2_1[101]}
   );
   gpc1_1 gpc2892 (
      {stage1_1[133]},
      {stage2_1[102]}
   );
   gpc1_1 gpc2893 (
      {stage1_1[134]},
      {stage2_1[103]}
   );
   gpc1_1 gpc2894 (
      {stage1_1[135]},
      {stage2_1[104]}
   );
   gpc1_1 gpc2895 (
      {stage1_1[136]},
      {stage2_1[105]}
   );
   gpc1_1 gpc2896 (
      {stage1_1[137]},
      {stage2_1[106]}
   );
   gpc1_1 gpc2897 (
      {stage1_2[225]},
      {stage2_2[48]}
   );
   gpc1_1 gpc2898 (
      {stage1_2[226]},
      {stage2_2[49]}
   );
   gpc1_1 gpc2899 (
      {stage1_2[227]},
      {stage2_2[50]}
   );
   gpc1_1 gpc2900 (
      {stage1_3[169]},
      {stage2_3[69]}
   );
   gpc1_1 gpc2901 (
      {stage1_3[170]},
      {stage2_3[70]}
   );
   gpc1_1 gpc2902 (
      {stage1_3[171]},
      {stage2_3[71]}
   );
   gpc1_1 gpc2903 (
      {stage1_3[172]},
      {stage2_3[72]}
   );
   gpc1_1 gpc2904 (
      {stage1_3[173]},
      {stage2_3[73]}
   );
   gpc1_1 gpc2905 (
      {stage1_3[174]},
      {stage2_3[74]}
   );
   gpc1_1 gpc2906 (
      {stage1_3[175]},
      {stage2_3[75]}
   );
   gpc1_1 gpc2907 (
      {stage1_3[176]},
      {stage2_3[76]}
   );
   gpc1_1 gpc2908 (
      {stage1_3[177]},
      {stage2_3[77]}
   );
   gpc1_1 gpc2909 (
      {stage1_3[178]},
      {stage2_3[78]}
   );
   gpc1_1 gpc2910 (
      {stage1_3[179]},
      {stage2_3[79]}
   );
   gpc1_1 gpc2911 (
      {stage1_3[180]},
      {stage2_3[80]}
   );
   gpc1_1 gpc2912 (
      {stage1_3[181]},
      {stage2_3[81]}
   );
   gpc1_1 gpc2913 (
      {stage1_3[182]},
      {stage2_3[82]}
   );
   gpc1_1 gpc2914 (
      {stage1_3[183]},
      {stage2_3[83]}
   );
   gpc1_1 gpc2915 (
      {stage1_3[184]},
      {stage2_3[84]}
   );
   gpc1_1 gpc2916 (
      {stage1_3[185]},
      {stage2_3[85]}
   );
   gpc1_1 gpc2917 (
      {stage1_3[186]},
      {stage2_3[86]}
   );
   gpc1_1 gpc2918 (
      {stage1_3[187]},
      {stage2_3[87]}
   );
   gpc1_1 gpc2919 (
      {stage1_5[213]},
      {stage2_5[79]}
   );
   gpc1_1 gpc2920 (
      {stage1_5[214]},
      {stage2_5[80]}
   );
   gpc1_1 gpc2921 (
      {stage1_5[215]},
      {stage2_5[81]}
   );
   gpc1_1 gpc2922 (
      {stage1_5[216]},
      {stage2_5[82]}
   );
   gpc1_1 gpc2923 (
      {stage1_5[217]},
      {stage2_5[83]}
   );
   gpc1_1 gpc2924 (
      {stage1_7[218]},
      {stage2_7[104]}
   );
   gpc1_1 gpc2925 (
      {stage1_7[219]},
      {stage2_7[105]}
   );
   gpc1_1 gpc2926 (
      {stage1_7[220]},
      {stage2_7[106]}
   );
   gpc1_1 gpc2927 (
      {stage1_7[221]},
      {stage2_7[107]}
   );
   gpc1_1 gpc2928 (
      {stage1_7[222]},
      {stage2_7[108]}
   );
   gpc1_1 gpc2929 (
      {stage1_7[223]},
      {stage2_7[109]}
   );
   gpc1_1 gpc2930 (
      {stage1_8[183]},
      {stage2_8[85]}
   );
   gpc1_1 gpc2931 (
      {stage1_8[184]},
      {stage2_8[86]}
   );
   gpc1_1 gpc2932 (
      {stage1_8[185]},
      {stage2_8[87]}
   );
   gpc1_1 gpc2933 (
      {stage1_8[186]},
      {stage2_8[88]}
   );
   gpc1_1 gpc2934 (
      {stage1_8[187]},
      {stage2_8[89]}
   );
   gpc1_1 gpc2935 (
      {stage1_8[188]},
      {stage2_8[90]}
   );
   gpc1_1 gpc2936 (
      {stage1_8[189]},
      {stage2_8[91]}
   );
   gpc1_1 gpc2937 (
      {stage1_8[190]},
      {stage2_8[92]}
   );
   gpc1_1 gpc2938 (
      {stage1_8[191]},
      {stage2_8[93]}
   );
   gpc1_1 gpc2939 (
      {stage1_8[192]},
      {stage2_8[94]}
   );
   gpc1_1 gpc2940 (
      {stage1_8[193]},
      {stage2_8[95]}
   );
   gpc1_1 gpc2941 (
      {stage1_8[194]},
      {stage2_8[96]}
   );
   gpc1_1 gpc2942 (
      {stage1_8[195]},
      {stage2_8[97]}
   );
   gpc1_1 gpc2943 (
      {stage1_8[196]},
      {stage2_8[98]}
   );
   gpc1_1 gpc2944 (
      {stage1_8[197]},
      {stage2_8[99]}
   );
   gpc1_1 gpc2945 (
      {stage1_8[198]},
      {stage2_8[100]}
   );
   gpc1_1 gpc2946 (
      {stage1_8[199]},
      {stage2_8[101]}
   );
   gpc1_1 gpc2947 (
      {stage1_8[200]},
      {stage2_8[102]}
   );
   gpc1_1 gpc2948 (
      {stage1_8[201]},
      {stage2_8[103]}
   );
   gpc1_1 gpc2949 (
      {stage1_8[202]},
      {stage2_8[104]}
   );
   gpc1_1 gpc2950 (
      {stage1_8[203]},
      {stage2_8[105]}
   );
   gpc1_1 gpc2951 (
      {stage1_8[204]},
      {stage2_8[106]}
   );
   gpc1_1 gpc2952 (
      {stage1_8[205]},
      {stage2_8[107]}
   );
   gpc1_1 gpc2953 (
      {stage1_9[211]},
      {stage2_9[72]}
   );
   gpc1_1 gpc2954 (
      {stage1_9[212]},
      {stage2_9[73]}
   );
   gpc1_1 gpc2955 (
      {stage1_9[213]},
      {stage2_9[74]}
   );
   gpc1_1 gpc2956 (
      {stage1_10[186]},
      {stage2_10[87]}
   );
   gpc1_1 gpc2957 (
      {stage1_10[187]},
      {stage2_10[88]}
   );
   gpc1_1 gpc2958 (
      {stage1_12[277]},
      {stage2_12[98]}
   );
   gpc1_1 gpc2959 (
      {stage1_12[278]},
      {stage2_12[99]}
   );
   gpc1_1 gpc2960 (
      {stage1_12[279]},
      {stage2_12[100]}
   );
   gpc1_1 gpc2961 (
      {stage1_12[280]},
      {stage2_12[101]}
   );
   gpc1_1 gpc2962 (
      {stage1_12[281]},
      {stage2_12[102]}
   );
   gpc1_1 gpc2963 (
      {stage1_14[238]},
      {stage2_14[80]}
   );
   gpc1_1 gpc2964 (
      {stage1_14[239]},
      {stage2_14[81]}
   );
   gpc1_1 gpc2965 (
      {stage1_14[240]},
      {stage2_14[82]}
   );
   gpc1_1 gpc2966 (
      {stage1_14[241]},
      {stage2_14[83]}
   );
   gpc1_1 gpc2967 (
      {stage1_14[242]},
      {stage2_14[84]}
   );
   gpc1_1 gpc2968 (
      {stage1_14[243]},
      {stage2_14[85]}
   );
   gpc1_1 gpc2969 (
      {stage1_14[244]},
      {stage2_14[86]}
   );
   gpc1_1 gpc2970 (
      {stage1_14[245]},
      {stage2_14[87]}
   );
   gpc1_1 gpc2971 (
      {stage1_14[246]},
      {stage2_14[88]}
   );
   gpc1_1 gpc2972 (
      {stage1_14[247]},
      {stage2_14[89]}
   );
   gpc1_1 gpc2973 (
      {stage1_14[248]},
      {stage2_14[90]}
   );
   gpc1_1 gpc2974 (
      {stage1_14[249]},
      {stage2_14[91]}
   );
   gpc1_1 gpc2975 (
      {stage1_14[250]},
      {stage2_14[92]}
   );
   gpc1_1 gpc2976 (
      {stage1_14[251]},
      {stage2_14[93]}
   );
   gpc1_1 gpc2977 (
      {stage1_14[252]},
      {stage2_14[94]}
   );
   gpc1_1 gpc2978 (
      {stage1_14[253]},
      {stage2_14[95]}
   );
   gpc1_1 gpc2979 (
      {stage1_14[254]},
      {stage2_14[96]}
   );
   gpc1_1 gpc2980 (
      {stage1_14[255]},
      {stage2_14[97]}
   );
   gpc1_1 gpc2981 (
      {stage1_14[256]},
      {stage2_14[98]}
   );
   gpc1_1 gpc2982 (
      {stage1_14[257]},
      {stage2_14[99]}
   );
   gpc1_1 gpc2983 (
      {stage1_14[258]},
      {stage2_14[100]}
   );
   gpc1_1 gpc2984 (
      {stage1_14[259]},
      {stage2_14[101]}
   );
   gpc1_1 gpc2985 (
      {stage1_14[260]},
      {stage2_14[102]}
   );
   gpc1_1 gpc2986 (
      {stage1_14[261]},
      {stage2_14[103]}
   );
   gpc1_1 gpc2987 (
      {stage1_14[262]},
      {stage2_14[104]}
   );
   gpc1_1 gpc2988 (
      {stage1_14[263]},
      {stage2_14[105]}
   );
   gpc1_1 gpc2989 (
      {stage1_14[264]},
      {stage2_14[106]}
   );
   gpc1_1 gpc2990 (
      {stage1_14[265]},
      {stage2_14[107]}
   );
   gpc1_1 gpc2991 (
      {stage1_14[266]},
      {stage2_14[108]}
   );
   gpc1_1 gpc2992 (
      {stage1_14[267]},
      {stage2_14[109]}
   );
   gpc1_1 gpc2993 (
      {stage1_14[268]},
      {stage2_14[110]}
   );
   gpc1_1 gpc2994 (
      {stage1_14[269]},
      {stage2_14[111]}
   );
   gpc1_1 gpc2995 (
      {stage1_14[270]},
      {stage2_14[112]}
   );
   gpc1_1 gpc2996 (
      {stage1_14[271]},
      {stage2_14[113]}
   );
   gpc1_1 gpc2997 (
      {stage1_14[272]},
      {stage2_14[114]}
   );
   gpc1_1 gpc2998 (
      {stage1_14[273]},
      {stage2_14[115]}
   );
   gpc1_1 gpc2999 (
      {stage1_14[274]},
      {stage2_14[116]}
   );
   gpc1_1 gpc3000 (
      {stage1_14[275]},
      {stage2_14[117]}
   );
   gpc1_1 gpc3001 (
      {stage1_14[276]},
      {stage2_14[118]}
   );
   gpc1_1 gpc3002 (
      {stage1_14[277]},
      {stage2_14[119]}
   );
   gpc1_1 gpc3003 (
      {stage1_14[278]},
      {stage2_14[120]}
   );
   gpc1_1 gpc3004 (
      {stage1_14[279]},
      {stage2_14[121]}
   );
   gpc1_1 gpc3005 (
      {stage1_14[280]},
      {stage2_14[122]}
   );
   gpc1_1 gpc3006 (
      {stage1_14[281]},
      {stage2_14[123]}
   );
   gpc1_1 gpc3007 (
      {stage1_14[282]},
      {stage2_14[124]}
   );
   gpc1_1 gpc3008 (
      {stage1_14[283]},
      {stage2_14[125]}
   );
   gpc1_1 gpc3009 (
      {stage1_14[284]},
      {stage2_14[126]}
   );
   gpc1_1 gpc3010 (
      {stage1_14[285]},
      {stage2_14[127]}
   );
   gpc1_1 gpc3011 (
      {stage1_14[286]},
      {stage2_14[128]}
   );
   gpc1_1 gpc3012 (
      {stage1_14[287]},
      {stage2_14[129]}
   );
   gpc1_1 gpc3013 (
      {stage1_14[288]},
      {stage2_14[130]}
   );
   gpc1_1 gpc3014 (
      {stage1_14[289]},
      {stage2_14[131]}
   );
   gpc1_1 gpc3015 (
      {stage1_14[290]},
      {stage2_14[132]}
   );
   gpc1_1 gpc3016 (
      {stage1_14[291]},
      {stage2_14[133]}
   );
   gpc1_1 gpc3017 (
      {stage1_14[292]},
      {stage2_14[134]}
   );
   gpc1_1 gpc3018 (
      {stage1_14[293]},
      {stage2_14[135]}
   );
   gpc1_1 gpc3019 (
      {stage1_14[294]},
      {stage2_14[136]}
   );
   gpc1_1 gpc3020 (
      {stage1_14[295]},
      {stage2_14[137]}
   );
   gpc1_1 gpc3021 (
      {stage1_14[296]},
      {stage2_14[138]}
   );
   gpc1_1 gpc3022 (
      {stage1_15[128]},
      {stage2_15[92]}
   );
   gpc1_1 gpc3023 (
      {stage1_15[129]},
      {stage2_15[93]}
   );
   gpc1_1 gpc3024 (
      {stage1_15[130]},
      {stage2_15[94]}
   );
   gpc1_1 gpc3025 (
      {stage1_15[131]},
      {stage2_15[95]}
   );
   gpc1_1 gpc3026 (
      {stage1_15[132]},
      {stage2_15[96]}
   );
   gpc1_1 gpc3027 (
      {stage1_15[133]},
      {stage2_15[97]}
   );
   gpc1_1 gpc3028 (
      {stage1_15[134]},
      {stage2_15[98]}
   );
   gpc1_1 gpc3029 (
      {stage1_15[135]},
      {stage2_15[99]}
   );
   gpc1_1 gpc3030 (
      {stage1_15[136]},
      {stage2_15[100]}
   );
   gpc1_1 gpc3031 (
      {stage1_15[137]},
      {stage2_15[101]}
   );
   gpc1_1 gpc3032 (
      {stage1_15[138]},
      {stage2_15[102]}
   );
   gpc1_1 gpc3033 (
      {stage1_15[139]},
      {stage2_15[103]}
   );
   gpc1_1 gpc3034 (
      {stage1_15[140]},
      {stage2_15[104]}
   );
   gpc1_1 gpc3035 (
      {stage1_15[141]},
      {stage2_15[105]}
   );
   gpc1_1 gpc3036 (
      {stage1_15[142]},
      {stage2_15[106]}
   );
   gpc1_1 gpc3037 (
      {stage1_15[143]},
      {stage2_15[107]}
   );
   gpc1_1 gpc3038 (
      {stage1_15[144]},
      {stage2_15[108]}
   );
   gpc1_1 gpc3039 (
      {stage1_15[145]},
      {stage2_15[109]}
   );
   gpc1_1 gpc3040 (
      {stage1_15[146]},
      {stage2_15[110]}
   );
   gpc1_1 gpc3041 (
      {stage1_15[147]},
      {stage2_15[111]}
   );
   gpc1_1 gpc3042 (
      {stage1_15[148]},
      {stage2_15[112]}
   );
   gpc1_1 gpc3043 (
      {stage1_15[149]},
      {stage2_15[113]}
   );
   gpc1_1 gpc3044 (
      {stage1_15[150]},
      {stage2_15[114]}
   );
   gpc1_1 gpc3045 (
      {stage1_15[151]},
      {stage2_15[115]}
   );
   gpc1_1 gpc3046 (
      {stage1_15[152]},
      {stage2_15[116]}
   );
   gpc1_1 gpc3047 (
      {stage1_15[153]},
      {stage2_15[117]}
   );
   gpc1_1 gpc3048 (
      {stage1_15[154]},
      {stage2_15[118]}
   );
   gpc1_1 gpc3049 (
      {stage1_15[155]},
      {stage2_15[119]}
   );
   gpc1_1 gpc3050 (
      {stage1_15[156]},
      {stage2_15[120]}
   );
   gpc1_1 gpc3051 (
      {stage1_15[157]},
      {stage2_15[121]}
   );
   gpc1_1 gpc3052 (
      {stage1_15[158]},
      {stage2_15[122]}
   );
   gpc1_1 gpc3053 (
      {stage1_15[159]},
      {stage2_15[123]}
   );
   gpc1_1 gpc3054 (
      {stage1_15[160]},
      {stage2_15[124]}
   );
   gpc1_1 gpc3055 (
      {stage1_15[161]},
      {stage2_15[125]}
   );
   gpc1_1 gpc3056 (
      {stage1_15[162]},
      {stage2_15[126]}
   );
   gpc1_1 gpc3057 (
      {stage1_15[163]},
      {stage2_15[127]}
   );
   gpc1_1 gpc3058 (
      {stage1_15[164]},
      {stage2_15[128]}
   );
   gpc1_1 gpc3059 (
      {stage1_15[165]},
      {stage2_15[129]}
   );
   gpc1_1 gpc3060 (
      {stage1_15[166]},
      {stage2_15[130]}
   );
   gpc1_1 gpc3061 (
      {stage1_15[167]},
      {stage2_15[131]}
   );
   gpc1_1 gpc3062 (
      {stage1_15[168]},
      {stage2_15[132]}
   );
   gpc1_1 gpc3063 (
      {stage1_15[169]},
      {stage2_15[133]}
   );
   gpc1_1 gpc3064 (
      {stage1_15[170]},
      {stage2_15[134]}
   );
   gpc1_1 gpc3065 (
      {stage1_15[171]},
      {stage2_15[135]}
   );
   gpc1_1 gpc3066 (
      {stage1_16[257]},
      {stage2_16[96]}
   );
   gpc1_1 gpc3067 (
      {stage1_16[258]},
      {stage2_16[97]}
   );
   gpc1_1 gpc3068 (
      {stage1_16[259]},
      {stage2_16[98]}
   );
   gpc1_1 gpc3069 (
      {stage1_16[260]},
      {stage2_16[99]}
   );
   gpc1_1 gpc3070 (
      {stage1_16[261]},
      {stage2_16[100]}
   );
   gpc1_1 gpc3071 (
      {stage1_16[262]},
      {stage2_16[101]}
   );
   gpc1_1 gpc3072 (
      {stage1_16[263]},
      {stage2_16[102]}
   );
   gpc1_1 gpc3073 (
      {stage1_16[264]},
      {stage2_16[103]}
   );
   gpc1_1 gpc3074 (
      {stage1_17[234]},
      {stage2_17[85]}
   );
   gpc1_1 gpc3075 (
      {stage1_17[235]},
      {stage2_17[86]}
   );
   gpc1_1 gpc3076 (
      {stage1_17[236]},
      {stage2_17[87]}
   );
   gpc1_1 gpc3077 (
      {stage1_17[237]},
      {stage2_17[88]}
   );
   gpc1_1 gpc3078 (
      {stage1_17[238]},
      {stage2_17[89]}
   );
   gpc1_1 gpc3079 (
      {stage1_17[239]},
      {stage2_17[90]}
   );
   gpc1_1 gpc3080 (
      {stage1_17[240]},
      {stage2_17[91]}
   );
   gpc1_1 gpc3081 (
      {stage1_17[241]},
      {stage2_17[92]}
   );
   gpc1_1 gpc3082 (
      {stage1_17[242]},
      {stage2_17[93]}
   );
   gpc1_1 gpc3083 (
      {stage1_17[243]},
      {stage2_17[94]}
   );
   gpc1_1 gpc3084 (
      {stage1_17[244]},
      {stage2_17[95]}
   );
   gpc1_1 gpc3085 (
      {stage1_17[245]},
      {stage2_17[96]}
   );
   gpc1_1 gpc3086 (
      {stage1_17[246]},
      {stage2_17[97]}
   );
   gpc1_1 gpc3087 (
      {stage1_17[247]},
      {stage2_17[98]}
   );
   gpc1_1 gpc3088 (
      {stage1_17[248]},
      {stage2_17[99]}
   );
   gpc1_1 gpc3089 (
      {stage1_17[249]},
      {stage2_17[100]}
   );
   gpc1_1 gpc3090 (
      {stage1_17[250]},
      {stage2_17[101]}
   );
   gpc1_1 gpc3091 (
      {stage1_17[251]},
      {stage2_17[102]}
   );
   gpc1_1 gpc3092 (
      {stage1_17[252]},
      {stage2_17[103]}
   );
   gpc1_1 gpc3093 (
      {stage1_17[253]},
      {stage2_17[104]}
   );
   gpc1_1 gpc3094 (
      {stage1_17[254]},
      {stage2_17[105]}
   );
   gpc1_1 gpc3095 (
      {stage1_17[255]},
      {stage2_17[106]}
   );
   gpc1_1 gpc3096 (
      {stage1_17[256]},
      {stage2_17[107]}
   );
   gpc1_1 gpc3097 (
      {stage1_17[257]},
      {stage2_17[108]}
   );
   gpc1_1 gpc3098 (
      {stage1_17[258]},
      {stage2_17[109]}
   );
   gpc1_1 gpc3099 (
      {stage1_17[259]},
      {stage2_17[110]}
   );
   gpc1_1 gpc3100 (
      {stage1_17[260]},
      {stage2_17[111]}
   );
   gpc1_1 gpc3101 (
      {stage1_17[261]},
      {stage2_17[112]}
   );
   gpc1_1 gpc3102 (
      {stage1_17[262]},
      {stage2_17[113]}
   );
   gpc1_1 gpc3103 (
      {stage1_17[263]},
      {stage2_17[114]}
   );
   gpc1_1 gpc3104 (
      {stage1_17[264]},
      {stage2_17[115]}
   );
   gpc1_1 gpc3105 (
      {stage1_17[265]},
      {stage2_17[116]}
   );
   gpc1_1 gpc3106 (
      {stage1_17[266]},
      {stage2_17[117]}
   );
   gpc1_1 gpc3107 (
      {stage1_17[267]},
      {stage2_17[118]}
   );
   gpc1_1 gpc3108 (
      {stage1_17[268]},
      {stage2_17[119]}
   );
   gpc1_1 gpc3109 (
      {stage1_17[269]},
      {stage2_17[120]}
   );
   gpc1_1 gpc3110 (
      {stage1_17[270]},
      {stage2_17[121]}
   );
   gpc1_1 gpc3111 (
      {stage1_18[198]},
      {stage2_18[79]}
   );
   gpc1_1 gpc3112 (
      {stage1_18[199]},
      {stage2_18[80]}
   );
   gpc1_1 gpc3113 (
      {stage1_18[200]},
      {stage2_18[81]}
   );
   gpc1_1 gpc3114 (
      {stage1_19[295]},
      {stage2_19[105]}
   );
   gpc1_1 gpc3115 (
      {stage1_19[296]},
      {stage2_19[106]}
   );
   gpc1_1 gpc3116 (
      {stage1_19[297]},
      {stage2_19[107]}
   );
   gpc1_1 gpc3117 (
      {stage1_19[298]},
      {stage2_19[108]}
   );
   gpc1_1 gpc3118 (
      {stage1_19[299]},
      {stage2_19[109]}
   );
   gpc1_1 gpc3119 (
      {stage1_20[172]},
      {stage2_20[111]}
   );
   gpc1_1 gpc3120 (
      {stage1_20[173]},
      {stage2_20[112]}
   );
   gpc1_1 gpc3121 (
      {stage1_20[174]},
      {stage2_20[113]}
   );
   gpc1_1 gpc3122 (
      {stage1_20[175]},
      {stage2_20[114]}
   );
   gpc1_1 gpc3123 (
      {stage1_20[176]},
      {stage2_20[115]}
   );
   gpc1_1 gpc3124 (
      {stage1_20[177]},
      {stage2_20[116]}
   );
   gpc1_1 gpc3125 (
      {stage1_20[178]},
      {stage2_20[117]}
   );
   gpc1_1 gpc3126 (
      {stage1_20[179]},
      {stage2_20[118]}
   );
   gpc1_1 gpc3127 (
      {stage1_20[180]},
      {stage2_20[119]}
   );
   gpc1_1 gpc3128 (
      {stage1_20[181]},
      {stage2_20[120]}
   );
   gpc1_1 gpc3129 (
      {stage1_20[182]},
      {stage2_20[121]}
   );
   gpc1_1 gpc3130 (
      {stage1_20[183]},
      {stage2_20[122]}
   );
   gpc1_1 gpc3131 (
      {stage1_20[184]},
      {stage2_20[123]}
   );
   gpc1_1 gpc3132 (
      {stage1_20[185]},
      {stage2_20[124]}
   );
   gpc1_1 gpc3133 (
      {stage1_20[186]},
      {stage2_20[125]}
   );
   gpc1_1 gpc3134 (
      {stage1_20[187]},
      {stage2_20[126]}
   );
   gpc1_1 gpc3135 (
      {stage1_20[188]},
      {stage2_20[127]}
   );
   gpc1_1 gpc3136 (
      {stage1_21[198]},
      {stage2_21[78]}
   );
   gpc1_1 gpc3137 (
      {stage1_24[194]},
      {stage2_24[82]}
   );
   gpc1_1 gpc3138 (
      {stage1_24[195]},
      {stage2_24[83]}
   );
   gpc1_1 gpc3139 (
      {stage1_24[196]},
      {stage2_24[84]}
   );
   gpc1_1 gpc3140 (
      {stage1_24[197]},
      {stage2_24[85]}
   );
   gpc1_1 gpc3141 (
      {stage1_24[198]},
      {stage2_24[86]}
   );
   gpc1_1 gpc3142 (
      {stage1_24[199]},
      {stage2_24[87]}
   );
   gpc1_1 gpc3143 (
      {stage1_24[200]},
      {stage2_24[88]}
   );
   gpc1_1 gpc3144 (
      {stage1_24[201]},
      {stage2_24[89]}
   );
   gpc1_1 gpc3145 (
      {stage1_24[202]},
      {stage2_24[90]}
   );
   gpc1_1 gpc3146 (
      {stage1_24[203]},
      {stage2_24[91]}
   );
   gpc1_1 gpc3147 (
      {stage1_24[204]},
      {stage2_24[92]}
   );
   gpc1_1 gpc3148 (
      {stage1_24[205]},
      {stage2_24[93]}
   );
   gpc1_1 gpc3149 (
      {stage1_24[206]},
      {stage2_24[94]}
   );
   gpc1_1 gpc3150 (
      {stage1_24[207]},
      {stage2_24[95]}
   );
   gpc1_1 gpc3151 (
      {stage1_24[208]},
      {stage2_24[96]}
   );
   gpc1_1 gpc3152 (
      {stage1_24[209]},
      {stage2_24[97]}
   );
   gpc1_1 gpc3153 (
      {stage1_24[210]},
      {stage2_24[98]}
   );
   gpc1_1 gpc3154 (
      {stage1_24[211]},
      {stage2_24[99]}
   );
   gpc1_1 gpc3155 (
      {stage1_25[209]},
      {stage2_25[62]}
   );
   gpc1_1 gpc3156 (
      {stage1_25[210]},
      {stage2_25[63]}
   );
   gpc1_1 gpc3157 (
      {stage1_25[211]},
      {stage2_25[64]}
   );
   gpc1_1 gpc3158 (
      {stage1_25[212]},
      {stage2_25[65]}
   );
   gpc1_1 gpc3159 (
      {stage1_25[213]},
      {stage2_25[66]}
   );
   gpc1_1 gpc3160 (
      {stage1_25[214]},
      {stage2_25[67]}
   );
   gpc1_1 gpc3161 (
      {stage1_25[215]},
      {stage2_25[68]}
   );
   gpc1_1 gpc3162 (
      {stage1_25[216]},
      {stage2_25[69]}
   );
   gpc1_1 gpc3163 (
      {stage1_25[217]},
      {stage2_25[70]}
   );
   gpc1_1 gpc3164 (
      {stage1_25[218]},
      {stage2_25[71]}
   );
   gpc1_1 gpc3165 (
      {stage1_25[219]},
      {stage2_25[72]}
   );
   gpc1_1 gpc3166 (
      {stage1_25[220]},
      {stage2_25[73]}
   );
   gpc1_1 gpc3167 (
      {stage1_25[221]},
      {stage2_25[74]}
   );
   gpc1_1 gpc3168 (
      {stage1_25[222]},
      {stage2_25[75]}
   );
   gpc1_1 gpc3169 (
      {stage1_25[223]},
      {stage2_25[76]}
   );
   gpc1_1 gpc3170 (
      {stage1_25[224]},
      {stage2_25[77]}
   );
   gpc1_1 gpc3171 (
      {stage1_25[225]},
      {stage2_25[78]}
   );
   gpc1_1 gpc3172 (
      {stage1_25[226]},
      {stage2_25[79]}
   );
   gpc1_1 gpc3173 (
      {stage1_25[227]},
      {stage2_25[80]}
   );
   gpc1_1 gpc3174 (
      {stage1_25[228]},
      {stage2_25[81]}
   );
   gpc1_1 gpc3175 (
      {stage1_25[229]},
      {stage2_25[82]}
   );
   gpc1_1 gpc3176 (
      {stage1_25[230]},
      {stage2_25[83]}
   );
   gpc1_1 gpc3177 (
      {stage1_25[231]},
      {stage2_25[84]}
   );
   gpc1_1 gpc3178 (
      {stage1_25[232]},
      {stage2_25[85]}
   );
   gpc1_1 gpc3179 (
      {stage1_25[233]},
      {stage2_25[86]}
   );
   gpc1_1 gpc3180 (
      {stage1_25[234]},
      {stage2_25[87]}
   );
   gpc1_1 gpc3181 (
      {stage1_28[243]},
      {stage2_28[66]}
   );
   gpc1_1 gpc3182 (
      {stage1_28[244]},
      {stage2_28[67]}
   );
   gpc1_1 gpc3183 (
      {stage1_28[245]},
      {stage2_28[68]}
   );
   gpc1_1 gpc3184 (
      {stage1_28[246]},
      {stage2_28[69]}
   );
   gpc1_1 gpc3185 (
      {stage1_28[247]},
      {stage2_28[70]}
   );
   gpc1_1 gpc3186 (
      {stage1_28[248]},
      {stage2_28[71]}
   );
   gpc1_1 gpc3187 (
      {stage1_28[249]},
      {stage2_28[72]}
   );
   gpc1_1 gpc3188 (
      {stage1_28[250]},
      {stage2_28[73]}
   );
   gpc1_1 gpc3189 (
      {stage1_28[251]},
      {stage2_28[74]}
   );
   gpc1_1 gpc3190 (
      {stage1_29[186]},
      {stage2_29[71]}
   );
   gpc1_1 gpc3191 (
      {stage1_29[187]},
      {stage2_29[72]}
   );
   gpc1_1 gpc3192 (
      {stage1_29[188]},
      {stage2_29[73]}
   );
   gpc1_1 gpc3193 (
      {stage1_29[189]},
      {stage2_29[74]}
   );
   gpc1_1 gpc3194 (
      {stage1_29[190]},
      {stage2_29[75]}
   );
   gpc1_1 gpc3195 (
      {stage1_29[191]},
      {stage2_29[76]}
   );
   gpc1_1 gpc3196 (
      {stage1_29[192]},
      {stage2_29[77]}
   );
   gpc1_1 gpc3197 (
      {stage1_29[193]},
      {stage2_29[78]}
   );
   gpc1_1 gpc3198 (
      {stage1_29[194]},
      {stage2_29[79]}
   );
   gpc1_1 gpc3199 (
      {stage1_29[195]},
      {stage2_29[80]}
   );
   gpc1_1 gpc3200 (
      {stage1_29[196]},
      {stage2_29[81]}
   );
   gpc1_1 gpc3201 (
      {stage1_29[197]},
      {stage2_29[82]}
   );
   gpc1_1 gpc3202 (
      {stage1_29[198]},
      {stage2_29[83]}
   );
   gpc1_1 gpc3203 (
      {stage1_29[199]},
      {stage2_29[84]}
   );
   gpc1_1 gpc3204 (
      {stage1_29[200]},
      {stage2_29[85]}
   );
   gpc1_1 gpc3205 (
      {stage1_29[201]},
      {stage2_29[86]}
   );
   gpc1_1 gpc3206 (
      {stage1_29[202]},
      {stage2_29[87]}
   );
   gpc1_1 gpc3207 (
      {stage1_29[203]},
      {stage2_29[88]}
   );
   gpc1_1 gpc3208 (
      {stage1_29[204]},
      {stage2_29[89]}
   );
   gpc1_1 gpc3209 (
      {stage1_29[205]},
      {stage2_29[90]}
   );
   gpc1_1 gpc3210 (
      {stage1_29[206]},
      {stage2_29[91]}
   );
   gpc1_1 gpc3211 (
      {stage1_29[207]},
      {stage2_29[92]}
   );
   gpc1_1 gpc3212 (
      {stage1_29[208]},
      {stage2_29[93]}
   );
   gpc1_1 gpc3213 (
      {stage1_29[209]},
      {stage2_29[94]}
   );
   gpc1_1 gpc3214 (
      {stage1_29[210]},
      {stage2_29[95]}
   );
   gpc1_1 gpc3215 (
      {stage1_29[211]},
      {stage2_29[96]}
   );
   gpc1_1 gpc3216 (
      {stage1_29[212]},
      {stage2_29[97]}
   );
   gpc1_1 gpc3217 (
      {stage1_29[213]},
      {stage2_29[98]}
   );
   gpc1_1 gpc3218 (
      {stage1_29[214]},
      {stage2_29[99]}
   );
   gpc1_1 gpc3219 (
      {stage1_29[215]},
      {stage2_29[100]}
   );
   gpc1_1 gpc3220 (
      {stage1_29[216]},
      {stage2_29[101]}
   );
   gpc1_1 gpc3221 (
      {stage1_29[217]},
      {stage2_29[102]}
   );
   gpc1_1 gpc3222 (
      {stage1_29[218]},
      {stage2_29[103]}
   );
   gpc1_1 gpc3223 (
      {stage1_29[219]},
      {stage2_29[104]}
   );
   gpc1_1 gpc3224 (
      {stage1_29[220]},
      {stage2_29[105]}
   );
   gpc1_1 gpc3225 (
      {stage1_29[221]},
      {stage2_29[106]}
   );
   gpc1_1 gpc3226 (
      {stage1_29[222]},
      {stage2_29[107]}
   );
   gpc1_1 gpc3227 (
      {stage1_29[223]},
      {stage2_29[108]}
   );
   gpc1_1 gpc3228 (
      {stage1_29[224]},
      {stage2_29[109]}
   );
   gpc1_1 gpc3229 (
      {stage1_29[225]},
      {stage2_29[110]}
   );
   gpc1_1 gpc3230 (
      {stage1_29[226]},
      {stage2_29[111]}
   );
   gpc1_1 gpc3231 (
      {stage1_29[227]},
      {stage2_29[112]}
   );
   gpc1_1 gpc3232 (
      {stage1_29[228]},
      {stage2_29[113]}
   );
   gpc1_1 gpc3233 (
      {stage1_29[229]},
      {stage2_29[114]}
   );
   gpc1_1 gpc3234 (
      {stage1_29[230]},
      {stage2_29[115]}
   );
   gpc1_1 gpc3235 (
      {stage1_29[231]},
      {stage2_29[116]}
   );
   gpc1_1 gpc3236 (
      {stage1_29[232]},
      {stage2_29[117]}
   );
   gpc1_1 gpc3237 (
      {stage1_29[233]},
      {stage2_29[118]}
   );
   gpc1_1 gpc3238 (
      {stage1_29[234]},
      {stage2_29[119]}
   );
   gpc1_1 gpc3239 (
      {stage1_29[235]},
      {stage2_29[120]}
   );
   gpc1_1 gpc3240 (
      {stage1_30[132]},
      {stage2_30[90]}
   );
   gpc1_1 gpc3241 (
      {stage1_30[133]},
      {stage2_30[91]}
   );
   gpc1_1 gpc3242 (
      {stage1_30[134]},
      {stage2_30[92]}
   );
   gpc1_1 gpc3243 (
      {stage1_30[135]},
      {stage2_30[93]}
   );
   gpc1_1 gpc3244 (
      {stage1_30[136]},
      {stage2_30[94]}
   );
   gpc1_1 gpc3245 (
      {stage1_30[137]},
      {stage2_30[95]}
   );
   gpc1_1 gpc3246 (
      {stage1_30[138]},
      {stage2_30[96]}
   );
   gpc1_1 gpc3247 (
      {stage1_30[139]},
      {stage2_30[97]}
   );
   gpc1_1 gpc3248 (
      {stage1_30[140]},
      {stage2_30[98]}
   );
   gpc1_1 gpc3249 (
      {stage1_30[141]},
      {stage2_30[99]}
   );
   gpc1_1 gpc3250 (
      {stage1_30[142]},
      {stage2_30[100]}
   );
   gpc1_1 gpc3251 (
      {stage1_30[143]},
      {stage2_30[101]}
   );
   gpc1_1 gpc3252 (
      {stage1_30[144]},
      {stage2_30[102]}
   );
   gpc1_1 gpc3253 (
      {stage1_30[145]},
      {stage2_30[103]}
   );
   gpc1_1 gpc3254 (
      {stage1_30[146]},
      {stage2_30[104]}
   );
   gpc1_1 gpc3255 (
      {stage1_30[147]},
      {stage2_30[105]}
   );
   gpc1_1 gpc3256 (
      {stage1_30[148]},
      {stage2_30[106]}
   );
   gpc1_1 gpc3257 (
      {stage1_30[149]},
      {stage2_30[107]}
   );
   gpc1_1 gpc3258 (
      {stage1_30[150]},
      {stage2_30[108]}
   );
   gpc1_1 gpc3259 (
      {stage1_30[151]},
      {stage2_30[109]}
   );
   gpc1_1 gpc3260 (
      {stage1_30[152]},
      {stage2_30[110]}
   );
   gpc1_1 gpc3261 (
      {stage1_30[153]},
      {stage2_30[111]}
   );
   gpc1_1 gpc3262 (
      {stage1_30[154]},
      {stage2_30[112]}
   );
   gpc1_1 gpc3263 (
      {stage1_30[155]},
      {stage2_30[113]}
   );
   gpc1_1 gpc3264 (
      {stage1_30[156]},
      {stage2_30[114]}
   );
   gpc1_1 gpc3265 (
      {stage1_30[157]},
      {stage2_30[115]}
   );
   gpc1_1 gpc3266 (
      {stage1_30[158]},
      {stage2_30[116]}
   );
   gpc1_1 gpc3267 (
      {stage1_30[159]},
      {stage2_30[117]}
   );
   gpc1_1 gpc3268 (
      {stage1_30[160]},
      {stage2_30[118]}
   );
   gpc1_1 gpc3269 (
      {stage1_30[161]},
      {stage2_30[119]}
   );
   gpc1_1 gpc3270 (
      {stage1_30[162]},
      {stage2_30[120]}
   );
   gpc1_1 gpc3271 (
      {stage1_30[163]},
      {stage2_30[121]}
   );
   gpc1_1 gpc3272 (
      {stage1_30[164]},
      {stage2_30[122]}
   );
   gpc1_1 gpc3273 (
      {stage1_30[165]},
      {stage2_30[123]}
   );
   gpc1_1 gpc3274 (
      {stage1_30[166]},
      {stage2_30[124]}
   );
   gpc1_1 gpc3275 (
      {stage1_30[167]},
      {stage2_30[125]}
   );
   gpc1_1 gpc3276 (
      {stage1_30[168]},
      {stage2_30[126]}
   );
   gpc1_1 gpc3277 (
      {stage1_30[169]},
      {stage2_30[127]}
   );
   gpc1_1 gpc3278 (
      {stage1_30[170]},
      {stage2_30[128]}
   );
   gpc1_1 gpc3279 (
      {stage1_30[171]},
      {stage2_30[129]}
   );
   gpc1_1 gpc3280 (
      {stage1_31[144]},
      {stage2_31[67]}
   );
   gpc1_1 gpc3281 (
      {stage1_31[145]},
      {stage2_31[68]}
   );
   gpc1_1 gpc3282 (
      {stage1_31[146]},
      {stage2_31[69]}
   );
   gpc1_1 gpc3283 (
      {stage1_31[147]},
      {stage2_31[70]}
   );
   gpc1_1 gpc3284 (
      {stage1_31[148]},
      {stage2_31[71]}
   );
   gpc1_1 gpc3285 (
      {stage1_31[149]},
      {stage2_31[72]}
   );
   gpc1_1 gpc3286 (
      {stage1_31[150]},
      {stage2_31[73]}
   );
   gpc1_1 gpc3287 (
      {stage1_31[151]},
      {stage2_31[74]}
   );
   gpc1_1 gpc3288 (
      {stage1_31[152]},
      {stage2_31[75]}
   );
   gpc1_1 gpc3289 (
      {stage1_31[153]},
      {stage2_31[76]}
   );
   gpc1_1 gpc3290 (
      {stage1_31[154]},
      {stage2_31[77]}
   );
   gpc1_1 gpc3291 (
      {stage1_31[155]},
      {stage2_31[78]}
   );
   gpc1_1 gpc3292 (
      {stage1_31[156]},
      {stage2_31[79]}
   );
   gpc1_1 gpc3293 (
      {stage1_31[157]},
      {stage2_31[80]}
   );
   gpc1_1 gpc3294 (
      {stage1_31[158]},
      {stage2_31[81]}
   );
   gpc1_1 gpc3295 (
      {stage1_31[159]},
      {stage2_31[82]}
   );
   gpc1_1 gpc3296 (
      {stage1_31[160]},
      {stage2_31[83]}
   );
   gpc1_1 gpc3297 (
      {stage1_32[132]},
      {stage2_32[46]}
   );
   gpc1_1 gpc3298 (
      {stage1_32[133]},
      {stage2_32[47]}
   );
   gpc1_1 gpc3299 (
      {stage1_32[134]},
      {stage2_32[48]}
   );
   gpc1_1 gpc3300 (
      {stage1_32[135]},
      {stage2_32[49]}
   );
   gpc1_1 gpc3301 (
      {stage1_32[136]},
      {stage2_32[50]}
   );
   gpc1_1 gpc3302 (
      {stage1_32[137]},
      {stage2_32[51]}
   );
   gpc1_1 gpc3303 (
      {stage1_32[138]},
      {stage2_32[52]}
   );
   gpc1_1 gpc3304 (
      {stage1_32[139]},
      {stage2_32[53]}
   );
   gpc1_1 gpc3305 (
      {stage1_32[140]},
      {stage2_32[54]}
   );
   gpc1_1 gpc3306 (
      {stage1_32[141]},
      {stage2_32[55]}
   );
   gpc1_1 gpc3307 (
      {stage1_32[142]},
      {stage2_32[56]}
   );
   gpc1_1 gpc3308 (
      {stage1_32[143]},
      {stage2_32[57]}
   );
   gpc1_1 gpc3309 (
      {stage1_32[144]},
      {stage2_32[58]}
   );
   gpc1_1 gpc3310 (
      {stage1_32[145]},
      {stage2_32[59]}
   );
   gpc1_1 gpc3311 (
      {stage1_32[146]},
      {stage2_32[60]}
   );
   gpc1_1 gpc3312 (
      {stage1_32[147]},
      {stage2_32[61]}
   );
   gpc1_1 gpc3313 (
      {stage1_32[148]},
      {stage2_32[62]}
   );
   gpc1_1 gpc3314 (
      {stage1_32[149]},
      {stage2_32[63]}
   );
   gpc1_1 gpc3315 (
      {stage1_32[150]},
      {stage2_32[64]}
   );
   gpc1163_5 gpc3316 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc3317 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1163_5 gpc3318 (
      {stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_2[2]},
      {stage2_3[2]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc1163_5 gpc3319 (
      {stage2_0[9], stage2_0[10], stage2_0[11]},
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_2[3]},
      {stage2_3[3]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc1163_5 gpc3320 (
      {stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_2[4]},
      {stage2_3[4]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc1163_5 gpc3321 (
      {stage2_0[15], stage2_0[16], stage2_0[17]},
      {stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35]},
      {stage2_2[5]},
      {stage2_3[5]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc1163_5 gpc3322 (
      {stage2_0[18], stage2_0[19], stage2_0[20]},
      {stage2_1[36], stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_2[6]},
      {stage2_3[6]},
      {stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6],stage3_0[6]}
   );
   gpc606_5 gpc3323 (
      {stage2_1[42], stage2_1[43], stage2_1[44], stage2_1[45], stage2_1[46], stage2_1[47]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[0],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc3324 (
      {stage2_1[48], stage2_1[49], stage2_1[50], stage2_1[51], stage2_1[52], stage2_1[53]},
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage3_5[1],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc3325 (
      {stage2_1[54], stage2_1[55], stage2_1[56], stage2_1[57], stage2_1[58], stage2_1[59]},
      {stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage3_5[2],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc606_5 gpc3326 (
      {stage2_1[60], stage2_1[61], stage2_1[62], stage2_1[63], stage2_1[64], stage2_1[65]},
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30]},
      {stage3_5[3],stage3_4[10],stage3_3[10],stage3_2[10],stage3_1[10]}
   );
   gpc606_5 gpc3327 (
      {stage2_1[66], stage2_1[67], stage2_1[68], stage2_1[69], stage2_1[70], stage2_1[71]},
      {stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35], stage2_3[36]},
      {stage3_5[4],stage3_4[11],stage3_3[11],stage3_2[11],stage3_1[11]}
   );
   gpc606_5 gpc3328 (
      {stage2_1[72], stage2_1[73], stage2_1[74], stage2_1[75], stage2_1[76], stage2_1[77]},
      {stage2_3[37], stage2_3[38], stage2_3[39], stage2_3[40], stage2_3[41], stage2_3[42]},
      {stage3_5[5],stage3_4[12],stage3_3[12],stage3_2[12],stage3_1[12]}
   );
   gpc606_5 gpc3329 (
      {stage2_1[78], stage2_1[79], stage2_1[80], stage2_1[81], stage2_1[82], stage2_1[83]},
      {stage2_3[43], stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48]},
      {stage3_5[6],stage3_4[13],stage3_3[13],stage3_2[13],stage3_1[13]}
   );
   gpc606_5 gpc3330 (
      {stage2_1[84], stage2_1[85], stage2_1[86], stage2_1[87], stage2_1[88], stage2_1[89]},
      {stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53], stage2_3[54]},
      {stage3_5[7],stage3_4[14],stage3_3[14],stage3_2[14],stage3_1[14]}
   );
   gpc606_5 gpc3331 (
      {stage2_1[90], stage2_1[91], stage2_1[92], stage2_1[93], stage2_1[94], stage2_1[95]},
      {stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58], stage2_3[59], stage2_3[60]},
      {stage3_5[8],stage3_4[15],stage3_3[15],stage3_2[15],stage3_1[15]}
   );
   gpc606_5 gpc3332 (
      {stage2_1[96], stage2_1[97], stage2_1[98], stage2_1[99], stage2_1[100], stage2_1[101]},
      {stage2_3[61], stage2_3[62], stage2_3[63], stage2_3[64], stage2_3[65], stage2_3[66]},
      {stage3_5[9],stage3_4[16],stage3_3[16],stage3_2[16],stage3_1[16]}
   );
   gpc606_5 gpc3333 (
      {stage2_1[102], stage2_1[103], stage2_1[104], stage2_1[105], stage2_1[106], 1'b0},
      {stage2_3[67], stage2_3[68], stage2_3[69], stage2_3[70], stage2_3[71], stage2_3[72]},
      {stage3_5[10],stage3_4[17],stage3_3[17],stage3_2[17],stage3_1[17]}
   );
   gpc606_5 gpc3334 (
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[11],stage3_4[18],stage3_3[18],stage3_2[18]}
   );
   gpc606_5 gpc3335 (
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[12],stage3_4[19],stage3_3[19],stage3_2[19]}
   );
   gpc606_5 gpc3336 (
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[13],stage3_4[20],stage3_3[20],stage3_2[20]}
   );
   gpc606_5 gpc3337 (
      {stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29], stage2_2[30]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[14],stage3_4[21],stage3_3[21],stage3_2[21]}
   );
   gpc606_5 gpc3338 (
      {stage2_2[31], stage2_2[32], stage2_2[33], stage2_2[34], stage2_2[35], stage2_2[36]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[15],stage3_4[22],stage3_3[22],stage3_2[22]}
   );
   gpc606_5 gpc3339 (
      {stage2_2[37], stage2_2[38], stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[16],stage3_4[23],stage3_3[23],stage3_2[23]}
   );
   gpc615_5 gpc3340 (
      {stage2_3[73], stage2_3[74], stage2_3[75], stage2_3[76], stage2_3[77]},
      {stage2_4[36]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[6],stage3_5[17],stage3_4[24],stage3_3[24]}
   );
   gpc615_5 gpc3341 (
      {stage2_3[78], stage2_3[79], stage2_3[80], stage2_3[81], stage2_3[82]},
      {stage2_4[37]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[7],stage3_5[18],stage3_4[25],stage3_3[25]}
   );
   gpc615_5 gpc3342 (
      {stage2_3[83], stage2_3[84], stage2_3[85], stage2_3[86], stage2_3[87]},
      {stage2_4[38]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[8],stage3_5[19],stage3_4[26],stage3_3[26]}
   );
   gpc606_5 gpc3343 (
      {stage2_4[39], stage2_4[40], stage2_4[41], stage2_4[42], stage2_4[43], stage2_4[44]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[9],stage3_5[20],stage3_4[27]}
   );
   gpc606_5 gpc3344 (
      {stage2_4[45], stage2_4[46], stage2_4[47], stage2_4[48], stage2_4[49], stage2_4[50]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[10],stage3_5[21],stage3_4[28]}
   );
   gpc606_5 gpc3345 (
      {stage2_4[51], stage2_4[52], stage2_4[53], stage2_4[54], stage2_4[55], stage2_4[56]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[11],stage3_5[22],stage3_4[29]}
   );
   gpc615_5 gpc3346 (
      {stage2_4[57], stage2_4[58], stage2_4[59], stage2_4[60], stage2_4[61]},
      {stage2_5[18]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[6],stage3_6[12],stage3_5[23],stage3_4[30]}
   );
   gpc615_5 gpc3347 (
      {stage2_4[62], stage2_4[63], stage2_4[64], stage2_4[65], stage2_4[66]},
      {stage2_5[19]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[7],stage3_6[13],stage3_5[24],stage3_4[31]}
   );
   gpc615_5 gpc3348 (
      {stage2_4[67], stage2_4[68], stage2_4[69], stage2_4[70], stage2_4[71]},
      {stage2_5[20]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[8],stage3_6[14],stage3_5[25],stage3_4[32]}
   );
   gpc615_5 gpc3349 (
      {stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75], stage2_4[76]},
      {stage2_5[21]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[9],stage3_6[15],stage3_5[26],stage3_4[33]}
   );
   gpc615_5 gpc3350 (
      {stage2_4[77], stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81]},
      {stage2_5[22]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[10],stage3_6[16],stage3_5[27],stage3_4[34]}
   );
   gpc606_5 gpc3351 (
      {stage2_5[23], stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[8],stage3_7[11],stage3_6[17],stage3_5[28]}
   );
   gpc606_5 gpc3352 (
      {stage2_5[29], stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[9],stage3_7[12],stage3_6[18],stage3_5[29]}
   );
   gpc606_5 gpc3353 (
      {stage2_5[35], stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[10],stage3_7[13],stage3_6[19],stage3_5[30]}
   );
   gpc606_5 gpc3354 (
      {stage2_5[41], stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[11],stage3_7[14],stage3_6[20],stage3_5[31]}
   );
   gpc606_5 gpc3355 (
      {stage2_5[47], stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[12],stage3_7[15],stage3_6[21],stage3_5[32]}
   );
   gpc606_5 gpc3356 (
      {stage2_5[53], stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58]},
      {stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35]},
      {stage3_9[5],stage3_8[13],stage3_7[16],stage3_6[22],stage3_5[33]}
   );
   gpc606_5 gpc3357 (
      {stage2_5[59], stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64]},
      {stage2_7[36], stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage3_9[6],stage3_8[14],stage3_7[17],stage3_6[23],stage3_5[34]}
   );
   gpc606_5 gpc3358 (
      {stage2_5[65], stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70]},
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46], stage2_7[47]},
      {stage3_9[7],stage3_8[15],stage3_7[18],stage3_6[24],stage3_5[35]}
   );
   gpc615_5 gpc3359 (
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52]},
      {stage2_7[48]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[8],stage3_8[16],stage3_7[19],stage3_6[25]}
   );
   gpc615_5 gpc3360 (
      {stage2_6[53], stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57]},
      {stage2_7[49]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[9],stage3_8[17],stage3_7[20],stage3_6[26]}
   );
   gpc615_5 gpc3361 (
      {stage2_6[58], stage2_6[59], stage2_6[60], stage2_6[61], stage2_6[62]},
      {stage2_7[50]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[10],stage3_8[18],stage3_7[21],stage3_6[27]}
   );
   gpc615_5 gpc3362 (
      {stage2_6[63], stage2_6[64], stage2_6[65], stage2_6[66], stage2_6[67]},
      {stage2_7[51]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[11],stage3_8[19],stage3_7[22],stage3_6[28]}
   );
   gpc615_5 gpc3363 (
      {stage2_6[68], stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72]},
      {stage2_7[52]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[12],stage3_8[20],stage3_7[23],stage3_6[29]}
   );
   gpc615_5 gpc3364 (
      {stage2_6[73], stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77]},
      {stage2_7[53]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[13],stage3_8[21],stage3_7[24],stage3_6[30]}
   );
   gpc615_5 gpc3365 (
      {stage2_6[78], stage2_6[79], stage2_6[80], stage2_6[81], stage2_6[82]},
      {stage2_7[54]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[14],stage3_8[22],stage3_7[25],stage3_6[31]}
   );
   gpc615_5 gpc3366 (
      {stage2_7[55], stage2_7[56], stage2_7[57], stage2_7[58], stage2_7[59]},
      {stage2_8[42]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[7],stage3_9[15],stage3_8[23],stage3_7[26]}
   );
   gpc615_5 gpc3367 (
      {stage2_7[60], stage2_7[61], stage2_7[62], stage2_7[63], stage2_7[64]},
      {stage2_8[43]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[8],stage3_9[16],stage3_8[24],stage3_7[27]}
   );
   gpc615_5 gpc3368 (
      {stage2_7[65], stage2_7[66], stage2_7[67], stage2_7[68], stage2_7[69]},
      {stage2_8[44]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[9],stage3_9[17],stage3_8[25],stage3_7[28]}
   );
   gpc1343_5 gpc3369 (
      {stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21]},
      {stage2_10[0], stage2_10[1], stage2_10[2]},
      {stage2_11[0]},
      {stage3_12[0],stage3_11[3],stage3_10[10],stage3_9[18],stage3_8[26]}
   );
   gpc1343_5 gpc3370 (
      {stage2_8[48], stage2_8[49], stage2_8[50]},
      {stage2_9[22], stage2_9[23], stage2_9[24], stage2_9[25]},
      {stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage2_11[1]},
      {stage3_12[1],stage3_11[4],stage3_10[11],stage3_9[19],stage3_8[27]}
   );
   gpc1343_5 gpc3371 (
      {stage2_8[51], stage2_8[52], stage2_8[53]},
      {stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage2_10[6], stage2_10[7], stage2_10[8]},
      {stage2_11[2]},
      {stage3_12[2],stage3_11[5],stage3_10[12],stage3_9[20],stage3_8[28]}
   );
   gpc606_5 gpc3372 (
      {stage2_8[54], stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59]},
      {stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12], stage2_10[13], stage2_10[14]},
      {stage3_12[3],stage3_11[6],stage3_10[13],stage3_9[21],stage3_8[29]}
   );
   gpc606_5 gpc3373 (
      {stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63], stage2_8[64], stage2_8[65]},
      {stage2_10[15], stage2_10[16], stage2_10[17], stage2_10[18], stage2_10[19], stage2_10[20]},
      {stage3_12[4],stage3_11[7],stage3_10[14],stage3_9[22],stage3_8[30]}
   );
   gpc606_5 gpc3374 (
      {stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70], stage2_8[71]},
      {stage2_10[21], stage2_10[22], stage2_10[23], stage2_10[24], stage2_10[25], stage2_10[26]},
      {stage3_12[5],stage3_11[8],stage3_10[15],stage3_9[23],stage3_8[31]}
   );
   gpc606_5 gpc3375 (
      {stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75], stage2_8[76], stage2_8[77]},
      {stage2_10[27], stage2_10[28], stage2_10[29], stage2_10[30], stage2_10[31], stage2_10[32]},
      {stage3_12[6],stage3_11[9],stage3_10[16],stage3_9[24],stage3_8[32]}
   );
   gpc606_5 gpc3376 (
      {stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81], stage2_8[82], stage2_8[83]},
      {stage2_10[33], stage2_10[34], stage2_10[35], stage2_10[36], stage2_10[37], stage2_10[38]},
      {stage3_12[7],stage3_11[10],stage3_10[17],stage3_9[25],stage3_8[33]}
   );
   gpc606_5 gpc3377 (
      {stage2_8[84], stage2_8[85], stage2_8[86], stage2_8[87], stage2_8[88], stage2_8[89]},
      {stage2_10[39], stage2_10[40], stage2_10[41], stage2_10[42], stage2_10[43], stage2_10[44]},
      {stage3_12[8],stage3_11[11],stage3_10[18],stage3_9[26],stage3_8[34]}
   );
   gpc606_5 gpc3378 (
      {stage2_8[90], stage2_8[91], stage2_8[92], stage2_8[93], stage2_8[94], stage2_8[95]},
      {stage2_10[45], stage2_10[46], stage2_10[47], stage2_10[48], stage2_10[49], stage2_10[50]},
      {stage3_12[9],stage3_11[12],stage3_10[19],stage3_9[27],stage3_8[35]}
   );
   gpc606_5 gpc3379 (
      {stage2_8[96], stage2_8[97], stage2_8[98], stage2_8[99], stage2_8[100], stage2_8[101]},
      {stage2_10[51], stage2_10[52], stage2_10[53], stage2_10[54], stage2_10[55], stage2_10[56]},
      {stage3_12[10],stage3_11[13],stage3_10[20],stage3_9[28],stage3_8[36]}
   );
   gpc606_5 gpc3380 (
      {stage2_8[102], stage2_8[103], stage2_8[104], stage2_8[105], stage2_8[106], stage2_8[107]},
      {stage2_10[57], stage2_10[58], stage2_10[59], stage2_10[60], stage2_10[61], stage2_10[62]},
      {stage3_12[11],stage3_11[14],stage3_10[21],stage3_9[29],stage3_8[37]}
   );
   gpc606_5 gpc3381 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8]},
      {stage3_13[0],stage3_12[12],stage3_11[15],stage3_10[22],stage3_9[30]}
   );
   gpc615_5 gpc3382 (
      {stage2_10[63], stage2_10[64], stage2_10[65], stage2_10[66], stage2_10[67]},
      {stage2_11[9]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[13],stage3_11[16],stage3_10[23]}
   );
   gpc615_5 gpc3383 (
      {stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71], stage2_10[72]},
      {stage2_11[10]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[2],stage3_12[14],stage3_11[17],stage3_10[24]}
   );
   gpc615_5 gpc3384 (
      {stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76], stage2_10[77]},
      {stage2_11[11]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[3],stage3_12[15],stage3_11[18],stage3_10[25]}
   );
   gpc615_5 gpc3385 (
      {stage2_10[78], stage2_10[79], stage2_10[80], stage2_10[81], stage2_10[82]},
      {stage2_11[12]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[3],stage3_13[4],stage3_12[16],stage3_11[19],stage3_10[26]}
   );
   gpc615_5 gpc3386 (
      {stage2_10[83], stage2_10[84], stage2_10[85], stage2_10[86], stage2_10[87]},
      {stage2_11[13]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[4],stage3_13[5],stage3_12[17],stage3_11[20],stage3_10[27]}
   );
   gpc606_5 gpc3387 (
      {stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[5],stage3_13[6],stage3_12[18],stage3_11[21]}
   );
   gpc606_5 gpc3388 (
      {stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[6],stage3_13[7],stage3_12[19],stage3_11[22]}
   );
   gpc606_5 gpc3389 (
      {stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[7],stage3_13[8],stage3_12[20],stage3_11[23]}
   );
   gpc606_5 gpc3390 (
      {stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[8],stage3_13[9],stage3_12[21],stage3_11[24]}
   );
   gpc606_5 gpc3391 (
      {stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[9],stage3_13[10],stage3_12[22],stage3_11[25]}
   );
   gpc606_5 gpc3392 (
      {stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48], stage2_11[49]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[10],stage3_13[11],stage3_12[23],stage3_11[26]}
   );
   gpc606_5 gpc3393 (
      {stage2_11[50], stage2_11[51], stage2_11[52], stage2_11[53], stage2_11[54], stage2_11[55]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[11],stage3_13[12],stage3_12[24],stage3_11[27]}
   );
   gpc606_5 gpc3394 (
      {stage2_11[56], stage2_11[57], stage2_11[58], stage2_11[59], stage2_11[60], stage2_11[61]},
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage3_15[7],stage3_14[12],stage3_13[13],stage3_12[25],stage3_11[28]}
   );
   gpc606_5 gpc3395 (
      {stage2_11[62], stage2_11[63], stage2_11[64], stage2_11[65], stage2_11[66], stage2_11[67]},
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage3_15[8],stage3_14[13],stage3_13[14],stage3_12[26],stage3_11[29]}
   );
   gpc606_5 gpc3396 (
      {stage2_11[68], stage2_11[69], stage2_11[70], stage2_11[71], stage2_11[72], stage2_11[73]},
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage3_15[9],stage3_14[14],stage3_13[15],stage3_12[27],stage3_11[30]}
   );
   gpc606_5 gpc3397 (
      {stage2_11[74], stage2_11[75], stage2_11[76], stage2_11[77], stage2_11[78], stage2_11[79]},
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage3_15[10],stage3_14[15],stage3_13[16],stage3_12[28],stage3_11[31]}
   );
   gpc606_5 gpc3398 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[11],stage3_14[16],stage3_13[17],stage3_12[29]}
   );
   gpc606_5 gpc3399 (
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[12],stage3_14[17],stage3_13[18],stage3_12[30]}
   );
   gpc606_5 gpc3400 (
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[13],stage3_14[18],stage3_13[19],stage3_12[31]}
   );
   gpc606_5 gpc3401 (
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[14],stage3_14[19],stage3_13[20],stage3_12[32]}
   );
   gpc606_5 gpc3402 (
      {stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[15],stage3_14[20],stage3_13[21],stage3_12[33]}
   );
   gpc606_5 gpc3403 (
      {stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[16],stage3_14[21],stage3_13[22],stage3_12[34]}
   );
   gpc606_5 gpc3404 (
      {stage2_12[66], stage2_12[67], stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[17],stage3_14[22],stage3_13[23],stage3_12[35]}
   );
   gpc606_5 gpc3405 (
      {stage2_12[72], stage2_12[73], stage2_12[74], stage2_12[75], stage2_12[76], stage2_12[77]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[18],stage3_14[23],stage3_13[24],stage3_12[36]}
   );
   gpc606_5 gpc3406 (
      {stage2_12[78], stage2_12[79], stage2_12[80], stage2_12[81], stage2_12[82], stage2_12[83]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[19],stage3_14[24],stage3_13[25],stage3_12[37]}
   );
   gpc606_5 gpc3407 (
      {stage2_12[84], stage2_12[85], stage2_12[86], stage2_12[87], stage2_12[88], stage2_12[89]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[20],stage3_14[25],stage3_13[26],stage3_12[38]}
   );
   gpc606_5 gpc3408 (
      {stage2_12[90], stage2_12[91], stage2_12[92], stage2_12[93], stage2_12[94], stage2_12[95]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[21],stage3_14[26],stage3_13[27],stage3_12[39]}
   );
   gpc606_5 gpc3409 (
      {stage2_12[96], stage2_12[97], stage2_12[98], stage2_12[99], stage2_12[100], stage2_12[101]},
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage3_16[11],stage3_15[22],stage3_14[27],stage3_13[28],stage3_12[40]}
   );
   gpc606_5 gpc3410 (
      {stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69], stage2_13[70], stage2_13[71]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[12],stage3_15[23],stage3_14[28],stage3_13[29]}
   );
   gpc606_5 gpc3411 (
      {stage2_13[72], stage2_13[73], stage2_13[74], stage2_13[75], stage2_13[76], stage2_13[77]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[13],stage3_15[24],stage3_14[29],stage3_13[30]}
   );
   gpc606_5 gpc3412 (
      {stage2_13[78], stage2_13[79], stage2_13[80], stage2_13[81], stage2_13[82], stage2_13[83]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[14],stage3_15[25],stage3_14[30],stage3_13[31]}
   );
   gpc606_5 gpc3413 (
      {stage2_13[84], stage2_13[85], stage2_13[86], stage2_13[87], stage2_13[88], stage2_13[89]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[15],stage3_15[26],stage3_14[31],stage3_13[32]}
   );
   gpc615_5 gpc3414 (
      {stage2_13[90], stage2_13[91], stage2_13[92], stage2_13[93], stage2_13[94]},
      {stage2_14[72]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[16],stage3_15[27],stage3_14[32],stage3_13[33]}
   );
   gpc615_5 gpc3415 (
      {stage2_14[73], stage2_14[74], stage2_14[75], stage2_14[76], stage2_14[77]},
      {stage2_15[30]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[5],stage3_16[17],stage3_15[28],stage3_14[33]}
   );
   gpc615_5 gpc3416 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82]},
      {stage2_15[31]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[6],stage3_16[18],stage3_15[29],stage3_14[34]}
   );
   gpc615_5 gpc3417 (
      {stage2_14[83], stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87]},
      {stage2_15[32]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[7],stage3_16[19],stage3_15[30],stage3_14[35]}
   );
   gpc615_5 gpc3418 (
      {stage2_14[88], stage2_14[89], stage2_14[90], stage2_14[91], stage2_14[92]},
      {stage2_15[33]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[8],stage3_16[20],stage3_15[31],stage3_14[36]}
   );
   gpc615_5 gpc3419 (
      {stage2_14[93], stage2_14[94], stage2_14[95], stage2_14[96], stage2_14[97]},
      {stage2_15[34]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[9],stage3_16[21],stage3_15[32],stage3_14[37]}
   );
   gpc615_5 gpc3420 (
      {stage2_14[98], stage2_14[99], stage2_14[100], stage2_14[101], stage2_14[102]},
      {stage2_15[35]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[10],stage3_16[22],stage3_15[33],stage3_14[38]}
   );
   gpc615_5 gpc3421 (
      {stage2_14[103], stage2_14[104], stage2_14[105], stage2_14[106], stage2_14[107]},
      {stage2_15[36]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[11],stage3_16[23],stage3_15[34],stage3_14[39]}
   );
   gpc615_5 gpc3422 (
      {stage2_14[108], stage2_14[109], stage2_14[110], stage2_14[111], stage2_14[112]},
      {stage2_15[37]},
      {stage2_16[42], stage2_16[43], stage2_16[44], stage2_16[45], stage2_16[46], stage2_16[47]},
      {stage3_18[7],stage3_17[12],stage3_16[24],stage3_15[35],stage3_14[40]}
   );
   gpc615_5 gpc3423 (
      {stage2_14[113], stage2_14[114], stage2_14[115], stage2_14[116], stage2_14[117]},
      {stage2_15[38]},
      {stage2_16[48], stage2_16[49], stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53]},
      {stage3_18[8],stage3_17[13],stage3_16[25],stage3_15[36],stage3_14[41]}
   );
   gpc615_5 gpc3424 (
      {stage2_14[118], stage2_14[119], stage2_14[120], stage2_14[121], stage2_14[122]},
      {stage2_15[39]},
      {stage2_16[54], stage2_16[55], stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59]},
      {stage3_18[9],stage3_17[14],stage3_16[26],stage3_15[37],stage3_14[42]}
   );
   gpc615_5 gpc3425 (
      {stage2_14[123], stage2_14[124], stage2_14[125], stage2_14[126], stage2_14[127]},
      {stage2_15[40]},
      {stage2_16[60], stage2_16[61], stage2_16[62], stage2_16[63], stage2_16[64], stage2_16[65]},
      {stage3_18[10],stage3_17[15],stage3_16[27],stage3_15[38],stage3_14[43]}
   );
   gpc615_5 gpc3426 (
      {stage2_14[128], stage2_14[129], stage2_14[130], stage2_14[131], stage2_14[132]},
      {stage2_15[41]},
      {stage2_16[66], stage2_16[67], stage2_16[68], stage2_16[69], stage2_16[70], stage2_16[71]},
      {stage3_18[11],stage3_17[16],stage3_16[28],stage3_15[39],stage3_14[44]}
   );
   gpc2135_5 gpc3427 (
      {stage2_15[42], stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46]},
      {stage2_16[72], stage2_16[73], stage2_16[74]},
      {stage2_17[0]},
      {stage2_18[0], stage2_18[1]},
      {stage3_19[0],stage3_18[12],stage3_17[17],stage3_16[29],stage3_15[40]}
   );
   gpc606_5 gpc3428 (
      {stage2_15[47], stage2_15[48], stage2_15[49], stage2_15[50], stage2_15[51], stage2_15[52]},
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6]},
      {stage3_19[1],stage3_18[13],stage3_17[18],stage3_16[30],stage3_15[41]}
   );
   gpc606_5 gpc3429 (
      {stage2_15[53], stage2_15[54], stage2_15[55], stage2_15[56], stage2_15[57], stage2_15[58]},
      {stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12]},
      {stage3_19[2],stage3_18[14],stage3_17[19],stage3_16[31],stage3_15[42]}
   );
   gpc606_5 gpc3430 (
      {stage2_15[59], stage2_15[60], stage2_15[61], stage2_15[62], stage2_15[63], stage2_15[64]},
      {stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17], stage2_17[18]},
      {stage3_19[3],stage3_18[15],stage3_17[20],stage3_16[32],stage3_15[43]}
   );
   gpc606_5 gpc3431 (
      {stage2_15[65], stage2_15[66], stage2_15[67], stage2_15[68], stage2_15[69], stage2_15[70]},
      {stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23], stage2_17[24]},
      {stage3_19[4],stage3_18[16],stage3_17[21],stage3_16[33],stage3_15[44]}
   );
   gpc606_5 gpc3432 (
      {stage2_15[71], stage2_15[72], stage2_15[73], stage2_15[74], stage2_15[75], stage2_15[76]},
      {stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29], stage2_17[30]},
      {stage3_19[5],stage3_18[17],stage3_17[22],stage3_16[34],stage3_15[45]}
   );
   gpc606_5 gpc3433 (
      {stage2_15[77], stage2_15[78], stage2_15[79], stage2_15[80], stage2_15[81], stage2_15[82]},
      {stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35], stage2_17[36]},
      {stage3_19[6],stage3_18[18],stage3_17[23],stage3_16[35],stage3_15[46]}
   );
   gpc606_5 gpc3434 (
      {stage2_15[83], stage2_15[84], stage2_15[85], stage2_15[86], stage2_15[87], stage2_15[88]},
      {stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41], stage2_17[42]},
      {stage3_19[7],stage3_18[19],stage3_17[24],stage3_16[36],stage3_15[47]}
   );
   gpc606_5 gpc3435 (
      {stage2_15[89], stage2_15[90], stage2_15[91], stage2_15[92], stage2_15[93], stage2_15[94]},
      {stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47], stage2_17[48]},
      {stage3_19[8],stage3_18[20],stage3_17[25],stage3_16[37],stage3_15[48]}
   );
   gpc606_5 gpc3436 (
      {stage2_16[75], stage2_16[76], stage2_16[77], stage2_16[78], stage2_16[79], stage2_16[80]},
      {stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6], stage2_18[7]},
      {stage3_20[0],stage3_19[9],stage3_18[21],stage3_17[26],stage3_16[38]}
   );
   gpc606_5 gpc3437 (
      {stage2_17[49], stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53], stage2_17[54]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[1],stage3_19[10],stage3_18[22],stage3_17[27]}
   );
   gpc606_5 gpc3438 (
      {stage2_17[55], stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59], stage2_17[60]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[2],stage3_19[11],stage3_18[23],stage3_17[28]}
   );
   gpc606_5 gpc3439 (
      {stage2_17[61], stage2_17[62], stage2_17[63], stage2_17[64], stage2_17[65], stage2_17[66]},
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage3_21[2],stage3_20[3],stage3_19[12],stage3_18[24],stage3_17[29]}
   );
   gpc606_5 gpc3440 (
      {stage2_17[67], stage2_17[68], stage2_17[69], stage2_17[70], stage2_17[71], stage2_17[72]},
      {stage2_19[18], stage2_19[19], stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage3_21[3],stage3_20[4],stage3_19[13],stage3_18[25],stage3_17[30]}
   );
   gpc606_5 gpc3441 (
      {stage2_17[73], stage2_17[74], stage2_17[75], stage2_17[76], stage2_17[77], stage2_17[78]},
      {stage2_19[24], stage2_19[25], stage2_19[26], stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage3_21[4],stage3_20[5],stage3_19[14],stage3_18[26],stage3_17[31]}
   );
   gpc606_5 gpc3442 (
      {stage2_17[79], stage2_17[80], stage2_17[81], stage2_17[82], stage2_17[83], stage2_17[84]},
      {stage2_19[30], stage2_19[31], stage2_19[32], stage2_19[33], stage2_19[34], stage2_19[35]},
      {stage3_21[5],stage3_20[6],stage3_19[15],stage3_18[27],stage3_17[32]}
   );
   gpc606_5 gpc3443 (
      {stage2_17[85], stage2_17[86], stage2_17[87], stage2_17[88], stage2_17[89], stage2_17[90]},
      {stage2_19[36], stage2_19[37], stage2_19[38], stage2_19[39], stage2_19[40], stage2_19[41]},
      {stage3_21[6],stage3_20[7],stage3_19[16],stage3_18[28],stage3_17[33]}
   );
   gpc606_5 gpc3444 (
      {stage2_17[91], stage2_17[92], stage2_17[93], stage2_17[94], stage2_17[95], stage2_17[96]},
      {stage2_19[42], stage2_19[43], stage2_19[44], stage2_19[45], stage2_19[46], stage2_19[47]},
      {stage3_21[7],stage3_20[8],stage3_19[17],stage3_18[29],stage3_17[34]}
   );
   gpc606_5 gpc3445 (
      {stage2_17[97], stage2_17[98], stage2_17[99], stage2_17[100], stage2_17[101], stage2_17[102]},
      {stage2_19[48], stage2_19[49], stage2_19[50], stage2_19[51], stage2_19[52], stage2_19[53]},
      {stage3_21[8],stage3_20[9],stage3_19[18],stage3_18[30],stage3_17[35]}
   );
   gpc606_5 gpc3446 (
      {stage2_17[103], stage2_17[104], stage2_17[105], stage2_17[106], stage2_17[107], stage2_17[108]},
      {stage2_19[54], stage2_19[55], stage2_19[56], stage2_19[57], stage2_19[58], stage2_19[59]},
      {stage3_21[9],stage3_20[10],stage3_19[19],stage3_18[31],stage3_17[36]}
   );
   gpc1343_5 gpc3447 (
      {stage2_18[8], stage2_18[9], stage2_18[10]},
      {stage2_19[60], stage2_19[61], stage2_19[62], stage2_19[63]},
      {stage2_20[0], stage2_20[1], stage2_20[2]},
      {stage2_21[0]},
      {stage3_22[0],stage3_21[10],stage3_20[11],stage3_19[20],stage3_18[32]}
   );
   gpc1343_5 gpc3448 (
      {stage2_18[11], stage2_18[12], stage2_18[13]},
      {stage2_19[64], stage2_19[65], stage2_19[66], stage2_19[67]},
      {stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage2_21[1]},
      {stage3_22[1],stage3_21[11],stage3_20[12],stage3_19[21],stage3_18[33]}
   );
   gpc1343_5 gpc3449 (
      {stage2_18[14], stage2_18[15], stage2_18[16]},
      {stage2_19[68], stage2_19[69], stage2_19[70], stage2_19[71]},
      {stage2_20[6], stage2_20[7], stage2_20[8]},
      {stage2_21[2]},
      {stage3_22[2],stage3_21[12],stage3_20[13],stage3_19[22],stage3_18[34]}
   );
   gpc1343_5 gpc3450 (
      {stage2_18[17], stage2_18[18], stage2_18[19]},
      {stage2_19[72], stage2_19[73], stage2_19[74], stage2_19[75]},
      {stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage2_21[3]},
      {stage3_22[3],stage3_21[13],stage3_20[14],stage3_19[23],stage3_18[35]}
   );
   gpc615_5 gpc3451 (
      {stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24]},
      {stage2_19[76]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[4],stage3_21[14],stage3_20[15],stage3_19[24],stage3_18[36]}
   );
   gpc615_5 gpc3452 (
      {stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29]},
      {stage2_19[77]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[5],stage3_21[15],stage3_20[16],stage3_19[25],stage3_18[37]}
   );
   gpc615_5 gpc3453 (
      {stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34]},
      {stage2_19[78]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[6],stage3_21[16],stage3_20[17],stage3_19[26],stage3_18[38]}
   );
   gpc615_5 gpc3454 (
      {stage2_18[35], stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39]},
      {stage2_19[79]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[7],stage3_21[17],stage3_20[18],stage3_19[27],stage3_18[39]}
   );
   gpc615_5 gpc3455 (
      {stage2_18[40], stage2_18[41], stage2_18[42], stage2_18[43], stage2_18[44]},
      {stage2_19[80]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[8],stage3_21[18],stage3_20[19],stage3_19[28],stage3_18[40]}
   );
   gpc615_5 gpc3456 (
      {stage2_18[45], stage2_18[46], stage2_18[47], stage2_18[48], stage2_18[49]},
      {stage2_19[81]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[9],stage3_21[19],stage3_20[20],stage3_19[29],stage3_18[41]}
   );
   gpc615_5 gpc3457 (
      {stage2_18[50], stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54]},
      {stage2_19[82]},
      {stage2_20[48], stage2_20[49], stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53]},
      {stage3_22[10],stage3_21[20],stage3_20[21],stage3_19[30],stage3_18[42]}
   );
   gpc615_5 gpc3458 (
      {stage2_18[55], stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59]},
      {stage2_19[83]},
      {stage2_20[54], stage2_20[55], stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59]},
      {stage3_22[11],stage3_21[21],stage3_20[22],stage3_19[31],stage3_18[43]}
   );
   gpc615_5 gpc3459 (
      {stage2_18[60], stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64]},
      {stage2_19[84]},
      {stage2_20[60], stage2_20[61], stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65]},
      {stage3_22[12],stage3_21[22],stage3_20[23],stage3_19[32],stage3_18[44]}
   );
   gpc615_5 gpc3460 (
      {stage2_18[65], stage2_18[66], stage2_18[67], stage2_18[68], stage2_18[69]},
      {stage2_19[85]},
      {stage2_20[66], stage2_20[67], stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71]},
      {stage3_22[13],stage3_21[23],stage3_20[24],stage3_19[33],stage3_18[45]}
   );
   gpc615_5 gpc3461 (
      {stage2_18[70], stage2_18[71], stage2_18[72], stage2_18[73], stage2_18[74]},
      {stage2_19[86]},
      {stage2_20[72], stage2_20[73], stage2_20[74], stage2_20[75], stage2_20[76], stage2_20[77]},
      {stage3_22[14],stage3_21[24],stage3_20[25],stage3_19[34],stage3_18[46]}
   );
   gpc615_5 gpc3462 (
      {stage2_18[75], stage2_18[76], stage2_18[77], stage2_18[78], stage2_18[79]},
      {stage2_19[87]},
      {stage2_20[78], stage2_20[79], stage2_20[80], stage2_20[81], stage2_20[82], stage2_20[83]},
      {stage3_22[15],stage3_21[25],stage3_20[26],stage3_19[35],stage3_18[47]}
   );
   gpc615_5 gpc3463 (
      {stage2_19[88], stage2_19[89], stage2_19[90], stage2_19[91], stage2_19[92]},
      {stage2_20[84]},
      {stage2_21[4], stage2_21[5], stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9]},
      {stage3_23[0],stage3_22[16],stage3_21[26],stage3_20[27],stage3_19[36]}
   );
   gpc615_5 gpc3464 (
      {stage2_19[93], stage2_19[94], stage2_19[95], stage2_19[96], stage2_19[97]},
      {stage2_20[85]},
      {stage2_21[10], stage2_21[11], stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15]},
      {stage3_23[1],stage3_22[17],stage3_21[27],stage3_20[28],stage3_19[37]}
   );
   gpc606_5 gpc3465 (
      {stage2_20[86], stage2_20[87], stage2_20[88], stage2_20[89], stage2_20[90], stage2_20[91]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[2],stage3_22[18],stage3_21[28],stage3_20[29]}
   );
   gpc606_5 gpc3466 (
      {stage2_20[92], stage2_20[93], stage2_20[94], stage2_20[95], stage2_20[96], stage2_20[97]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[1],stage3_23[3],stage3_22[19],stage3_21[29],stage3_20[30]}
   );
   gpc606_5 gpc3467 (
      {stage2_20[98], stage2_20[99], stage2_20[100], stage2_20[101], stage2_20[102], stage2_20[103]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[2],stage3_23[4],stage3_22[20],stage3_21[30],stage3_20[31]}
   );
   gpc606_5 gpc3468 (
      {stage2_20[104], stage2_20[105], stage2_20[106], stage2_20[107], stage2_20[108], stage2_20[109]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage3_24[3],stage3_23[5],stage3_22[21],stage3_21[31],stage3_20[32]}
   );
   gpc606_5 gpc3469 (
      {stage2_20[110], stage2_20[111], stage2_20[112], stage2_20[113], stage2_20[114], stage2_20[115]},
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage3_24[4],stage3_23[6],stage3_22[22],stage3_21[32],stage3_20[33]}
   );
   gpc1163_5 gpc3470 (
      {stage2_21[16], stage2_21[17], stage2_21[18]},
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34], stage2_22[35]},
      {stage2_23[0]},
      {stage2_24[0]},
      {stage3_25[0],stage3_24[5],stage3_23[7],stage3_22[23],stage3_21[33]}
   );
   gpc1163_5 gpc3471 (
      {stage2_21[19], stage2_21[20], stage2_21[21]},
      {stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39], stage2_22[40], stage2_22[41]},
      {stage2_23[1]},
      {stage2_24[1]},
      {stage3_25[1],stage3_24[6],stage3_23[8],stage3_22[24],stage3_21[34]}
   );
   gpc1163_5 gpc3472 (
      {stage2_21[22], stage2_21[23], stage2_21[24]},
      {stage2_22[42], stage2_22[43], stage2_22[44], stage2_22[45], stage2_22[46], stage2_22[47]},
      {stage2_23[2]},
      {stage2_24[2]},
      {stage3_25[2],stage3_24[7],stage3_23[9],stage3_22[25],stage3_21[35]}
   );
   gpc1163_5 gpc3473 (
      {stage2_21[25], stage2_21[26], stage2_21[27]},
      {stage2_22[48], stage2_22[49], stage2_22[50], stage2_22[51], stage2_22[52], stage2_22[53]},
      {stage2_23[3]},
      {stage2_24[3]},
      {stage3_25[3],stage3_24[8],stage3_23[10],stage3_22[26],stage3_21[36]}
   );
   gpc1163_5 gpc3474 (
      {stage2_21[28], stage2_21[29], stage2_21[30]},
      {stage2_22[54], stage2_22[55], stage2_22[56], stage2_22[57], stage2_22[58], stage2_22[59]},
      {stage2_23[4]},
      {stage2_24[4]},
      {stage3_25[4],stage3_24[9],stage3_23[11],stage3_22[27],stage3_21[37]}
   );
   gpc1163_5 gpc3475 (
      {stage2_21[31], stage2_21[32], stage2_21[33]},
      {stage2_22[60], stage2_22[61], stage2_22[62], stage2_22[63], stage2_22[64], stage2_22[65]},
      {stage2_23[5]},
      {stage2_24[5]},
      {stage3_25[5],stage3_24[10],stage3_23[12],stage3_22[28],stage3_21[38]}
   );
   gpc606_5 gpc3476 (
      {stage2_21[34], stage2_21[35], stage2_21[36], stage2_21[37], stage2_21[38], stage2_21[39]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[6],stage3_24[11],stage3_23[13],stage3_22[29],stage3_21[39]}
   );
   gpc606_5 gpc3477 (
      {stage2_21[40], stage2_21[41], stage2_21[42], stage2_21[43], stage2_21[44], stage2_21[45]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[7],stage3_24[12],stage3_23[14],stage3_22[30],stage3_21[40]}
   );
   gpc606_5 gpc3478 (
      {stage2_21[46], stage2_21[47], stage2_21[48], stage2_21[49], stage2_21[50], stage2_21[51]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[8],stage3_24[13],stage3_23[15],stage3_22[31],stage3_21[41]}
   );
   gpc606_5 gpc3479 (
      {stage2_21[52], stage2_21[53], stage2_21[54], stage2_21[55], stage2_21[56], stage2_21[57]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[9],stage3_24[14],stage3_23[16],stage3_22[32],stage3_21[42]}
   );
   gpc606_5 gpc3480 (
      {stage2_21[58], stage2_21[59], stage2_21[60], stage2_21[61], stage2_21[62], stage2_21[63]},
      {stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35]},
      {stage3_25[10],stage3_24[15],stage3_23[17],stage3_22[33],stage3_21[43]}
   );
   gpc615_5 gpc3481 (
      {stage2_23[36], stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40]},
      {stage2_24[6]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[0],stage3_25[11],stage3_24[16],stage3_23[18]}
   );
   gpc615_5 gpc3482 (
      {stage2_23[41], stage2_23[42], stage2_23[43], stage2_23[44], stage2_23[45]},
      {stage2_24[7]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[1],stage3_25[12],stage3_24[17],stage3_23[19]}
   );
   gpc615_5 gpc3483 (
      {stage2_23[46], stage2_23[47], stage2_23[48], stage2_23[49], stage2_23[50]},
      {stage2_24[8]},
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage3_27[2],stage3_26[2],stage3_25[13],stage3_24[18],stage3_23[20]}
   );
   gpc615_5 gpc3484 (
      {stage2_23[51], stage2_23[52], stage2_23[53], stage2_23[54], stage2_23[55]},
      {stage2_24[9]},
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage3_27[3],stage3_26[3],stage3_25[14],stage3_24[19],stage3_23[21]}
   );
   gpc615_5 gpc3485 (
      {stage2_23[56], stage2_23[57], stage2_23[58], stage2_23[59], stage2_23[60]},
      {stage2_24[10]},
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage3_27[4],stage3_26[4],stage3_25[15],stage3_24[20],stage3_23[22]}
   );
   gpc615_5 gpc3486 (
      {stage2_23[61], stage2_23[62], stage2_23[63], stage2_23[64], stage2_23[65]},
      {stage2_24[11]},
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage3_27[5],stage3_26[5],stage3_25[16],stage3_24[21],stage3_23[23]}
   );
   gpc615_5 gpc3487 (
      {stage2_23[66], stage2_23[67], stage2_23[68], stage2_23[69], stage2_23[70]},
      {stage2_24[12]},
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage3_27[6],stage3_26[6],stage3_25[17],stage3_24[22],stage3_23[24]}
   );
   gpc615_5 gpc3488 (
      {stage2_23[71], stage2_23[72], stage2_23[73], stage2_23[74], stage2_23[75]},
      {stage2_24[13]},
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46], stage2_25[47]},
      {stage3_27[7],stage3_26[7],stage3_25[18],stage3_24[23],stage3_23[25]}
   );
   gpc615_5 gpc3489 (
      {stage2_23[76], stage2_23[77], stage2_23[78], stage2_23[79], stage2_23[80]},
      {stage2_24[14]},
      {stage2_25[48], stage2_25[49], stage2_25[50], stage2_25[51], stage2_25[52], stage2_25[53]},
      {stage3_27[8],stage3_26[8],stage3_25[19],stage3_24[24],stage3_23[26]}
   );
   gpc615_5 gpc3490 (
      {stage2_23[81], stage2_23[82], stage2_23[83], stage2_23[84], stage2_23[85]},
      {stage2_24[15]},
      {stage2_25[54], stage2_25[55], stage2_25[56], stage2_25[57], stage2_25[58], stage2_25[59]},
      {stage3_27[9],stage3_26[9],stage3_25[20],stage3_24[25],stage3_23[27]}
   );
   gpc615_5 gpc3491 (
      {stage2_23[86], stage2_23[87], stage2_23[88], stage2_23[89], stage2_23[90]},
      {stage2_24[16]},
      {stage2_25[60], stage2_25[61], stage2_25[62], stage2_25[63], stage2_25[64], stage2_25[65]},
      {stage3_27[10],stage3_26[10],stage3_25[21],stage3_24[26],stage3_23[28]}
   );
   gpc606_5 gpc3492 (
      {stage2_24[17], stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[11],stage3_26[11],stage3_25[22],stage3_24[27]}
   );
   gpc606_5 gpc3493 (
      {stage2_24[23], stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[12],stage3_26[12],stage3_25[23],stage3_24[28]}
   );
   gpc606_5 gpc3494 (
      {stage2_24[29], stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[13],stage3_26[13],stage3_25[24],stage3_24[29]}
   );
   gpc606_5 gpc3495 (
      {stage2_24[35], stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40]},
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23]},
      {stage3_28[3],stage3_27[14],stage3_26[14],stage3_25[25],stage3_24[30]}
   );
   gpc606_5 gpc3496 (
      {stage2_24[41], stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46]},
      {stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29]},
      {stage3_28[4],stage3_27[15],stage3_26[15],stage3_25[26],stage3_24[31]}
   );
   gpc606_5 gpc3497 (
      {stage2_24[47], stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52]},
      {stage2_26[30], stage2_26[31], stage2_26[32], stage2_26[33], stage2_26[34], stage2_26[35]},
      {stage3_28[5],stage3_27[16],stage3_26[16],stage3_25[27],stage3_24[32]}
   );
   gpc606_5 gpc3498 (
      {stage2_24[53], stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58]},
      {stage2_26[36], stage2_26[37], stage2_26[38], stage2_26[39], stage2_26[40], stage2_26[41]},
      {stage3_28[6],stage3_27[17],stage3_26[17],stage3_25[28],stage3_24[33]}
   );
   gpc606_5 gpc3499 (
      {stage2_24[59], stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64]},
      {stage2_26[42], stage2_26[43], stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47]},
      {stage3_28[7],stage3_27[18],stage3_26[18],stage3_25[29],stage3_24[34]}
   );
   gpc606_5 gpc3500 (
      {stage2_24[65], stage2_24[66], stage2_24[67], stage2_24[68], stage2_24[69], stage2_24[70]},
      {stage2_26[48], stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52], stage2_26[53]},
      {stage3_28[8],stage3_27[19],stage3_26[19],stage3_25[30],stage3_24[35]}
   );
   gpc606_5 gpc3501 (
      {stage2_24[71], stage2_24[72], stage2_24[73], stage2_24[74], stage2_24[75], stage2_24[76]},
      {stage2_26[54], stage2_26[55], stage2_26[56], stage2_26[57], stage2_26[58], stage2_26[59]},
      {stage3_28[9],stage3_27[20],stage3_26[20],stage3_25[31],stage3_24[36]}
   );
   gpc606_5 gpc3502 (
      {stage2_24[77], stage2_24[78], stage2_24[79], stage2_24[80], stage2_24[81], stage2_24[82]},
      {stage2_26[60], stage2_26[61], stage2_26[62], stage2_26[63], stage2_26[64], stage2_26[65]},
      {stage3_28[10],stage3_27[21],stage3_26[21],stage3_25[32],stage3_24[37]}
   );
   gpc606_5 gpc3503 (
      {stage2_24[83], stage2_24[84], stage2_24[85], stage2_24[86], stage2_24[87], stage2_24[88]},
      {stage2_26[66], stage2_26[67], stage2_26[68], stage2_26[69], stage2_26[70], stage2_26[71]},
      {stage3_28[11],stage3_27[22],stage3_26[22],stage3_25[33],stage3_24[38]}
   );
   gpc606_5 gpc3504 (
      {stage2_24[89], stage2_24[90], stage2_24[91], stage2_24[92], stage2_24[93], stage2_24[94]},
      {stage2_26[72], stage2_26[73], stage2_26[74], stage2_26[75], stage2_26[76], stage2_26[77]},
      {stage3_28[12],stage3_27[23],stage3_26[23],stage3_25[34],stage3_24[39]}
   );
   gpc606_5 gpc3505 (
      {stage2_24[95], stage2_24[96], stage2_24[97], stage2_24[98], stage2_24[99], 1'b0},
      {stage2_26[78], stage2_26[79], stage2_26[80], stage2_26[81], stage2_26[82], stage2_26[83]},
      {stage3_28[13],stage3_27[24],stage3_26[24],stage3_25[35],stage3_24[40]}
   );
   gpc606_5 gpc3506 (
      {stage2_25[66], stage2_25[67], stage2_25[68], stage2_25[69], stage2_25[70], stage2_25[71]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[14],stage3_27[25],stage3_26[25],stage3_25[36]}
   );
   gpc606_5 gpc3507 (
      {stage2_25[72], stage2_25[73], stage2_25[74], stage2_25[75], stage2_25[76], stage2_25[77]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[15],stage3_27[26],stage3_26[26],stage3_25[37]}
   );
   gpc606_5 gpc3508 (
      {stage2_25[78], stage2_25[79], stage2_25[80], stage2_25[81], stage2_25[82], stage2_25[83]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[16],stage3_27[27],stage3_26[27],stage3_25[38]}
   );
   gpc606_5 gpc3509 (
      {stage2_25[84], stage2_25[85], stage2_25[86], stage2_25[87], 1'b0, 1'b0},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[17],stage3_27[28],stage3_26[28],stage3_25[39]}
   );
   gpc615_5 gpc3510 (
      {stage2_26[84], stage2_26[85], stage2_26[86], stage2_26[87], stage2_26[88]},
      {stage2_27[24]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[4],stage3_28[18],stage3_27[29],stage3_26[29]}
   );
   gpc615_5 gpc3511 (
      {stage2_26[89], stage2_26[90], stage2_26[91], stage2_26[92], stage2_26[93]},
      {stage2_27[25]},
      {stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11]},
      {stage3_30[1],stage3_29[5],stage3_28[19],stage3_27[30],stage3_26[30]}
   );
   gpc615_5 gpc3512 (
      {stage2_26[94], stage2_26[95], stage2_26[96], stage2_26[97], stage2_26[98]},
      {stage2_27[26]},
      {stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17]},
      {stage3_30[2],stage3_29[6],stage3_28[20],stage3_27[31],stage3_26[31]}
   );
   gpc606_5 gpc3513 (
      {stage2_27[27], stage2_27[28], stage2_27[29], stage2_27[30], stage2_27[31], stage2_27[32]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[3],stage3_29[7],stage3_28[21],stage3_27[32]}
   );
   gpc606_5 gpc3514 (
      {stage2_27[33], stage2_27[34], stage2_27[35], stage2_27[36], stage2_27[37], stage2_27[38]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[4],stage3_29[8],stage3_28[22],stage3_27[33]}
   );
   gpc606_5 gpc3515 (
      {stage2_27[39], stage2_27[40], stage2_27[41], stage2_27[42], stage2_27[43], stage2_27[44]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[5],stage3_29[9],stage3_28[23],stage3_27[34]}
   );
   gpc615_5 gpc3516 (
      {stage2_27[45], stage2_27[46], stage2_27[47], stage2_27[48], stage2_27[49]},
      {stage2_28[18]},
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage3_31[3],stage3_30[6],stage3_29[10],stage3_28[24],stage3_27[35]}
   );
   gpc615_5 gpc3517 (
      {stage2_27[50], stage2_27[51], stage2_27[52], stage2_27[53], stage2_27[54]},
      {stage2_28[19]},
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage3_31[4],stage3_30[7],stage3_29[11],stage3_28[25],stage3_27[36]}
   );
   gpc615_5 gpc3518 (
      {stage2_27[55], stage2_27[56], stage2_27[57], stage2_27[58], stage2_27[59]},
      {stage2_28[20]},
      {stage2_29[30], stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage3_31[5],stage3_30[8],stage3_29[12],stage3_28[26],stage3_27[37]}
   );
   gpc615_5 gpc3519 (
      {stage2_27[60], stage2_27[61], stage2_27[62], stage2_27[63], stage2_27[64]},
      {stage2_28[21]},
      {stage2_29[36], stage2_29[37], stage2_29[38], stage2_29[39], stage2_29[40], stage2_29[41]},
      {stage3_31[6],stage3_30[9],stage3_29[13],stage3_28[27],stage3_27[38]}
   );
   gpc615_5 gpc3520 (
      {stage2_27[65], stage2_27[66], stage2_27[67], stage2_27[68], stage2_27[69]},
      {stage2_28[22]},
      {stage2_29[42], stage2_29[43], stage2_29[44], stage2_29[45], stage2_29[46], stage2_29[47]},
      {stage3_31[7],stage3_30[10],stage3_29[14],stage3_28[28],stage3_27[39]}
   );
   gpc606_5 gpc3521 (
      {stage2_28[23], stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[8],stage3_30[11],stage3_29[15],stage3_28[29]}
   );
   gpc606_5 gpc3522 (
      {stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[9],stage3_30[12],stage3_29[16],stage3_28[30]}
   );
   gpc606_5 gpc3523 (
      {stage2_28[35], stage2_28[36], stage2_28[37], stage2_28[38], stage2_28[39], stage2_28[40]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[10],stage3_30[13],stage3_29[17],stage3_28[31]}
   );
   gpc606_5 gpc3524 (
      {stage2_28[41], stage2_28[42], stage2_28[43], stage2_28[44], stage2_28[45], stage2_28[46]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[11],stage3_30[14],stage3_29[18],stage3_28[32]}
   );
   gpc606_5 gpc3525 (
      {stage2_28[47], stage2_28[48], stage2_28[49], stage2_28[50], stage2_28[51], stage2_28[52]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[12],stage3_30[15],stage3_29[19],stage3_28[33]}
   );
   gpc606_5 gpc3526 (
      {stage2_28[53], stage2_28[54], stage2_28[55], stage2_28[56], stage2_28[57], stage2_28[58]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage3_32[5],stage3_31[13],stage3_30[16],stage3_29[20],stage3_28[34]}
   );
   gpc615_5 gpc3527 (
      {stage2_28[59], stage2_28[60], stage2_28[61], stage2_28[62], stage2_28[63]},
      {stage2_29[48]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage3_32[6],stage3_31[14],stage3_30[17],stage3_29[21],stage3_28[35]}
   );
   gpc615_5 gpc3528 (
      {stage2_28[64], stage2_28[65], stage2_28[66], stage2_28[67], stage2_28[68]},
      {stage2_29[49]},
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage3_32[7],stage3_31[15],stage3_30[18],stage3_29[22],stage3_28[36]}
   );
   gpc1163_5 gpc3529 (
      {stage2_29[50], stage2_29[51], stage2_29[52]},
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], stage2_30[52], stage2_30[53]},
      {stage2_31[0]},
      {stage2_32[0]},
      {stage3_33[0],stage3_32[8],stage3_31[16],stage3_30[19],stage3_29[23]}
   );
   gpc1163_5 gpc3530 (
      {stage2_29[53], stage2_29[54], stage2_29[55]},
      {stage2_30[54], stage2_30[55], stage2_30[56], stage2_30[57], stage2_30[58], stage2_30[59]},
      {stage2_31[1]},
      {stage2_32[1]},
      {stage3_33[1],stage3_32[9],stage3_31[17],stage3_30[20],stage3_29[24]}
   );
   gpc1163_5 gpc3531 (
      {stage2_29[56], stage2_29[57], stage2_29[58]},
      {stage2_30[60], stage2_30[61], stage2_30[62], stage2_30[63], stage2_30[64], stage2_30[65]},
      {stage2_31[2]},
      {stage2_32[2]},
      {stage3_33[2],stage3_32[10],stage3_31[18],stage3_30[21],stage3_29[25]}
   );
   gpc1163_5 gpc3532 (
      {stage2_29[59], stage2_29[60], stage2_29[61]},
      {stage2_30[66], stage2_30[67], stage2_30[68], stage2_30[69], stage2_30[70], stage2_30[71]},
      {stage2_31[3]},
      {stage2_32[3]},
      {stage3_33[3],stage3_32[11],stage3_31[19],stage3_30[22],stage3_29[26]}
   );
   gpc1163_5 gpc3533 (
      {stage2_29[62], stage2_29[63], stage2_29[64]},
      {stage2_30[72], stage2_30[73], stage2_30[74], stage2_30[75], stage2_30[76], stage2_30[77]},
      {stage2_31[4]},
      {stage2_32[4]},
      {stage3_33[4],stage3_32[12],stage3_31[20],stage3_30[23],stage3_29[27]}
   );
   gpc606_5 gpc3534 (
      {stage2_29[65], stage2_29[66], stage2_29[67], stage2_29[68], stage2_29[69], stage2_29[70]},
      {stage2_31[5], stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10]},
      {stage3_33[5],stage3_32[13],stage3_31[21],stage3_30[24],stage3_29[28]}
   );
   gpc606_5 gpc3535 (
      {stage2_29[71], stage2_29[72], stage2_29[73], stage2_29[74], stage2_29[75], stage2_29[76]},
      {stage2_31[11], stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16]},
      {stage3_33[6],stage3_32[14],stage3_31[22],stage3_30[25],stage3_29[29]}
   );
   gpc606_5 gpc3536 (
      {stage2_29[77], stage2_29[78], stage2_29[79], stage2_29[80], stage2_29[81], stage2_29[82]},
      {stage2_31[17], stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22]},
      {stage3_33[7],stage3_32[15],stage3_31[23],stage3_30[26],stage3_29[30]}
   );
   gpc606_5 gpc3537 (
      {stage2_29[83], stage2_29[84], stage2_29[85], stage2_29[86], stage2_29[87], stage2_29[88]},
      {stage2_31[23], stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28]},
      {stage3_33[8],stage3_32[16],stage3_31[24],stage3_30[27],stage3_29[31]}
   );
   gpc606_5 gpc3538 (
      {stage2_29[89], stage2_29[90], stage2_29[91], stage2_29[92], stage2_29[93], stage2_29[94]},
      {stage2_31[29], stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], stage2_31[34]},
      {stage3_33[9],stage3_32[17],stage3_31[25],stage3_30[28],stage3_29[32]}
   );
   gpc606_5 gpc3539 (
      {stage2_29[95], stage2_29[96], stage2_29[97], stage2_29[98], stage2_29[99], stage2_29[100]},
      {stage2_31[35], stage2_31[36], stage2_31[37], stage2_31[38], stage2_31[39], stage2_31[40]},
      {stage3_33[10],stage3_32[18],stage3_31[26],stage3_30[29],stage3_29[33]}
   );
   gpc606_5 gpc3540 (
      {stage2_29[101], stage2_29[102], stage2_29[103], stage2_29[104], stage2_29[105], stage2_29[106]},
      {stage2_31[41], stage2_31[42], stage2_31[43], stage2_31[44], stage2_31[45], stage2_31[46]},
      {stage3_33[11],stage3_32[19],stage3_31[27],stage3_30[30],stage3_29[34]}
   );
   gpc606_5 gpc3541 (
      {stage2_29[107], stage2_29[108], stage2_29[109], stage2_29[110], stage2_29[111], stage2_29[112]},
      {stage2_31[47], stage2_31[48], stage2_31[49], stage2_31[50], stage2_31[51], stage2_31[52]},
      {stage3_33[12],stage3_32[20],stage3_31[28],stage3_30[31],stage3_29[35]}
   );
   gpc606_5 gpc3542 (
      {stage2_29[113], stage2_29[114], stage2_29[115], stage2_29[116], stage2_29[117], stage2_29[118]},
      {stage2_31[53], stage2_31[54], stage2_31[55], stage2_31[56], stage2_31[57], stage2_31[58]},
      {stage3_33[13],stage3_32[21],stage3_31[29],stage3_30[32],stage3_29[36]}
   );
   gpc606_5 gpc3543 (
      {stage2_30[78], stage2_30[79], stage2_30[80], stage2_30[81], stage2_30[82], stage2_30[83]},
      {stage2_32[5], stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10]},
      {stage3_34[0],stage3_33[14],stage3_32[22],stage3_31[30],stage3_30[33]}
   );
   gpc606_5 gpc3544 (
      {stage2_30[84], stage2_30[85], stage2_30[86], stage2_30[87], stage2_30[88], stage2_30[89]},
      {stage2_32[11], stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16]},
      {stage3_34[1],stage3_33[15],stage3_32[23],stage3_31[31],stage3_30[34]}
   );
   gpc606_5 gpc3545 (
      {stage2_30[90], stage2_30[91], stage2_30[92], stage2_30[93], stage2_30[94], stage2_30[95]},
      {stage2_32[17], stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22]},
      {stage3_34[2],stage3_33[16],stage3_32[24],stage3_31[32],stage3_30[35]}
   );
   gpc606_5 gpc3546 (
      {stage2_30[96], stage2_30[97], stage2_30[98], stage2_30[99], stage2_30[100], stage2_30[101]},
      {stage2_32[23], stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28]},
      {stage3_34[3],stage3_33[17],stage3_32[25],stage3_31[33],stage3_30[36]}
   );
   gpc606_5 gpc3547 (
      {stage2_30[102], stage2_30[103], stage2_30[104], stage2_30[105], stage2_30[106], stage2_30[107]},
      {stage2_32[29], stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34]},
      {stage3_34[4],stage3_33[18],stage3_32[26],stage3_31[34],stage3_30[37]}
   );
   gpc606_5 gpc3548 (
      {stage2_31[59], stage2_31[60], stage2_31[61], stage2_31[62], stage2_31[63], stage2_31[64]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[5],stage3_33[19],stage3_32[27],stage3_31[35]}
   );
   gpc606_5 gpc3549 (
      {stage2_31[65], stage2_31[66], stage2_31[67], stage2_31[68], stage2_31[69], stage2_31[70]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[6],stage3_33[20],stage3_32[28],stage3_31[36]}
   );
   gpc606_5 gpc3550 (
      {stage2_31[71], stage2_31[72], stage2_31[73], stage2_31[74], stage2_31[75], stage2_31[76]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[7],stage3_33[21],stage3_32[29],stage3_31[37]}
   );
   gpc606_5 gpc3551 (
      {stage2_31[77], stage2_31[78], stage2_31[79], stage2_31[80], stage2_31[81], stage2_31[82]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[8],stage3_33[22],stage3_32[30],stage3_31[38]}
   );
   gpc606_5 gpc3552 (
      {stage2_32[35], stage2_32[36], stage2_32[37], stage2_32[38], stage2_32[39], stage2_32[40]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[4],stage3_34[9],stage3_33[23],stage3_32[31]}
   );
   gpc606_5 gpc3553 (
      {stage2_32[41], stage2_32[42], stage2_32[43], stage2_32[44], stage2_32[45], stage2_32[46]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[5],stage3_34[10],stage3_33[24],stage3_32[32]}
   );
   gpc606_5 gpc3554 (
      {stage2_32[47], stage2_32[48], stage2_32[49], stage2_32[50], stage2_32[51], stage2_32[52]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17]},
      {stage3_36[2],stage3_35[6],stage3_34[11],stage3_33[25],stage3_32[33]}
   );
   gpc606_5 gpc3555 (
      {stage2_32[53], stage2_32[54], stage2_32[55], stage2_32[56], stage2_32[57], stage2_32[58]},
      {stage2_34[18], stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23]},
      {stage3_36[3],stage3_35[7],stage3_34[12],stage3_33[26],stage3_32[34]}
   );
   gpc606_5 gpc3556 (
      {stage2_32[59], stage2_32[60], stage2_32[61], stage2_32[62], stage2_32[63], stage2_32[64]},
      {stage2_34[24], stage2_34[25], stage2_34[26], stage2_34[27], stage2_34[28], stage2_34[29]},
      {stage3_36[4],stage3_35[8],stage3_34[13],stage3_33[27],stage3_32[35]}
   );
   gpc606_5 gpc3557 (
      {stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[5],stage3_35[9],stage3_34[14],stage3_33[28]}
   );
   gpc606_5 gpc3558 (
      {stage2_33[30], stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35]},
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage3_37[1],stage3_36[6],stage3_35[10],stage3_34[15],stage3_33[29]}
   );
   gpc1_1 gpc3559 (
      {stage2_0[21]},
      {stage3_0[7]}
   );
   gpc1_1 gpc3560 (
      {stage2_2[43]},
      {stage3_2[24]}
   );
   gpc1_1 gpc3561 (
      {stage2_2[44]},
      {stage3_2[25]}
   );
   gpc1_1 gpc3562 (
      {stage2_2[45]},
      {stage3_2[26]}
   );
   gpc1_1 gpc3563 (
      {stage2_2[46]},
      {stage3_2[27]}
   );
   gpc1_1 gpc3564 (
      {stage2_2[47]},
      {stage3_2[28]}
   );
   gpc1_1 gpc3565 (
      {stage2_2[48]},
      {stage3_2[29]}
   );
   gpc1_1 gpc3566 (
      {stage2_2[49]},
      {stage3_2[30]}
   );
   gpc1_1 gpc3567 (
      {stage2_2[50]},
      {stage3_2[31]}
   );
   gpc1_1 gpc3568 (
      {stage2_4[82]},
      {stage3_4[35]}
   );
   gpc1_1 gpc3569 (
      {stage2_4[83]},
      {stage3_4[36]}
   );
   gpc1_1 gpc3570 (
      {stage2_4[84]},
      {stage3_4[37]}
   );
   gpc1_1 gpc3571 (
      {stage2_4[85]},
      {stage3_4[38]}
   );
   gpc1_1 gpc3572 (
      {stage2_4[86]},
      {stage3_4[39]}
   );
   gpc1_1 gpc3573 (
      {stage2_4[87]},
      {stage3_4[40]}
   );
   gpc1_1 gpc3574 (
      {stage2_4[88]},
      {stage3_4[41]}
   );
   gpc1_1 gpc3575 (
      {stage2_4[89]},
      {stage3_4[42]}
   );
   gpc1_1 gpc3576 (
      {stage2_4[90]},
      {stage3_4[43]}
   );
   gpc1_1 gpc3577 (
      {stage2_5[71]},
      {stage3_5[36]}
   );
   gpc1_1 gpc3578 (
      {stage2_5[72]},
      {stage3_5[37]}
   );
   gpc1_1 gpc3579 (
      {stage2_5[73]},
      {stage3_5[38]}
   );
   gpc1_1 gpc3580 (
      {stage2_5[74]},
      {stage3_5[39]}
   );
   gpc1_1 gpc3581 (
      {stage2_5[75]},
      {stage3_5[40]}
   );
   gpc1_1 gpc3582 (
      {stage2_5[76]},
      {stage3_5[41]}
   );
   gpc1_1 gpc3583 (
      {stage2_5[77]},
      {stage3_5[42]}
   );
   gpc1_1 gpc3584 (
      {stage2_5[78]},
      {stage3_5[43]}
   );
   gpc1_1 gpc3585 (
      {stage2_5[79]},
      {stage3_5[44]}
   );
   gpc1_1 gpc3586 (
      {stage2_5[80]},
      {stage3_5[45]}
   );
   gpc1_1 gpc3587 (
      {stage2_5[81]},
      {stage3_5[46]}
   );
   gpc1_1 gpc3588 (
      {stage2_5[82]},
      {stage3_5[47]}
   );
   gpc1_1 gpc3589 (
      {stage2_5[83]},
      {stage3_5[48]}
   );
   gpc1_1 gpc3590 (
      {stage2_6[83]},
      {stage3_6[32]}
   );
   gpc1_1 gpc3591 (
      {stage2_6[84]},
      {stage3_6[33]}
   );
   gpc1_1 gpc3592 (
      {stage2_6[85]},
      {stage3_6[34]}
   );
   gpc1_1 gpc3593 (
      {stage2_6[86]},
      {stage3_6[35]}
   );
   gpc1_1 gpc3594 (
      {stage2_6[87]},
      {stage3_6[36]}
   );
   gpc1_1 gpc3595 (
      {stage2_6[88]},
      {stage3_6[37]}
   );
   gpc1_1 gpc3596 (
      {stage2_6[89]},
      {stage3_6[38]}
   );
   gpc1_1 gpc3597 (
      {stage2_6[90]},
      {stage3_6[39]}
   );
   gpc1_1 gpc3598 (
      {stage2_6[91]},
      {stage3_6[40]}
   );
   gpc1_1 gpc3599 (
      {stage2_6[92]},
      {stage3_6[41]}
   );
   gpc1_1 gpc3600 (
      {stage2_6[93]},
      {stage3_6[42]}
   );
   gpc1_1 gpc3601 (
      {stage2_7[70]},
      {stage3_7[29]}
   );
   gpc1_1 gpc3602 (
      {stage2_7[71]},
      {stage3_7[30]}
   );
   gpc1_1 gpc3603 (
      {stage2_7[72]},
      {stage3_7[31]}
   );
   gpc1_1 gpc3604 (
      {stage2_7[73]},
      {stage3_7[32]}
   );
   gpc1_1 gpc3605 (
      {stage2_7[74]},
      {stage3_7[33]}
   );
   gpc1_1 gpc3606 (
      {stage2_7[75]},
      {stage3_7[34]}
   );
   gpc1_1 gpc3607 (
      {stage2_7[76]},
      {stage3_7[35]}
   );
   gpc1_1 gpc3608 (
      {stage2_7[77]},
      {stage3_7[36]}
   );
   gpc1_1 gpc3609 (
      {stage2_7[78]},
      {stage3_7[37]}
   );
   gpc1_1 gpc3610 (
      {stage2_7[79]},
      {stage3_7[38]}
   );
   gpc1_1 gpc3611 (
      {stage2_7[80]},
      {stage3_7[39]}
   );
   gpc1_1 gpc3612 (
      {stage2_7[81]},
      {stage3_7[40]}
   );
   gpc1_1 gpc3613 (
      {stage2_7[82]},
      {stage3_7[41]}
   );
   gpc1_1 gpc3614 (
      {stage2_7[83]},
      {stage3_7[42]}
   );
   gpc1_1 gpc3615 (
      {stage2_7[84]},
      {stage3_7[43]}
   );
   gpc1_1 gpc3616 (
      {stage2_7[85]},
      {stage3_7[44]}
   );
   gpc1_1 gpc3617 (
      {stage2_7[86]},
      {stage3_7[45]}
   );
   gpc1_1 gpc3618 (
      {stage2_7[87]},
      {stage3_7[46]}
   );
   gpc1_1 gpc3619 (
      {stage2_7[88]},
      {stage3_7[47]}
   );
   gpc1_1 gpc3620 (
      {stage2_7[89]},
      {stage3_7[48]}
   );
   gpc1_1 gpc3621 (
      {stage2_7[90]},
      {stage3_7[49]}
   );
   gpc1_1 gpc3622 (
      {stage2_7[91]},
      {stage3_7[50]}
   );
   gpc1_1 gpc3623 (
      {stage2_7[92]},
      {stage3_7[51]}
   );
   gpc1_1 gpc3624 (
      {stage2_7[93]},
      {stage3_7[52]}
   );
   gpc1_1 gpc3625 (
      {stage2_7[94]},
      {stage3_7[53]}
   );
   gpc1_1 gpc3626 (
      {stage2_7[95]},
      {stage3_7[54]}
   );
   gpc1_1 gpc3627 (
      {stage2_7[96]},
      {stage3_7[55]}
   );
   gpc1_1 gpc3628 (
      {stage2_7[97]},
      {stage3_7[56]}
   );
   gpc1_1 gpc3629 (
      {stage2_7[98]},
      {stage3_7[57]}
   );
   gpc1_1 gpc3630 (
      {stage2_7[99]},
      {stage3_7[58]}
   );
   gpc1_1 gpc3631 (
      {stage2_7[100]},
      {stage3_7[59]}
   );
   gpc1_1 gpc3632 (
      {stage2_7[101]},
      {stage3_7[60]}
   );
   gpc1_1 gpc3633 (
      {stage2_7[102]},
      {stage3_7[61]}
   );
   gpc1_1 gpc3634 (
      {stage2_7[103]},
      {stage3_7[62]}
   );
   gpc1_1 gpc3635 (
      {stage2_7[104]},
      {stage3_7[63]}
   );
   gpc1_1 gpc3636 (
      {stage2_7[105]},
      {stage3_7[64]}
   );
   gpc1_1 gpc3637 (
      {stage2_7[106]},
      {stage3_7[65]}
   );
   gpc1_1 gpc3638 (
      {stage2_7[107]},
      {stage3_7[66]}
   );
   gpc1_1 gpc3639 (
      {stage2_7[108]},
      {stage3_7[67]}
   );
   gpc1_1 gpc3640 (
      {stage2_7[109]},
      {stage3_7[68]}
   );
   gpc1_1 gpc3641 (
      {stage2_9[36]},
      {stage3_9[31]}
   );
   gpc1_1 gpc3642 (
      {stage2_9[37]},
      {stage3_9[32]}
   );
   gpc1_1 gpc3643 (
      {stage2_9[38]},
      {stage3_9[33]}
   );
   gpc1_1 gpc3644 (
      {stage2_9[39]},
      {stage3_9[34]}
   );
   gpc1_1 gpc3645 (
      {stage2_9[40]},
      {stage3_9[35]}
   );
   gpc1_1 gpc3646 (
      {stage2_9[41]},
      {stage3_9[36]}
   );
   gpc1_1 gpc3647 (
      {stage2_9[42]},
      {stage3_9[37]}
   );
   gpc1_1 gpc3648 (
      {stage2_9[43]},
      {stage3_9[38]}
   );
   gpc1_1 gpc3649 (
      {stage2_9[44]},
      {stage3_9[39]}
   );
   gpc1_1 gpc3650 (
      {stage2_9[45]},
      {stage3_9[40]}
   );
   gpc1_1 gpc3651 (
      {stage2_9[46]},
      {stage3_9[41]}
   );
   gpc1_1 gpc3652 (
      {stage2_9[47]},
      {stage3_9[42]}
   );
   gpc1_1 gpc3653 (
      {stage2_9[48]},
      {stage3_9[43]}
   );
   gpc1_1 gpc3654 (
      {stage2_9[49]},
      {stage3_9[44]}
   );
   gpc1_1 gpc3655 (
      {stage2_9[50]},
      {stage3_9[45]}
   );
   gpc1_1 gpc3656 (
      {stage2_9[51]},
      {stage3_9[46]}
   );
   gpc1_1 gpc3657 (
      {stage2_9[52]},
      {stage3_9[47]}
   );
   gpc1_1 gpc3658 (
      {stage2_9[53]},
      {stage3_9[48]}
   );
   gpc1_1 gpc3659 (
      {stage2_9[54]},
      {stage3_9[49]}
   );
   gpc1_1 gpc3660 (
      {stage2_9[55]},
      {stage3_9[50]}
   );
   gpc1_1 gpc3661 (
      {stage2_9[56]},
      {stage3_9[51]}
   );
   gpc1_1 gpc3662 (
      {stage2_9[57]},
      {stage3_9[52]}
   );
   gpc1_1 gpc3663 (
      {stage2_9[58]},
      {stage3_9[53]}
   );
   gpc1_1 gpc3664 (
      {stage2_9[59]},
      {stage3_9[54]}
   );
   gpc1_1 gpc3665 (
      {stage2_9[60]},
      {stage3_9[55]}
   );
   gpc1_1 gpc3666 (
      {stage2_9[61]},
      {stage3_9[56]}
   );
   gpc1_1 gpc3667 (
      {stage2_9[62]},
      {stage3_9[57]}
   );
   gpc1_1 gpc3668 (
      {stage2_9[63]},
      {stage3_9[58]}
   );
   gpc1_1 gpc3669 (
      {stage2_9[64]},
      {stage3_9[59]}
   );
   gpc1_1 gpc3670 (
      {stage2_9[65]},
      {stage3_9[60]}
   );
   gpc1_1 gpc3671 (
      {stage2_9[66]},
      {stage3_9[61]}
   );
   gpc1_1 gpc3672 (
      {stage2_9[67]},
      {stage3_9[62]}
   );
   gpc1_1 gpc3673 (
      {stage2_9[68]},
      {stage3_9[63]}
   );
   gpc1_1 gpc3674 (
      {stage2_9[69]},
      {stage3_9[64]}
   );
   gpc1_1 gpc3675 (
      {stage2_9[70]},
      {stage3_9[65]}
   );
   gpc1_1 gpc3676 (
      {stage2_9[71]},
      {stage3_9[66]}
   );
   gpc1_1 gpc3677 (
      {stage2_9[72]},
      {stage3_9[67]}
   );
   gpc1_1 gpc3678 (
      {stage2_9[73]},
      {stage3_9[68]}
   );
   gpc1_1 gpc3679 (
      {stage2_9[74]},
      {stage3_9[69]}
   );
   gpc1_1 gpc3680 (
      {stage2_10[88]},
      {stage3_10[28]}
   );
   gpc1_1 gpc3681 (
      {stage2_11[80]},
      {stage3_11[32]}
   );
   gpc1_1 gpc3682 (
      {stage2_11[81]},
      {stage3_11[33]}
   );
   gpc1_1 gpc3683 (
      {stage2_11[82]},
      {stage3_11[34]}
   );
   gpc1_1 gpc3684 (
      {stage2_11[83]},
      {stage3_11[35]}
   );
   gpc1_1 gpc3685 (
      {stage2_11[84]},
      {stage3_11[36]}
   );
   gpc1_1 gpc3686 (
      {stage2_11[85]},
      {stage3_11[37]}
   );
   gpc1_1 gpc3687 (
      {stage2_11[86]},
      {stage3_11[38]}
   );
   gpc1_1 gpc3688 (
      {stage2_11[87]},
      {stage3_11[39]}
   );
   gpc1_1 gpc3689 (
      {stage2_11[88]},
      {stage3_11[40]}
   );
   gpc1_1 gpc3690 (
      {stage2_11[89]},
      {stage3_11[41]}
   );
   gpc1_1 gpc3691 (
      {stage2_11[90]},
      {stage3_11[42]}
   );
   gpc1_1 gpc3692 (
      {stage2_11[91]},
      {stage3_11[43]}
   );
   gpc1_1 gpc3693 (
      {stage2_12[102]},
      {stage3_12[41]}
   );
   gpc1_1 gpc3694 (
      {stage2_13[95]},
      {stage3_13[34]}
   );
   gpc1_1 gpc3695 (
      {stage2_13[96]},
      {stage3_13[35]}
   );
   gpc1_1 gpc3696 (
      {stage2_13[97]},
      {stage3_13[36]}
   );
   gpc1_1 gpc3697 (
      {stage2_13[98]},
      {stage3_13[37]}
   );
   gpc1_1 gpc3698 (
      {stage2_13[99]},
      {stage3_13[38]}
   );
   gpc1_1 gpc3699 (
      {stage2_13[100]},
      {stage3_13[39]}
   );
   gpc1_1 gpc3700 (
      {stage2_13[101]},
      {stage3_13[40]}
   );
   gpc1_1 gpc3701 (
      {stage2_14[133]},
      {stage3_14[45]}
   );
   gpc1_1 gpc3702 (
      {stage2_14[134]},
      {stage3_14[46]}
   );
   gpc1_1 gpc3703 (
      {stage2_14[135]},
      {stage3_14[47]}
   );
   gpc1_1 gpc3704 (
      {stage2_14[136]},
      {stage3_14[48]}
   );
   gpc1_1 gpc3705 (
      {stage2_14[137]},
      {stage3_14[49]}
   );
   gpc1_1 gpc3706 (
      {stage2_14[138]},
      {stage3_14[50]}
   );
   gpc1_1 gpc3707 (
      {stage2_15[95]},
      {stage3_15[49]}
   );
   gpc1_1 gpc3708 (
      {stage2_15[96]},
      {stage3_15[50]}
   );
   gpc1_1 gpc3709 (
      {stage2_15[97]},
      {stage3_15[51]}
   );
   gpc1_1 gpc3710 (
      {stage2_15[98]},
      {stage3_15[52]}
   );
   gpc1_1 gpc3711 (
      {stage2_15[99]},
      {stage3_15[53]}
   );
   gpc1_1 gpc3712 (
      {stage2_15[100]},
      {stage3_15[54]}
   );
   gpc1_1 gpc3713 (
      {stage2_15[101]},
      {stage3_15[55]}
   );
   gpc1_1 gpc3714 (
      {stage2_15[102]},
      {stage3_15[56]}
   );
   gpc1_1 gpc3715 (
      {stage2_15[103]},
      {stage3_15[57]}
   );
   gpc1_1 gpc3716 (
      {stage2_15[104]},
      {stage3_15[58]}
   );
   gpc1_1 gpc3717 (
      {stage2_15[105]},
      {stage3_15[59]}
   );
   gpc1_1 gpc3718 (
      {stage2_15[106]},
      {stage3_15[60]}
   );
   gpc1_1 gpc3719 (
      {stage2_15[107]},
      {stage3_15[61]}
   );
   gpc1_1 gpc3720 (
      {stage2_15[108]},
      {stage3_15[62]}
   );
   gpc1_1 gpc3721 (
      {stage2_15[109]},
      {stage3_15[63]}
   );
   gpc1_1 gpc3722 (
      {stage2_15[110]},
      {stage3_15[64]}
   );
   gpc1_1 gpc3723 (
      {stage2_15[111]},
      {stage3_15[65]}
   );
   gpc1_1 gpc3724 (
      {stage2_15[112]},
      {stage3_15[66]}
   );
   gpc1_1 gpc3725 (
      {stage2_15[113]},
      {stage3_15[67]}
   );
   gpc1_1 gpc3726 (
      {stage2_15[114]},
      {stage3_15[68]}
   );
   gpc1_1 gpc3727 (
      {stage2_15[115]},
      {stage3_15[69]}
   );
   gpc1_1 gpc3728 (
      {stage2_15[116]},
      {stage3_15[70]}
   );
   gpc1_1 gpc3729 (
      {stage2_15[117]},
      {stage3_15[71]}
   );
   gpc1_1 gpc3730 (
      {stage2_15[118]},
      {stage3_15[72]}
   );
   gpc1_1 gpc3731 (
      {stage2_15[119]},
      {stage3_15[73]}
   );
   gpc1_1 gpc3732 (
      {stage2_15[120]},
      {stage3_15[74]}
   );
   gpc1_1 gpc3733 (
      {stage2_15[121]},
      {stage3_15[75]}
   );
   gpc1_1 gpc3734 (
      {stage2_15[122]},
      {stage3_15[76]}
   );
   gpc1_1 gpc3735 (
      {stage2_15[123]},
      {stage3_15[77]}
   );
   gpc1_1 gpc3736 (
      {stage2_15[124]},
      {stage3_15[78]}
   );
   gpc1_1 gpc3737 (
      {stage2_15[125]},
      {stage3_15[79]}
   );
   gpc1_1 gpc3738 (
      {stage2_15[126]},
      {stage3_15[80]}
   );
   gpc1_1 gpc3739 (
      {stage2_15[127]},
      {stage3_15[81]}
   );
   gpc1_1 gpc3740 (
      {stage2_15[128]},
      {stage3_15[82]}
   );
   gpc1_1 gpc3741 (
      {stage2_15[129]},
      {stage3_15[83]}
   );
   gpc1_1 gpc3742 (
      {stage2_15[130]},
      {stage3_15[84]}
   );
   gpc1_1 gpc3743 (
      {stage2_15[131]},
      {stage3_15[85]}
   );
   gpc1_1 gpc3744 (
      {stage2_15[132]},
      {stage3_15[86]}
   );
   gpc1_1 gpc3745 (
      {stage2_15[133]},
      {stage3_15[87]}
   );
   gpc1_1 gpc3746 (
      {stage2_15[134]},
      {stage3_15[88]}
   );
   gpc1_1 gpc3747 (
      {stage2_15[135]},
      {stage3_15[89]}
   );
   gpc1_1 gpc3748 (
      {stage2_16[81]},
      {stage3_16[39]}
   );
   gpc1_1 gpc3749 (
      {stage2_16[82]},
      {stage3_16[40]}
   );
   gpc1_1 gpc3750 (
      {stage2_16[83]},
      {stage3_16[41]}
   );
   gpc1_1 gpc3751 (
      {stage2_16[84]},
      {stage3_16[42]}
   );
   gpc1_1 gpc3752 (
      {stage2_16[85]},
      {stage3_16[43]}
   );
   gpc1_1 gpc3753 (
      {stage2_16[86]},
      {stage3_16[44]}
   );
   gpc1_1 gpc3754 (
      {stage2_16[87]},
      {stage3_16[45]}
   );
   gpc1_1 gpc3755 (
      {stage2_16[88]},
      {stage3_16[46]}
   );
   gpc1_1 gpc3756 (
      {stage2_16[89]},
      {stage3_16[47]}
   );
   gpc1_1 gpc3757 (
      {stage2_16[90]},
      {stage3_16[48]}
   );
   gpc1_1 gpc3758 (
      {stage2_16[91]},
      {stage3_16[49]}
   );
   gpc1_1 gpc3759 (
      {stage2_16[92]},
      {stage3_16[50]}
   );
   gpc1_1 gpc3760 (
      {stage2_16[93]},
      {stage3_16[51]}
   );
   gpc1_1 gpc3761 (
      {stage2_16[94]},
      {stage3_16[52]}
   );
   gpc1_1 gpc3762 (
      {stage2_16[95]},
      {stage3_16[53]}
   );
   gpc1_1 gpc3763 (
      {stage2_16[96]},
      {stage3_16[54]}
   );
   gpc1_1 gpc3764 (
      {stage2_16[97]},
      {stage3_16[55]}
   );
   gpc1_1 gpc3765 (
      {stage2_16[98]},
      {stage3_16[56]}
   );
   gpc1_1 gpc3766 (
      {stage2_16[99]},
      {stage3_16[57]}
   );
   gpc1_1 gpc3767 (
      {stage2_16[100]},
      {stage3_16[58]}
   );
   gpc1_1 gpc3768 (
      {stage2_16[101]},
      {stage3_16[59]}
   );
   gpc1_1 gpc3769 (
      {stage2_16[102]},
      {stage3_16[60]}
   );
   gpc1_1 gpc3770 (
      {stage2_16[103]},
      {stage3_16[61]}
   );
   gpc1_1 gpc3771 (
      {stage2_17[109]},
      {stage3_17[37]}
   );
   gpc1_1 gpc3772 (
      {stage2_17[110]},
      {stage3_17[38]}
   );
   gpc1_1 gpc3773 (
      {stage2_17[111]},
      {stage3_17[39]}
   );
   gpc1_1 gpc3774 (
      {stage2_17[112]},
      {stage3_17[40]}
   );
   gpc1_1 gpc3775 (
      {stage2_17[113]},
      {stage3_17[41]}
   );
   gpc1_1 gpc3776 (
      {stage2_17[114]},
      {stage3_17[42]}
   );
   gpc1_1 gpc3777 (
      {stage2_17[115]},
      {stage3_17[43]}
   );
   gpc1_1 gpc3778 (
      {stage2_17[116]},
      {stage3_17[44]}
   );
   gpc1_1 gpc3779 (
      {stage2_17[117]},
      {stage3_17[45]}
   );
   gpc1_1 gpc3780 (
      {stage2_17[118]},
      {stage3_17[46]}
   );
   gpc1_1 gpc3781 (
      {stage2_17[119]},
      {stage3_17[47]}
   );
   gpc1_1 gpc3782 (
      {stage2_17[120]},
      {stage3_17[48]}
   );
   gpc1_1 gpc3783 (
      {stage2_17[121]},
      {stage3_17[49]}
   );
   gpc1_1 gpc3784 (
      {stage2_18[80]},
      {stage3_18[48]}
   );
   gpc1_1 gpc3785 (
      {stage2_18[81]},
      {stage3_18[49]}
   );
   gpc1_1 gpc3786 (
      {stage2_19[98]},
      {stage3_19[38]}
   );
   gpc1_1 gpc3787 (
      {stage2_19[99]},
      {stage3_19[39]}
   );
   gpc1_1 gpc3788 (
      {stage2_19[100]},
      {stage3_19[40]}
   );
   gpc1_1 gpc3789 (
      {stage2_19[101]},
      {stage3_19[41]}
   );
   gpc1_1 gpc3790 (
      {stage2_19[102]},
      {stage3_19[42]}
   );
   gpc1_1 gpc3791 (
      {stage2_19[103]},
      {stage3_19[43]}
   );
   gpc1_1 gpc3792 (
      {stage2_19[104]},
      {stage3_19[44]}
   );
   gpc1_1 gpc3793 (
      {stage2_19[105]},
      {stage3_19[45]}
   );
   gpc1_1 gpc3794 (
      {stage2_19[106]},
      {stage3_19[46]}
   );
   gpc1_1 gpc3795 (
      {stage2_19[107]},
      {stage3_19[47]}
   );
   gpc1_1 gpc3796 (
      {stage2_19[108]},
      {stage3_19[48]}
   );
   gpc1_1 gpc3797 (
      {stage2_19[109]},
      {stage3_19[49]}
   );
   gpc1_1 gpc3798 (
      {stage2_20[116]},
      {stage3_20[34]}
   );
   gpc1_1 gpc3799 (
      {stage2_20[117]},
      {stage3_20[35]}
   );
   gpc1_1 gpc3800 (
      {stage2_20[118]},
      {stage3_20[36]}
   );
   gpc1_1 gpc3801 (
      {stage2_20[119]},
      {stage3_20[37]}
   );
   gpc1_1 gpc3802 (
      {stage2_20[120]},
      {stage3_20[38]}
   );
   gpc1_1 gpc3803 (
      {stage2_20[121]},
      {stage3_20[39]}
   );
   gpc1_1 gpc3804 (
      {stage2_20[122]},
      {stage3_20[40]}
   );
   gpc1_1 gpc3805 (
      {stage2_20[123]},
      {stage3_20[41]}
   );
   gpc1_1 gpc3806 (
      {stage2_20[124]},
      {stage3_20[42]}
   );
   gpc1_1 gpc3807 (
      {stage2_20[125]},
      {stage3_20[43]}
   );
   gpc1_1 gpc3808 (
      {stage2_20[126]},
      {stage3_20[44]}
   );
   gpc1_1 gpc3809 (
      {stage2_20[127]},
      {stage3_20[45]}
   );
   gpc1_1 gpc3810 (
      {stage2_21[64]},
      {stage3_21[44]}
   );
   gpc1_1 gpc3811 (
      {stage2_21[65]},
      {stage3_21[45]}
   );
   gpc1_1 gpc3812 (
      {stage2_21[66]},
      {stage3_21[46]}
   );
   gpc1_1 gpc3813 (
      {stage2_21[67]},
      {stage3_21[47]}
   );
   gpc1_1 gpc3814 (
      {stage2_21[68]},
      {stage3_21[48]}
   );
   gpc1_1 gpc3815 (
      {stage2_21[69]},
      {stage3_21[49]}
   );
   gpc1_1 gpc3816 (
      {stage2_21[70]},
      {stage3_21[50]}
   );
   gpc1_1 gpc3817 (
      {stage2_21[71]},
      {stage3_21[51]}
   );
   gpc1_1 gpc3818 (
      {stage2_21[72]},
      {stage3_21[52]}
   );
   gpc1_1 gpc3819 (
      {stage2_21[73]},
      {stage3_21[53]}
   );
   gpc1_1 gpc3820 (
      {stage2_21[74]},
      {stage3_21[54]}
   );
   gpc1_1 gpc3821 (
      {stage2_21[75]},
      {stage3_21[55]}
   );
   gpc1_1 gpc3822 (
      {stage2_21[76]},
      {stage3_21[56]}
   );
   gpc1_1 gpc3823 (
      {stage2_21[77]},
      {stage3_21[57]}
   );
   gpc1_1 gpc3824 (
      {stage2_21[78]},
      {stage3_21[58]}
   );
   gpc1_1 gpc3825 (
      {stage2_22[66]},
      {stage3_22[34]}
   );
   gpc1_1 gpc3826 (
      {stage2_22[67]},
      {stage3_22[35]}
   );
   gpc1_1 gpc3827 (
      {stage2_22[68]},
      {stage3_22[36]}
   );
   gpc1_1 gpc3828 (
      {stage2_22[69]},
      {stage3_22[37]}
   );
   gpc1_1 gpc3829 (
      {stage2_22[70]},
      {stage3_22[38]}
   );
   gpc1_1 gpc3830 (
      {stage2_22[71]},
      {stage3_22[39]}
   );
   gpc1_1 gpc3831 (
      {stage2_22[72]},
      {stage3_22[40]}
   );
   gpc1_1 gpc3832 (
      {stage2_22[73]},
      {stage3_22[41]}
   );
   gpc1_1 gpc3833 (
      {stage2_22[74]},
      {stage3_22[42]}
   );
   gpc1_1 gpc3834 (
      {stage2_22[75]},
      {stage3_22[43]}
   );
   gpc1_1 gpc3835 (
      {stage2_22[76]},
      {stage3_22[44]}
   );
   gpc1_1 gpc3836 (
      {stage2_22[77]},
      {stage3_22[45]}
   );
   gpc1_1 gpc3837 (
      {stage2_22[78]},
      {stage3_22[46]}
   );
   gpc1_1 gpc3838 (
      {stage2_23[91]},
      {stage3_23[29]}
   );
   gpc1_1 gpc3839 (
      {stage2_23[92]},
      {stage3_23[30]}
   );
   gpc1_1 gpc3840 (
      {stage2_23[93]},
      {stage3_23[31]}
   );
   gpc1_1 gpc3841 (
      {stage2_23[94]},
      {stage3_23[32]}
   );
   gpc1_1 gpc3842 (
      {stage2_23[95]},
      {stage3_23[33]}
   );
   gpc1_1 gpc3843 (
      {stage2_23[96]},
      {stage3_23[34]}
   );
   gpc1_1 gpc3844 (
      {stage2_23[97]},
      {stage3_23[35]}
   );
   gpc1_1 gpc3845 (
      {stage2_23[98]},
      {stage3_23[36]}
   );
   gpc1_1 gpc3846 (
      {stage2_23[99]},
      {stage3_23[37]}
   );
   gpc1_1 gpc3847 (
      {stage2_23[100]},
      {stage3_23[38]}
   );
   gpc1_1 gpc3848 (
      {stage2_23[101]},
      {stage3_23[39]}
   );
   gpc1_1 gpc3849 (
      {stage2_23[102]},
      {stage3_23[40]}
   );
   gpc1_1 gpc3850 (
      {stage2_23[103]},
      {stage3_23[41]}
   );
   gpc1_1 gpc3851 (
      {stage2_23[104]},
      {stage3_23[42]}
   );
   gpc1_1 gpc3852 (
      {stage2_23[105]},
      {stage3_23[43]}
   );
   gpc1_1 gpc3853 (
      {stage2_23[106]},
      {stage3_23[44]}
   );
   gpc1_1 gpc3854 (
      {stage2_23[107]},
      {stage3_23[45]}
   );
   gpc1_1 gpc3855 (
      {stage2_23[108]},
      {stage3_23[46]}
   );
   gpc1_1 gpc3856 (
      {stage2_23[109]},
      {stage3_23[47]}
   );
   gpc1_1 gpc3857 (
      {stage2_27[70]},
      {stage3_27[40]}
   );
   gpc1_1 gpc3858 (
      {stage2_27[71]},
      {stage3_27[41]}
   );
   gpc1_1 gpc3859 (
      {stage2_27[72]},
      {stage3_27[42]}
   );
   gpc1_1 gpc3860 (
      {stage2_27[73]},
      {stage3_27[43]}
   );
   gpc1_1 gpc3861 (
      {stage2_27[74]},
      {stage3_27[44]}
   );
   gpc1_1 gpc3862 (
      {stage2_27[75]},
      {stage3_27[45]}
   );
   gpc1_1 gpc3863 (
      {stage2_27[76]},
      {stage3_27[46]}
   );
   gpc1_1 gpc3864 (
      {stage2_27[77]},
      {stage3_27[47]}
   );
   gpc1_1 gpc3865 (
      {stage2_27[78]},
      {stage3_27[48]}
   );
   gpc1_1 gpc3866 (
      {stage2_27[79]},
      {stage3_27[49]}
   );
   gpc1_1 gpc3867 (
      {stage2_27[80]},
      {stage3_27[50]}
   );
   gpc1_1 gpc3868 (
      {stage2_27[81]},
      {stage3_27[51]}
   );
   gpc1_1 gpc3869 (
      {stage2_27[82]},
      {stage3_27[52]}
   );
   gpc1_1 gpc3870 (
      {stage2_27[83]},
      {stage3_27[53]}
   );
   gpc1_1 gpc3871 (
      {stage2_27[84]},
      {stage3_27[54]}
   );
   gpc1_1 gpc3872 (
      {stage2_27[85]},
      {stage3_27[55]}
   );
   gpc1_1 gpc3873 (
      {stage2_27[86]},
      {stage3_27[56]}
   );
   gpc1_1 gpc3874 (
      {stage2_27[87]},
      {stage3_27[57]}
   );
   gpc1_1 gpc3875 (
      {stage2_27[88]},
      {stage3_27[58]}
   );
   gpc1_1 gpc3876 (
      {stage2_27[89]},
      {stage3_27[59]}
   );
   gpc1_1 gpc3877 (
      {stage2_27[90]},
      {stage3_27[60]}
   );
   gpc1_1 gpc3878 (
      {stage2_27[91]},
      {stage3_27[61]}
   );
   gpc1_1 gpc3879 (
      {stage2_27[92]},
      {stage3_27[62]}
   );
   gpc1_1 gpc3880 (
      {stage2_27[93]},
      {stage3_27[63]}
   );
   gpc1_1 gpc3881 (
      {stage2_27[94]},
      {stage3_27[64]}
   );
   gpc1_1 gpc3882 (
      {stage2_27[95]},
      {stage3_27[65]}
   );
   gpc1_1 gpc3883 (
      {stage2_27[96]},
      {stage3_27[66]}
   );
   gpc1_1 gpc3884 (
      {stage2_28[69]},
      {stage3_28[37]}
   );
   gpc1_1 gpc3885 (
      {stage2_28[70]},
      {stage3_28[38]}
   );
   gpc1_1 gpc3886 (
      {stage2_28[71]},
      {stage3_28[39]}
   );
   gpc1_1 gpc3887 (
      {stage2_28[72]},
      {stage3_28[40]}
   );
   gpc1_1 gpc3888 (
      {stage2_28[73]},
      {stage3_28[41]}
   );
   gpc1_1 gpc3889 (
      {stage2_28[74]},
      {stage3_28[42]}
   );
   gpc1_1 gpc3890 (
      {stage2_29[119]},
      {stage3_29[37]}
   );
   gpc1_1 gpc3891 (
      {stage2_29[120]},
      {stage3_29[38]}
   );
   gpc1_1 gpc3892 (
      {stage2_30[108]},
      {stage3_30[38]}
   );
   gpc1_1 gpc3893 (
      {stage2_30[109]},
      {stage3_30[39]}
   );
   gpc1_1 gpc3894 (
      {stage2_30[110]},
      {stage3_30[40]}
   );
   gpc1_1 gpc3895 (
      {stage2_30[111]},
      {stage3_30[41]}
   );
   gpc1_1 gpc3896 (
      {stage2_30[112]},
      {stage3_30[42]}
   );
   gpc1_1 gpc3897 (
      {stage2_30[113]},
      {stage3_30[43]}
   );
   gpc1_1 gpc3898 (
      {stage2_30[114]},
      {stage3_30[44]}
   );
   gpc1_1 gpc3899 (
      {stage2_30[115]},
      {stage3_30[45]}
   );
   gpc1_1 gpc3900 (
      {stage2_30[116]},
      {stage3_30[46]}
   );
   gpc1_1 gpc3901 (
      {stage2_30[117]},
      {stage3_30[47]}
   );
   gpc1_1 gpc3902 (
      {stage2_30[118]},
      {stage3_30[48]}
   );
   gpc1_1 gpc3903 (
      {stage2_30[119]},
      {stage3_30[49]}
   );
   gpc1_1 gpc3904 (
      {stage2_30[120]},
      {stage3_30[50]}
   );
   gpc1_1 gpc3905 (
      {stage2_30[121]},
      {stage3_30[51]}
   );
   gpc1_1 gpc3906 (
      {stage2_30[122]},
      {stage3_30[52]}
   );
   gpc1_1 gpc3907 (
      {stage2_30[123]},
      {stage3_30[53]}
   );
   gpc1_1 gpc3908 (
      {stage2_30[124]},
      {stage3_30[54]}
   );
   gpc1_1 gpc3909 (
      {stage2_30[125]},
      {stage3_30[55]}
   );
   gpc1_1 gpc3910 (
      {stage2_30[126]},
      {stage3_30[56]}
   );
   gpc1_1 gpc3911 (
      {stage2_30[127]},
      {stage3_30[57]}
   );
   gpc1_1 gpc3912 (
      {stage2_30[128]},
      {stage3_30[58]}
   );
   gpc1_1 gpc3913 (
      {stage2_30[129]},
      {stage3_30[59]}
   );
   gpc1_1 gpc3914 (
      {stage2_31[83]},
      {stage3_31[39]}
   );
   gpc1_1 gpc3915 (
      {stage2_33[36]},
      {stage3_33[30]}
   );
   gpc1_1 gpc3916 (
      {stage2_33[37]},
      {stage3_33[31]}
   );
   gpc1_1 gpc3917 (
      {stage2_33[38]},
      {stage3_33[32]}
   );
   gpc1_1 gpc3918 (
      {stage2_33[39]},
      {stage3_33[33]}
   );
   gpc1_1 gpc3919 (
      {stage2_33[40]},
      {stage3_33[34]}
   );
   gpc1_1 gpc3920 (
      {stage2_33[41]},
      {stage3_33[35]}
   );
   gpc1_1 gpc3921 (
      {stage2_33[42]},
      {stage3_33[36]}
   );
   gpc1_1 gpc3922 (
      {stage2_33[43]},
      {stage3_33[37]}
   );
   gpc1_1 gpc3923 (
      {stage2_33[44]},
      {stage3_33[38]}
   );
   gpc1_1 gpc3924 (
      {stage2_33[45]},
      {stage3_33[39]}
   );
   gpc1_1 gpc3925 (
      {stage2_34[30]},
      {stage3_34[16]}
   );
   gpc1_1 gpc3926 (
      {stage2_34[31]},
      {stage3_34[17]}
   );
   gpc1_1 gpc3927 (
      {stage2_34[32]},
      {stage3_34[18]}
   );
   gpc1_1 gpc3928 (
      {stage2_34[33]},
      {stage3_34[19]}
   );
   gpc1_1 gpc3929 (
      {stage2_34[34]},
      {stage3_34[20]}
   );
   gpc1_1 gpc3930 (
      {stage2_34[35]},
      {stage3_34[21]}
   );
   gpc1_1 gpc3931 (
      {stage2_35[12]},
      {stage3_35[11]}
   );
   gpc1_1 gpc3932 (
      {stage2_35[13]},
      {stage3_35[12]}
   );
   gpc606_5 gpc3933 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc3934 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc3935 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc3936 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10], stage3_2[11]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[2],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc606_5 gpc3937 (
      {stage3_2[12], stage3_2[13], stage3_2[14], stage3_2[15], stage3_2[16], stage3_2[17]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[3],stage4_4[4],stage4_3[4],stage4_2[4]}
   );
   gpc606_5 gpc3938 (
      {stage3_2[18], stage3_2[19], stage3_2[20], stage3_2[21], stage3_2[22], stage3_2[23]},
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17]},
      {stage4_6[2],stage4_5[4],stage4_4[5],stage4_3[5],stage4_2[5]}
   );
   gpc606_5 gpc3939 (
      {stage3_2[24], stage3_2[25], stage3_2[26], stage3_2[27], stage3_2[28], stage3_2[29]},
      {stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22], stage3_4[23]},
      {stage4_6[3],stage4_5[5],stage4_4[6],stage4_3[6],stage4_2[6]}
   );
   gpc615_5 gpc3940 (
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16]},
      {stage3_4[24]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[4],stage4_5[6],stage4_4[7],stage4_3[7]}
   );
   gpc615_5 gpc3941 (
      {stage3_3[17], stage3_3[18], stage3_3[19], stage3_3[20], stage3_3[21]},
      {stage3_4[25]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[5],stage4_5[7],stage4_4[8],stage4_3[8]}
   );
   gpc615_5 gpc3942 (
      {stage3_3[22], stage3_3[23], stage3_3[24], stage3_3[25], stage3_3[26]},
      {stage3_4[26]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage4_7[2],stage4_6[6],stage4_5[8],stage4_4[9],stage4_3[9]}
   );
   gpc606_5 gpc3943 (
      {stage3_4[27], stage3_4[28], stage3_4[29], stage3_4[30], stage3_4[31], stage3_4[32]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[3],stage4_6[7],stage4_5[9],stage4_4[10]}
   );
   gpc606_5 gpc3944 (
      {stage3_4[33], stage3_4[34], stage3_4[35], stage3_4[36], stage3_4[37], stage3_4[38]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[4],stage4_6[8],stage4_5[10],stage4_4[11]}
   );
   gpc1163_5 gpc3945 (
      {stage3_5[18], stage3_5[19], stage3_5[20]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage3_7[0]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[2],stage4_7[5],stage4_6[9],stage4_5[11]}
   );
   gpc1163_5 gpc3946 (
      {stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage3_7[1]},
      {stage3_8[1]},
      {stage4_9[1],stage4_8[3],stage4_7[6],stage4_6[10],stage4_5[12]}
   );
   gpc606_5 gpc3947 (
      {stage3_5[24], stage3_5[25], stage3_5[26], stage3_5[27], stage3_5[28], stage3_5[29]},
      {stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage4_9[2],stage4_8[4],stage4_7[7],stage4_6[11],stage4_5[13]}
   );
   gpc606_5 gpc3948 (
      {stage3_5[30], stage3_5[31], stage3_5[32], stage3_5[33], stage3_5[34], stage3_5[35]},
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13]},
      {stage4_9[3],stage4_8[5],stage4_7[8],stage4_6[12],stage4_5[14]}
   );
   gpc606_5 gpc3949 (
      {stage3_5[36], stage3_5[37], stage3_5[38], stage3_5[39], stage3_5[40], stage3_5[41]},
      {stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17], stage3_7[18], stage3_7[19]},
      {stage4_9[4],stage4_8[6],stage4_7[9],stage4_6[13],stage4_5[15]}
   );
   gpc615_5 gpc3950 (
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28]},
      {stage3_7[20]},
      {stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5], stage3_8[6], stage3_8[7]},
      {stage4_10[0],stage4_9[5],stage4_8[7],stage4_7[10],stage4_6[14]}
   );
   gpc615_5 gpc3951 (
      {stage3_6[29], stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33]},
      {stage3_7[21]},
      {stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11], stage3_8[12], stage3_8[13]},
      {stage4_10[1],stage4_9[6],stage4_8[8],stage4_7[11],stage4_6[15]}
   );
   gpc615_5 gpc3952 (
      {stage3_6[34], stage3_6[35], stage3_6[36], stage3_6[37], stage3_6[38]},
      {stage3_7[22]},
      {stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17], stage3_8[18], stage3_8[19]},
      {stage4_10[2],stage4_9[7],stage4_8[9],stage4_7[12],stage4_6[16]}
   );
   gpc615_5 gpc3953 (
      {stage3_7[23], stage3_7[24], stage3_7[25], stage3_7[26], stage3_7[27]},
      {stage3_8[20]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[3],stage4_9[8],stage4_8[10],stage4_7[13]}
   );
   gpc615_5 gpc3954 (
      {stage3_7[28], stage3_7[29], stage3_7[30], stage3_7[31], stage3_7[32]},
      {stage3_8[21]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[4],stage4_9[9],stage4_8[11],stage4_7[14]}
   );
   gpc615_5 gpc3955 (
      {stage3_7[33], stage3_7[34], stage3_7[35], stage3_7[36], stage3_7[37]},
      {stage3_8[22]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[5],stage4_9[10],stage4_8[12],stage4_7[15]}
   );
   gpc615_5 gpc3956 (
      {stage3_7[38], stage3_7[39], stage3_7[40], stage3_7[41], stage3_7[42]},
      {stage3_8[23]},
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage4_11[3],stage4_10[6],stage4_9[11],stage4_8[13],stage4_7[16]}
   );
   gpc615_5 gpc3957 (
      {stage3_7[43], stage3_7[44], stage3_7[45], stage3_7[46], stage3_7[47]},
      {stage3_8[24]},
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage4_11[4],stage4_10[7],stage4_9[12],stage4_8[14],stage4_7[17]}
   );
   gpc615_5 gpc3958 (
      {stage3_7[48], stage3_7[49], stage3_7[50], stage3_7[51], stage3_7[52]},
      {stage3_8[25]},
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage4_11[5],stage4_10[8],stage4_9[13],stage4_8[15],stage4_7[18]}
   );
   gpc615_5 gpc3959 (
      {stage3_7[53], stage3_7[54], stage3_7[55], stage3_7[56], stage3_7[57]},
      {stage3_8[26]},
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage4_11[6],stage4_10[9],stage4_9[14],stage4_8[16],stage4_7[19]}
   );
   gpc615_5 gpc3960 (
      {stage3_7[58], stage3_7[59], stage3_7[60], stage3_7[61], stage3_7[62]},
      {stage3_8[27]},
      {stage3_9[42], stage3_9[43], stage3_9[44], stage3_9[45], stage3_9[46], stage3_9[47]},
      {stage4_11[7],stage4_10[10],stage4_9[15],stage4_8[17],stage4_7[20]}
   );
   gpc606_5 gpc3961 (
      {stage3_8[28], stage3_8[29], stage3_8[30], stage3_8[31], stage3_8[32], stage3_8[33]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[8],stage4_10[11],stage4_9[16],stage4_8[18]}
   );
   gpc623_5 gpc3962 (
      {stage3_9[48], stage3_9[49], stage3_9[50]},
      {stage3_10[6], stage3_10[7]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[1],stage4_11[9],stage4_10[12],stage4_9[17]}
   );
   gpc623_5 gpc3963 (
      {stage3_9[51], stage3_9[52], stage3_9[53]},
      {stage3_10[8], stage3_10[9]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[2],stage4_11[10],stage4_10[13],stage4_9[18]}
   );
   gpc623_5 gpc3964 (
      {stage3_9[54], stage3_9[55], stage3_9[56]},
      {stage3_10[10], stage3_10[11]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[3],stage4_11[11],stage4_10[14],stage4_9[19]}
   );
   gpc623_5 gpc3965 (
      {stage3_9[57], stage3_9[58], stage3_9[59]},
      {stage3_10[12], stage3_10[13]},
      {stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage4_13[3],stage4_12[4],stage4_11[12],stage4_10[15],stage4_9[20]}
   );
   gpc623_5 gpc3966 (
      {stage3_9[60], stage3_9[61], stage3_9[62]},
      {stage3_10[14], stage3_10[15]},
      {stage3_11[24], stage3_11[25], stage3_11[26], stage3_11[27], stage3_11[28], stage3_11[29]},
      {stage4_13[4],stage4_12[5],stage4_11[13],stage4_10[16],stage4_9[21]}
   );
   gpc623_5 gpc3967 (
      {stage3_9[63], stage3_9[64], stage3_9[65]},
      {stage3_10[16], stage3_10[17]},
      {stage3_11[30], stage3_11[31], stage3_11[32], stage3_11[33], stage3_11[34], stage3_11[35]},
      {stage4_13[5],stage4_12[6],stage4_11[14],stage4_10[17],stage4_9[22]}
   );
   gpc1163_5 gpc3968 (
      {stage3_11[36], stage3_11[37], stage3_11[38]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[0]},
      {stage3_14[0]},
      {stage4_15[0],stage4_14[0],stage4_13[6],stage4_12[7],stage4_11[15]}
   );
   gpc606_5 gpc3969 (
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6]},
      {stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[7],stage4_12[8]}
   );
   gpc606_5 gpc3970 (
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11], stage3_14[12]},
      {stage4_16[1],stage4_15[2],stage4_14[2],stage4_13[8],stage4_12[9]}
   );
   gpc606_5 gpc3971 (
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17], stage3_14[18]},
      {stage4_16[2],stage4_15[3],stage4_14[3],stage4_13[9],stage4_12[10]}
   );
   gpc606_5 gpc3972 (
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23], stage3_14[24]},
      {stage4_16[3],stage4_15[4],stage4_14[4],stage4_13[10],stage4_12[11]}
   );
   gpc606_5 gpc3973 (
      {stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35]},
      {stage3_14[25], stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29], stage3_14[30]},
      {stage4_16[4],stage4_15[5],stage4_14[5],stage4_13[11],stage4_12[12]}
   );
   gpc606_5 gpc3974 (
      {stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40], stage3_12[41]},
      {stage3_14[31], stage3_14[32], stage3_14[33], stage3_14[34], stage3_14[35], stage3_14[36]},
      {stage4_16[5],stage4_15[6],stage4_14[6],stage4_13[12],stage4_12[13]}
   );
   gpc2135_5 gpc3975 (
      {stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_14[37], stage3_14[38], stage3_14[39]},
      {stage3_15[0]},
      {stage3_16[0], stage3_16[1]},
      {stage4_17[0],stage4_16[6],stage4_15[7],stage4_14[7],stage4_13[13]}
   );
   gpc2135_5 gpc3976 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10]},
      {stage3_14[40], stage3_14[41], stage3_14[42]},
      {stage3_15[1]},
      {stage3_16[2], stage3_16[3]},
      {stage4_17[1],stage4_16[7],stage4_15[8],stage4_14[8],stage4_13[14]}
   );
   gpc2135_5 gpc3977 (
      {stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15]},
      {stage3_14[43], stage3_14[44], stage3_14[45]},
      {stage3_15[2]},
      {stage3_16[4], stage3_16[5]},
      {stage4_17[2],stage4_16[8],stage4_15[9],stage4_14[9],stage4_13[15]}
   );
   gpc2135_5 gpc3978 (
      {stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20]},
      {stage3_14[46], stage3_14[47], stage3_14[48]},
      {stage3_15[3]},
      {stage3_16[6], stage3_16[7]},
      {stage4_17[3],stage4_16[9],stage4_15[10],stage4_14[10],stage4_13[16]}
   );
   gpc2135_5 gpc3979 (
      {stage3_13[21], stage3_13[22], stage3_13[23], stage3_13[24], stage3_13[25]},
      {stage3_14[49], stage3_14[50], 1'b0},
      {stage3_15[4]},
      {stage3_16[8], stage3_16[9]},
      {stage4_17[4],stage4_16[10],stage4_15[11],stage4_14[11],stage4_13[17]}
   );
   gpc606_5 gpc3980 (
      {stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30], stage3_13[31]},
      {stage3_15[5], stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10]},
      {stage4_17[5],stage4_16[11],stage4_15[12],stage4_14[12],stage4_13[18]}
   );
   gpc2135_5 gpc3981 (
      {stage3_15[11], stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15]},
      {stage3_16[10], stage3_16[11], stage3_16[12]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1]},
      {stage4_19[0],stage4_18[0],stage4_17[6],stage4_16[12],stage4_15[13]}
   );
   gpc2135_5 gpc3982 (
      {stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19], stage3_15[20]},
      {stage3_16[13], stage3_16[14], stage3_16[15]},
      {stage3_17[1]},
      {stage3_18[2], stage3_18[3]},
      {stage4_19[1],stage4_18[1],stage4_17[7],stage4_16[13],stage4_15[14]}
   );
   gpc2135_5 gpc3983 (
      {stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25]},
      {stage3_16[16], stage3_16[17], stage3_16[18]},
      {stage3_17[2]},
      {stage3_18[4], stage3_18[5]},
      {stage4_19[2],stage4_18[2],stage4_17[8],stage4_16[14],stage4_15[15]}
   );
   gpc2135_5 gpc3984 (
      {stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29], stage3_15[30]},
      {stage3_16[19], stage3_16[20], stage3_16[21]},
      {stage3_17[3]},
      {stage3_18[6], stage3_18[7]},
      {stage4_19[3],stage4_18[3],stage4_17[9],stage4_16[15],stage4_15[16]}
   );
   gpc2135_5 gpc3985 (
      {stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34], stage3_15[35]},
      {stage3_16[22], stage3_16[23], stage3_16[24]},
      {stage3_17[4]},
      {stage3_18[8], stage3_18[9]},
      {stage4_19[4],stage4_18[4],stage4_17[10],stage4_16[16],stage4_15[17]}
   );
   gpc2135_5 gpc3986 (
      {stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39], stage3_15[40]},
      {stage3_16[25], stage3_16[26], stage3_16[27]},
      {stage3_17[5]},
      {stage3_18[10], stage3_18[11]},
      {stage4_19[5],stage4_18[5],stage4_17[11],stage4_16[17],stage4_15[18]}
   );
   gpc2135_5 gpc3987 (
      {stage3_15[41], stage3_15[42], stage3_15[43], stage3_15[44], stage3_15[45]},
      {stage3_16[28], stage3_16[29], stage3_16[30]},
      {stage3_17[6]},
      {stage3_18[12], stage3_18[13]},
      {stage4_19[6],stage4_18[6],stage4_17[12],stage4_16[18],stage4_15[19]}
   );
   gpc2135_5 gpc3988 (
      {stage3_15[46], stage3_15[47], stage3_15[48], stage3_15[49], stage3_15[50]},
      {stage3_16[31], stage3_16[32], stage3_16[33]},
      {stage3_17[7]},
      {stage3_18[14], stage3_18[15]},
      {stage4_19[7],stage4_18[7],stage4_17[13],stage4_16[19],stage4_15[20]}
   );
   gpc2135_5 gpc3989 (
      {stage3_15[51], stage3_15[52], stage3_15[53], stage3_15[54], stage3_15[55]},
      {stage3_16[34], stage3_16[35], stage3_16[36]},
      {stage3_17[8]},
      {stage3_18[16], stage3_18[17]},
      {stage4_19[8],stage4_18[8],stage4_17[14],stage4_16[20],stage4_15[21]}
   );
   gpc2135_5 gpc3990 (
      {stage3_15[56], stage3_15[57], stage3_15[58], stage3_15[59], stage3_15[60]},
      {stage3_16[37], stage3_16[38], stage3_16[39]},
      {stage3_17[9]},
      {stage3_18[18], stage3_18[19]},
      {stage4_19[9],stage4_18[9],stage4_17[15],stage4_16[21],stage4_15[22]}
   );
   gpc615_5 gpc3991 (
      {stage3_15[61], stage3_15[62], stage3_15[63], stage3_15[64], stage3_15[65]},
      {stage3_16[40]},
      {stage3_17[10], stage3_17[11], stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15]},
      {stage4_19[10],stage4_18[10],stage4_17[16],stage4_16[22],stage4_15[23]}
   );
   gpc606_5 gpc3992 (
      {stage3_16[41], stage3_16[42], stage3_16[43], stage3_16[44], stage3_16[45], stage3_16[46]},
      {stage3_18[20], stage3_18[21], stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25]},
      {stage4_20[0],stage4_19[11],stage4_18[11],stage4_17[17],stage4_16[23]}
   );
   gpc606_5 gpc3993 (
      {stage3_16[47], stage3_16[48], stage3_16[49], stage3_16[50], stage3_16[51], stage3_16[52]},
      {stage3_18[26], stage3_18[27], stage3_18[28], stage3_18[29], stage3_18[30], stage3_18[31]},
      {stage4_20[1],stage4_19[12],stage4_18[12],stage4_17[18],stage4_16[24]}
   );
   gpc606_5 gpc3994 (
      {stage3_16[53], stage3_16[54], stage3_16[55], stage3_16[56], stage3_16[57], stage3_16[58]},
      {stage3_18[32], stage3_18[33], stage3_18[34], stage3_18[35], stage3_18[36], stage3_18[37]},
      {stage4_20[2],stage4_19[13],stage4_18[13],stage4_17[19],stage4_16[25]}
   );
   gpc1163_5 gpc3995 (
      {stage3_17[16], stage3_17[17], stage3_17[18]},
      {stage3_18[38], stage3_18[39], stage3_18[40], stage3_18[41], stage3_18[42], stage3_18[43]},
      {stage3_19[0]},
      {stage3_20[0]},
      {stage4_21[0],stage4_20[3],stage4_19[14],stage4_18[14],stage4_17[20]}
   );
   gpc1163_5 gpc3996 (
      {stage3_17[19], stage3_17[20], stage3_17[21]},
      {stage3_18[44], stage3_18[45], stage3_18[46], stage3_18[47], stage3_18[48], stage3_18[49]},
      {stage3_19[1]},
      {stage3_20[1]},
      {stage4_21[1],stage4_20[4],stage4_19[15],stage4_18[15],stage4_17[21]}
   );
   gpc606_5 gpc3997 (
      {stage3_17[22], stage3_17[23], stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27]},
      {stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6], stage3_19[7]},
      {stage4_21[2],stage4_20[5],stage4_19[16],stage4_18[16],stage4_17[22]}
   );
   gpc606_5 gpc3998 (
      {stage3_17[28], stage3_17[29], stage3_17[30], stage3_17[31], stage3_17[32], stage3_17[33]},
      {stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11], stage3_19[12], stage3_19[13]},
      {stage4_21[3],stage4_20[6],stage4_19[17],stage4_18[17],stage4_17[23]}
   );
   gpc606_5 gpc3999 (
      {stage3_17[34], stage3_17[35], stage3_17[36], stage3_17[37], stage3_17[38], stage3_17[39]},
      {stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17], stage3_19[18], stage3_19[19]},
      {stage4_21[4],stage4_20[7],stage4_19[18],stage4_18[18],stage4_17[24]}
   );
   gpc615_5 gpc4000 (
      {stage3_19[20], stage3_19[21], stage3_19[22], stage3_19[23], stage3_19[24]},
      {stage3_20[2]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[5],stage4_20[8],stage4_19[19]}
   );
   gpc615_5 gpc4001 (
      {stage3_19[25], stage3_19[26], stage3_19[27], stage3_19[28], stage3_19[29]},
      {stage3_20[3]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[1],stage4_21[6],stage4_20[9],stage4_19[20]}
   );
   gpc615_5 gpc4002 (
      {stage3_19[30], stage3_19[31], stage3_19[32], stage3_19[33], stage3_19[34]},
      {stage3_20[4]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[2],stage4_21[7],stage4_20[10],stage4_19[21]}
   );
   gpc615_5 gpc4003 (
      {stage3_19[35], stage3_19[36], stage3_19[37], stage3_19[38], stage3_19[39]},
      {stage3_20[5]},
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage4_23[3],stage4_22[3],stage4_21[8],stage4_20[11],stage4_19[22]}
   );
   gpc1325_5 gpc4004 (
      {stage3_19[40], stage3_19[41], stage3_19[42], stage3_19[43], stage3_19[44]},
      {stage3_20[6], stage3_20[7]},
      {stage3_21[24], stage3_21[25], stage3_21[26]},
      {stage3_22[0]},
      {stage4_23[4],stage4_22[4],stage4_21[9],stage4_20[12],stage4_19[23]}
   );
   gpc1406_5 gpc4005 (
      {stage3_20[8], stage3_20[9], stage3_20[10], stage3_20[11], stage3_20[12], stage3_20[13]},
      {stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4]},
      {stage3_23[0]},
      {stage4_24[0],stage4_23[5],stage4_22[5],stage4_21[10],stage4_20[13]}
   );
   gpc606_5 gpc4006 (
      {stage3_20[14], stage3_20[15], stage3_20[16], stage3_20[17], stage3_20[18], stage3_20[19]},
      {stage3_22[5], stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10]},
      {stage4_24[1],stage4_23[6],stage4_22[6],stage4_21[11],stage4_20[14]}
   );
   gpc606_5 gpc4007 (
      {stage3_20[20], stage3_20[21], stage3_20[22], stage3_20[23], stage3_20[24], stage3_20[25]},
      {stage3_22[11], stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16]},
      {stage4_24[2],stage4_23[7],stage4_22[7],stage4_21[12],stage4_20[15]}
   );
   gpc606_5 gpc4008 (
      {stage3_20[26], stage3_20[27], stage3_20[28], stage3_20[29], stage3_20[30], stage3_20[31]},
      {stage3_22[17], stage3_22[18], stage3_22[19], stage3_22[20], stage3_22[21], stage3_22[22]},
      {stage4_24[3],stage4_23[8],stage4_22[8],stage4_21[13],stage4_20[16]}
   );
   gpc606_5 gpc4009 (
      {stage3_20[32], stage3_20[33], stage3_20[34], stage3_20[35], stage3_20[36], stage3_20[37]},
      {stage3_22[23], stage3_22[24], stage3_22[25], stage3_22[26], stage3_22[27], stage3_22[28]},
      {stage4_24[4],stage4_23[9],stage4_22[9],stage4_21[14],stage4_20[17]}
   );
   gpc606_5 gpc4010 (
      {stage3_21[27], stage3_21[28], stage3_21[29], stage3_21[30], stage3_21[31], stage3_21[32]},
      {stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5], stage3_23[6]},
      {stage4_25[0],stage4_24[5],stage4_23[10],stage4_22[10],stage4_21[15]}
   );
   gpc606_5 gpc4011 (
      {stage3_21[33], stage3_21[34], stage3_21[35], stage3_21[36], stage3_21[37], stage3_21[38]},
      {stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11], stage3_23[12]},
      {stage4_25[1],stage4_24[6],stage4_23[11],stage4_22[11],stage4_21[16]}
   );
   gpc606_5 gpc4012 (
      {stage3_21[39], stage3_21[40], stage3_21[41], stage3_21[42], stage3_21[43], stage3_21[44]},
      {stage3_23[13], stage3_23[14], stage3_23[15], stage3_23[16], stage3_23[17], stage3_23[18]},
      {stage4_25[2],stage4_24[7],stage4_23[12],stage4_22[12],stage4_21[17]}
   );
   gpc606_5 gpc4013 (
      {stage3_21[45], stage3_21[46], stage3_21[47], stage3_21[48], stage3_21[49], stage3_21[50]},
      {stage3_23[19], stage3_23[20], stage3_23[21], stage3_23[22], stage3_23[23], stage3_23[24]},
      {stage4_25[3],stage4_24[8],stage4_23[13],stage4_22[13],stage4_21[18]}
   );
   gpc606_5 gpc4014 (
      {stage3_21[51], stage3_21[52], stage3_21[53], stage3_21[54], stage3_21[55], stage3_21[56]},
      {stage3_23[25], stage3_23[26], stage3_23[27], stage3_23[28], stage3_23[29], stage3_23[30]},
      {stage4_25[4],stage4_24[9],stage4_23[14],stage4_22[14],stage4_21[19]}
   );
   gpc606_5 gpc4015 (
      {stage3_22[29], stage3_22[30], stage3_22[31], stage3_22[32], stage3_22[33], stage3_22[34]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[5],stage4_24[10],stage4_23[15],stage4_22[15]}
   );
   gpc606_5 gpc4016 (
      {stage3_22[35], stage3_22[36], stage3_22[37], stage3_22[38], stage3_22[39], stage3_22[40]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[6],stage4_24[11],stage4_23[16],stage4_22[16]}
   );
   gpc615_5 gpc4017 (
      {stage3_23[31], stage3_23[32], stage3_23[33], stage3_23[34], stage3_23[35]},
      {stage3_24[12]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[2],stage4_25[7],stage4_24[12],stage4_23[17]}
   );
   gpc615_5 gpc4018 (
      {stage3_23[36], stage3_23[37], stage3_23[38], stage3_23[39], stage3_23[40]},
      {stage3_24[13]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[3],stage4_25[8],stage4_24[13],stage4_23[18]}
   );
   gpc615_5 gpc4019 (
      {stage3_23[41], stage3_23[42], stage3_23[43], stage3_23[44], stage3_23[45]},
      {stage3_24[14]},
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage4_27[2],stage4_26[4],stage4_25[9],stage4_24[14],stage4_23[19]}
   );
   gpc606_5 gpc4020 (
      {stage3_24[15], stage3_24[16], stage3_24[17], stage3_24[18], stage3_24[19], stage3_24[20]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage4_28[0],stage4_27[3],stage4_26[5],stage4_25[10],stage4_24[15]}
   );
   gpc606_5 gpc4021 (
      {stage3_24[21], stage3_24[22], stage3_24[23], stage3_24[24], stage3_24[25], stage3_24[26]},
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage4_28[1],stage4_27[4],stage4_26[6],stage4_25[11],stage4_24[16]}
   );
   gpc606_5 gpc4022 (
      {stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21], stage3_25[22], stage3_25[23]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[2],stage4_27[5],stage4_26[7],stage4_25[12]}
   );
   gpc615_5 gpc4023 (
      {stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27], stage3_25[28]},
      {stage3_26[12]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[3],stage4_27[6],stage4_26[8],stage4_25[13]}
   );
   gpc615_5 gpc4024 (
      {stage3_25[29], stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33]},
      {stage3_26[13]},
      {stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17]},
      {stage4_29[2],stage4_28[4],stage4_27[7],stage4_26[9],stage4_25[14]}
   );
   gpc615_5 gpc4025 (
      {stage3_25[34], stage3_25[35], stage3_25[36], stage3_25[37], stage3_25[38]},
      {stage3_26[14]},
      {stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21], stage3_27[22], stage3_27[23]},
      {stage4_29[3],stage4_28[5],stage4_27[8],stage4_26[10],stage4_25[15]}
   );
   gpc615_5 gpc4026 (
      {stage3_26[15], stage3_26[16], stage3_26[17], stage3_26[18], stage3_26[19]},
      {stage3_27[24]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage4_30[0],stage4_29[4],stage4_28[6],stage4_27[9],stage4_26[11]}
   );
   gpc606_5 gpc4027 (
      {stage3_27[25], stage3_27[26], stage3_27[27], stage3_27[28], stage3_27[29], stage3_27[30]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[1],stage4_29[5],stage4_28[7],stage4_27[10]}
   );
   gpc606_5 gpc4028 (
      {stage3_27[31], stage3_27[32], stage3_27[33], stage3_27[34], stage3_27[35], stage3_27[36]},
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage4_31[1],stage4_30[2],stage4_29[6],stage4_28[8],stage4_27[11]}
   );
   gpc606_5 gpc4029 (
      {stage3_27[37], stage3_27[38], stage3_27[39], stage3_27[40], stage3_27[41], stage3_27[42]},
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage4_31[2],stage4_30[3],stage4_29[7],stage4_28[9],stage4_27[12]}
   );
   gpc606_5 gpc4030 (
      {stage3_27[43], stage3_27[44], stage3_27[45], stage3_27[46], stage3_27[47], stage3_27[48]},
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage4_31[3],stage4_30[4],stage4_29[8],stage4_28[10],stage4_27[13]}
   );
   gpc615_5 gpc4031 (
      {stage3_27[49], stage3_27[50], stage3_27[51], stage3_27[52], stage3_27[53]},
      {stage3_28[6]},
      {stage3_29[24], stage3_29[25], stage3_29[26], stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage4_31[4],stage4_30[5],stage4_29[9],stage4_28[11],stage4_27[14]}
   );
   gpc606_5 gpc4032 (
      {stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11], stage3_28[12]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[5],stage4_30[6],stage4_29[10],stage4_28[12]}
   );
   gpc606_5 gpc4033 (
      {stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], stage3_28[17], stage3_28[18]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[6],stage4_30[7],stage4_29[11],stage4_28[13]}
   );
   gpc606_5 gpc4034 (
      {stage3_28[19], stage3_28[20], stage3_28[21], stage3_28[22], stage3_28[23], stage3_28[24]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage4_32[2],stage4_31[7],stage4_30[8],stage4_29[12],stage4_28[14]}
   );
   gpc606_5 gpc4035 (
      {stage3_28[25], stage3_28[26], stage3_28[27], stage3_28[28], stage3_28[29], stage3_28[30]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage4_32[3],stage4_31[8],stage4_30[9],stage4_29[13],stage4_28[15]}
   );
   gpc606_5 gpc4036 (
      {stage3_28[31], stage3_28[32], stage3_28[33], stage3_28[34], stage3_28[35], stage3_28[36]},
      {stage3_30[24], stage3_30[25], stage3_30[26], stage3_30[27], stage3_30[28], stage3_30[29]},
      {stage4_32[4],stage4_31[9],stage4_30[10],stage4_29[14],stage4_28[16]}
   );
   gpc606_5 gpc4037 (
      {stage3_28[37], stage3_28[38], stage3_28[39], stage3_28[40], stage3_28[41], stage3_28[42]},
      {stage3_30[30], stage3_30[31], stage3_30[32], stage3_30[33], stage3_30[34], stage3_30[35]},
      {stage4_32[5],stage4_31[10],stage4_30[11],stage4_29[15],stage4_28[17]}
   );
   gpc615_5 gpc4038 (
      {stage3_29[30], stage3_29[31], stage3_29[32], stage3_29[33], stage3_29[34]},
      {stage3_30[36]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[6],stage4_31[11],stage4_30[12],stage4_29[16]}
   );
   gpc606_5 gpc4039 (
      {stage3_30[37], stage3_30[38], stage3_30[39], stage3_30[40], stage3_30[41], stage3_30[42]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[1],stage4_32[7],stage4_31[12],stage4_30[13]}
   );
   gpc615_5 gpc4040 (
      {stage3_30[43], stage3_30[44], stage3_30[45], stage3_30[46], stage3_30[47]},
      {stage3_31[6]},
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage4_34[1],stage4_33[2],stage4_32[8],stage4_31[13],stage4_30[14]}
   );
   gpc615_5 gpc4041 (
      {stage3_30[48], stage3_30[49], stage3_30[50], stage3_30[51], stage3_30[52]},
      {stage3_31[7]},
      {stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15], stage3_32[16], stage3_32[17]},
      {stage4_34[2],stage4_33[3],stage4_32[9],stage4_31[14],stage4_30[15]}
   );
   gpc606_5 gpc4042 (
      {stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11], stage3_31[12], stage3_31[13]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[3],stage4_33[4],stage4_32[10],stage4_31[15]}
   );
   gpc606_5 gpc4043 (
      {stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17], stage3_31[18], stage3_31[19]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage4_35[1],stage4_34[4],stage4_33[5],stage4_32[11],stage4_31[16]}
   );
   gpc615_5 gpc4044 (
      {stage3_31[20], stage3_31[21], stage3_31[22], stage3_31[23], stage3_31[24]},
      {stage3_32[18]},
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage4_35[2],stage4_34[5],stage4_33[6],stage4_32[12],stage4_31[17]}
   );
   gpc615_5 gpc4045 (
      {stage3_31[25], stage3_31[26], stage3_31[27], stage3_31[28], stage3_31[29]},
      {stage3_32[19]},
      {stage3_33[18], stage3_33[19], stage3_33[20], stage3_33[21], stage3_33[22], stage3_33[23]},
      {stage4_35[3],stage4_34[6],stage4_33[7],stage4_32[13],stage4_31[18]}
   );
   gpc615_5 gpc4046 (
      {stage3_31[30], stage3_31[31], stage3_31[32], stage3_31[33], stage3_31[34]},
      {stage3_32[20]},
      {stage3_33[24], stage3_33[25], stage3_33[26], stage3_33[27], stage3_33[28], stage3_33[29]},
      {stage4_35[4],stage4_34[7],stage4_33[8],stage4_32[14],stage4_31[19]}
   );
   gpc1325_5 gpc4047 (
      {stage3_31[35], stage3_31[36], stage3_31[37], stage3_31[38], stage3_31[39]},
      {stage3_32[21], stage3_32[22]},
      {stage3_33[30], stage3_33[31], stage3_33[32]},
      {stage3_34[0]},
      {stage4_35[5],stage4_34[8],stage4_33[9],stage4_32[15],stage4_31[20]}
   );
   gpc606_5 gpc4048 (
      {stage3_32[23], stage3_32[24], stage3_32[25], stage3_32[26], stage3_32[27], stage3_32[28]},
      {stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5], stage3_34[6]},
      {stage4_36[0],stage4_35[6],stage4_34[9],stage4_33[10],stage4_32[16]}
   );
   gpc606_5 gpc4049 (
      {stage3_32[29], stage3_32[30], stage3_32[31], stage3_32[32], stage3_32[33], stage3_32[34]},
      {stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11], stage3_34[12]},
      {stage4_36[1],stage4_35[7],stage4_34[10],stage4_33[11],stage4_32[17]}
   );
   gpc606_5 gpc4050 (
      {stage3_33[33], stage3_33[34], stage3_33[35], stage3_33[36], stage3_33[37], stage3_33[38]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[2],stage4_35[8],stage4_34[11],stage4_33[12]}
   );
   gpc2135_5 gpc4051 (
      {stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage3_35[6], stage3_35[7], stage3_35[8]},
      {stage3_36[0]},
      {stage3_37[0], stage3_37[1]},
      {stage4_38[0],stage4_37[1],stage4_36[3],stage4_35[9],stage4_34[12]}
   );
   gpc1_1 gpc4052 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc4053 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc4054 (
      {stage3_1[12]},
      {stage4_1[3]}
   );
   gpc1_1 gpc4055 (
      {stage3_1[13]},
      {stage4_1[4]}
   );
   gpc1_1 gpc4056 (
      {stage3_1[14]},
      {stage4_1[5]}
   );
   gpc1_1 gpc4057 (
      {stage3_1[15]},
      {stage4_1[6]}
   );
   gpc1_1 gpc4058 (
      {stage3_1[16]},
      {stage4_1[7]}
   );
   gpc1_1 gpc4059 (
      {stage3_1[17]},
      {stage4_1[8]}
   );
   gpc1_1 gpc4060 (
      {stage3_2[30]},
      {stage4_2[7]}
   );
   gpc1_1 gpc4061 (
      {stage3_2[31]},
      {stage4_2[8]}
   );
   gpc1_1 gpc4062 (
      {stage3_4[39]},
      {stage4_4[12]}
   );
   gpc1_1 gpc4063 (
      {stage3_4[40]},
      {stage4_4[13]}
   );
   gpc1_1 gpc4064 (
      {stage3_4[41]},
      {stage4_4[14]}
   );
   gpc1_1 gpc4065 (
      {stage3_4[42]},
      {stage4_4[15]}
   );
   gpc1_1 gpc4066 (
      {stage3_4[43]},
      {stage4_4[16]}
   );
   gpc1_1 gpc4067 (
      {stage3_5[42]},
      {stage4_5[16]}
   );
   gpc1_1 gpc4068 (
      {stage3_5[43]},
      {stage4_5[17]}
   );
   gpc1_1 gpc4069 (
      {stage3_5[44]},
      {stage4_5[18]}
   );
   gpc1_1 gpc4070 (
      {stage3_5[45]},
      {stage4_5[19]}
   );
   gpc1_1 gpc4071 (
      {stage3_5[46]},
      {stage4_5[20]}
   );
   gpc1_1 gpc4072 (
      {stage3_5[47]},
      {stage4_5[21]}
   );
   gpc1_1 gpc4073 (
      {stage3_5[48]},
      {stage4_5[22]}
   );
   gpc1_1 gpc4074 (
      {stage3_6[39]},
      {stage4_6[17]}
   );
   gpc1_1 gpc4075 (
      {stage3_6[40]},
      {stage4_6[18]}
   );
   gpc1_1 gpc4076 (
      {stage3_6[41]},
      {stage4_6[19]}
   );
   gpc1_1 gpc4077 (
      {stage3_6[42]},
      {stage4_6[20]}
   );
   gpc1_1 gpc4078 (
      {stage3_7[63]},
      {stage4_7[21]}
   );
   gpc1_1 gpc4079 (
      {stage3_7[64]},
      {stage4_7[22]}
   );
   gpc1_1 gpc4080 (
      {stage3_7[65]},
      {stage4_7[23]}
   );
   gpc1_1 gpc4081 (
      {stage3_7[66]},
      {stage4_7[24]}
   );
   gpc1_1 gpc4082 (
      {stage3_7[67]},
      {stage4_7[25]}
   );
   gpc1_1 gpc4083 (
      {stage3_7[68]},
      {stage4_7[26]}
   );
   gpc1_1 gpc4084 (
      {stage3_8[34]},
      {stage4_8[19]}
   );
   gpc1_1 gpc4085 (
      {stage3_8[35]},
      {stage4_8[20]}
   );
   gpc1_1 gpc4086 (
      {stage3_8[36]},
      {stage4_8[21]}
   );
   gpc1_1 gpc4087 (
      {stage3_8[37]},
      {stage4_8[22]}
   );
   gpc1_1 gpc4088 (
      {stage3_9[66]},
      {stage4_9[23]}
   );
   gpc1_1 gpc4089 (
      {stage3_9[67]},
      {stage4_9[24]}
   );
   gpc1_1 gpc4090 (
      {stage3_9[68]},
      {stage4_9[25]}
   );
   gpc1_1 gpc4091 (
      {stage3_9[69]},
      {stage4_9[26]}
   );
   gpc1_1 gpc4092 (
      {stage3_10[18]},
      {stage4_10[18]}
   );
   gpc1_1 gpc4093 (
      {stage3_10[19]},
      {stage4_10[19]}
   );
   gpc1_1 gpc4094 (
      {stage3_10[20]},
      {stage4_10[20]}
   );
   gpc1_1 gpc4095 (
      {stage3_10[21]},
      {stage4_10[21]}
   );
   gpc1_1 gpc4096 (
      {stage3_10[22]},
      {stage4_10[22]}
   );
   gpc1_1 gpc4097 (
      {stage3_10[23]},
      {stage4_10[23]}
   );
   gpc1_1 gpc4098 (
      {stage3_10[24]},
      {stage4_10[24]}
   );
   gpc1_1 gpc4099 (
      {stage3_10[25]},
      {stage4_10[25]}
   );
   gpc1_1 gpc4100 (
      {stage3_10[26]},
      {stage4_10[26]}
   );
   gpc1_1 gpc4101 (
      {stage3_10[27]},
      {stage4_10[27]}
   );
   gpc1_1 gpc4102 (
      {stage3_10[28]},
      {stage4_10[28]}
   );
   gpc1_1 gpc4103 (
      {stage3_11[39]},
      {stage4_11[16]}
   );
   gpc1_1 gpc4104 (
      {stage3_11[40]},
      {stage4_11[17]}
   );
   gpc1_1 gpc4105 (
      {stage3_11[41]},
      {stage4_11[18]}
   );
   gpc1_1 gpc4106 (
      {stage3_11[42]},
      {stage4_11[19]}
   );
   gpc1_1 gpc4107 (
      {stage3_11[43]},
      {stage4_11[20]}
   );
   gpc1_1 gpc4108 (
      {stage3_13[32]},
      {stage4_13[19]}
   );
   gpc1_1 gpc4109 (
      {stage3_13[33]},
      {stage4_13[20]}
   );
   gpc1_1 gpc4110 (
      {stage3_13[34]},
      {stage4_13[21]}
   );
   gpc1_1 gpc4111 (
      {stage3_13[35]},
      {stage4_13[22]}
   );
   gpc1_1 gpc4112 (
      {stage3_13[36]},
      {stage4_13[23]}
   );
   gpc1_1 gpc4113 (
      {stage3_13[37]},
      {stage4_13[24]}
   );
   gpc1_1 gpc4114 (
      {stage3_13[38]},
      {stage4_13[25]}
   );
   gpc1_1 gpc4115 (
      {stage3_13[39]},
      {stage4_13[26]}
   );
   gpc1_1 gpc4116 (
      {stage3_13[40]},
      {stage4_13[27]}
   );
   gpc1_1 gpc4117 (
      {stage3_15[66]},
      {stage4_15[24]}
   );
   gpc1_1 gpc4118 (
      {stage3_15[67]},
      {stage4_15[25]}
   );
   gpc1_1 gpc4119 (
      {stage3_15[68]},
      {stage4_15[26]}
   );
   gpc1_1 gpc4120 (
      {stage3_15[69]},
      {stage4_15[27]}
   );
   gpc1_1 gpc4121 (
      {stage3_15[70]},
      {stage4_15[28]}
   );
   gpc1_1 gpc4122 (
      {stage3_15[71]},
      {stage4_15[29]}
   );
   gpc1_1 gpc4123 (
      {stage3_15[72]},
      {stage4_15[30]}
   );
   gpc1_1 gpc4124 (
      {stage3_15[73]},
      {stage4_15[31]}
   );
   gpc1_1 gpc4125 (
      {stage3_15[74]},
      {stage4_15[32]}
   );
   gpc1_1 gpc4126 (
      {stage3_15[75]},
      {stage4_15[33]}
   );
   gpc1_1 gpc4127 (
      {stage3_15[76]},
      {stage4_15[34]}
   );
   gpc1_1 gpc4128 (
      {stage3_15[77]},
      {stage4_15[35]}
   );
   gpc1_1 gpc4129 (
      {stage3_15[78]},
      {stage4_15[36]}
   );
   gpc1_1 gpc4130 (
      {stage3_15[79]},
      {stage4_15[37]}
   );
   gpc1_1 gpc4131 (
      {stage3_15[80]},
      {stage4_15[38]}
   );
   gpc1_1 gpc4132 (
      {stage3_15[81]},
      {stage4_15[39]}
   );
   gpc1_1 gpc4133 (
      {stage3_15[82]},
      {stage4_15[40]}
   );
   gpc1_1 gpc4134 (
      {stage3_15[83]},
      {stage4_15[41]}
   );
   gpc1_1 gpc4135 (
      {stage3_15[84]},
      {stage4_15[42]}
   );
   gpc1_1 gpc4136 (
      {stage3_15[85]},
      {stage4_15[43]}
   );
   gpc1_1 gpc4137 (
      {stage3_15[86]},
      {stage4_15[44]}
   );
   gpc1_1 gpc4138 (
      {stage3_15[87]},
      {stage4_15[45]}
   );
   gpc1_1 gpc4139 (
      {stage3_15[88]},
      {stage4_15[46]}
   );
   gpc1_1 gpc4140 (
      {stage3_15[89]},
      {stage4_15[47]}
   );
   gpc1_1 gpc4141 (
      {stage3_16[59]},
      {stage4_16[26]}
   );
   gpc1_1 gpc4142 (
      {stage3_16[60]},
      {stage4_16[27]}
   );
   gpc1_1 gpc4143 (
      {stage3_16[61]},
      {stage4_16[28]}
   );
   gpc1_1 gpc4144 (
      {stage3_17[40]},
      {stage4_17[25]}
   );
   gpc1_1 gpc4145 (
      {stage3_17[41]},
      {stage4_17[26]}
   );
   gpc1_1 gpc4146 (
      {stage3_17[42]},
      {stage4_17[27]}
   );
   gpc1_1 gpc4147 (
      {stage3_17[43]},
      {stage4_17[28]}
   );
   gpc1_1 gpc4148 (
      {stage3_17[44]},
      {stage4_17[29]}
   );
   gpc1_1 gpc4149 (
      {stage3_17[45]},
      {stage4_17[30]}
   );
   gpc1_1 gpc4150 (
      {stage3_17[46]},
      {stage4_17[31]}
   );
   gpc1_1 gpc4151 (
      {stage3_17[47]},
      {stage4_17[32]}
   );
   gpc1_1 gpc4152 (
      {stage3_17[48]},
      {stage4_17[33]}
   );
   gpc1_1 gpc4153 (
      {stage3_17[49]},
      {stage4_17[34]}
   );
   gpc1_1 gpc4154 (
      {stage3_19[45]},
      {stage4_19[24]}
   );
   gpc1_1 gpc4155 (
      {stage3_19[46]},
      {stage4_19[25]}
   );
   gpc1_1 gpc4156 (
      {stage3_19[47]},
      {stage4_19[26]}
   );
   gpc1_1 gpc4157 (
      {stage3_19[48]},
      {stage4_19[27]}
   );
   gpc1_1 gpc4158 (
      {stage3_19[49]},
      {stage4_19[28]}
   );
   gpc1_1 gpc4159 (
      {stage3_20[38]},
      {stage4_20[18]}
   );
   gpc1_1 gpc4160 (
      {stage3_20[39]},
      {stage4_20[19]}
   );
   gpc1_1 gpc4161 (
      {stage3_20[40]},
      {stage4_20[20]}
   );
   gpc1_1 gpc4162 (
      {stage3_20[41]},
      {stage4_20[21]}
   );
   gpc1_1 gpc4163 (
      {stage3_20[42]},
      {stage4_20[22]}
   );
   gpc1_1 gpc4164 (
      {stage3_20[43]},
      {stage4_20[23]}
   );
   gpc1_1 gpc4165 (
      {stage3_20[44]},
      {stage4_20[24]}
   );
   gpc1_1 gpc4166 (
      {stage3_20[45]},
      {stage4_20[25]}
   );
   gpc1_1 gpc4167 (
      {stage3_21[57]},
      {stage4_21[20]}
   );
   gpc1_1 gpc4168 (
      {stage3_21[58]},
      {stage4_21[21]}
   );
   gpc1_1 gpc4169 (
      {stage3_22[41]},
      {stage4_22[17]}
   );
   gpc1_1 gpc4170 (
      {stage3_22[42]},
      {stage4_22[18]}
   );
   gpc1_1 gpc4171 (
      {stage3_22[43]},
      {stage4_22[19]}
   );
   gpc1_1 gpc4172 (
      {stage3_22[44]},
      {stage4_22[20]}
   );
   gpc1_1 gpc4173 (
      {stage3_22[45]},
      {stage4_22[21]}
   );
   gpc1_1 gpc4174 (
      {stage3_22[46]},
      {stage4_22[22]}
   );
   gpc1_1 gpc4175 (
      {stage3_23[46]},
      {stage4_23[20]}
   );
   gpc1_1 gpc4176 (
      {stage3_23[47]},
      {stage4_23[21]}
   );
   gpc1_1 gpc4177 (
      {stage3_24[27]},
      {stage4_24[17]}
   );
   gpc1_1 gpc4178 (
      {stage3_24[28]},
      {stage4_24[18]}
   );
   gpc1_1 gpc4179 (
      {stage3_24[29]},
      {stage4_24[19]}
   );
   gpc1_1 gpc4180 (
      {stage3_24[30]},
      {stage4_24[20]}
   );
   gpc1_1 gpc4181 (
      {stage3_24[31]},
      {stage4_24[21]}
   );
   gpc1_1 gpc4182 (
      {stage3_24[32]},
      {stage4_24[22]}
   );
   gpc1_1 gpc4183 (
      {stage3_24[33]},
      {stage4_24[23]}
   );
   gpc1_1 gpc4184 (
      {stage3_24[34]},
      {stage4_24[24]}
   );
   gpc1_1 gpc4185 (
      {stage3_24[35]},
      {stage4_24[25]}
   );
   gpc1_1 gpc4186 (
      {stage3_24[36]},
      {stage4_24[26]}
   );
   gpc1_1 gpc4187 (
      {stage3_24[37]},
      {stage4_24[27]}
   );
   gpc1_1 gpc4188 (
      {stage3_24[38]},
      {stage4_24[28]}
   );
   gpc1_1 gpc4189 (
      {stage3_24[39]},
      {stage4_24[29]}
   );
   gpc1_1 gpc4190 (
      {stage3_24[40]},
      {stage4_24[30]}
   );
   gpc1_1 gpc4191 (
      {stage3_25[39]},
      {stage4_25[16]}
   );
   gpc1_1 gpc4192 (
      {stage3_26[20]},
      {stage4_26[12]}
   );
   gpc1_1 gpc4193 (
      {stage3_26[21]},
      {stage4_26[13]}
   );
   gpc1_1 gpc4194 (
      {stage3_26[22]},
      {stage4_26[14]}
   );
   gpc1_1 gpc4195 (
      {stage3_26[23]},
      {stage4_26[15]}
   );
   gpc1_1 gpc4196 (
      {stage3_26[24]},
      {stage4_26[16]}
   );
   gpc1_1 gpc4197 (
      {stage3_26[25]},
      {stage4_26[17]}
   );
   gpc1_1 gpc4198 (
      {stage3_26[26]},
      {stage4_26[18]}
   );
   gpc1_1 gpc4199 (
      {stage3_26[27]},
      {stage4_26[19]}
   );
   gpc1_1 gpc4200 (
      {stage3_26[28]},
      {stage4_26[20]}
   );
   gpc1_1 gpc4201 (
      {stage3_26[29]},
      {stage4_26[21]}
   );
   gpc1_1 gpc4202 (
      {stage3_26[30]},
      {stage4_26[22]}
   );
   gpc1_1 gpc4203 (
      {stage3_26[31]},
      {stage4_26[23]}
   );
   gpc1_1 gpc4204 (
      {stage3_27[54]},
      {stage4_27[15]}
   );
   gpc1_1 gpc4205 (
      {stage3_27[55]},
      {stage4_27[16]}
   );
   gpc1_1 gpc4206 (
      {stage3_27[56]},
      {stage4_27[17]}
   );
   gpc1_1 gpc4207 (
      {stage3_27[57]},
      {stage4_27[18]}
   );
   gpc1_1 gpc4208 (
      {stage3_27[58]},
      {stage4_27[19]}
   );
   gpc1_1 gpc4209 (
      {stage3_27[59]},
      {stage4_27[20]}
   );
   gpc1_1 gpc4210 (
      {stage3_27[60]},
      {stage4_27[21]}
   );
   gpc1_1 gpc4211 (
      {stage3_27[61]},
      {stage4_27[22]}
   );
   gpc1_1 gpc4212 (
      {stage3_27[62]},
      {stage4_27[23]}
   );
   gpc1_1 gpc4213 (
      {stage3_27[63]},
      {stage4_27[24]}
   );
   gpc1_1 gpc4214 (
      {stage3_27[64]},
      {stage4_27[25]}
   );
   gpc1_1 gpc4215 (
      {stage3_27[65]},
      {stage4_27[26]}
   );
   gpc1_1 gpc4216 (
      {stage3_27[66]},
      {stage4_27[27]}
   );
   gpc1_1 gpc4217 (
      {stage3_29[35]},
      {stage4_29[17]}
   );
   gpc1_1 gpc4218 (
      {stage3_29[36]},
      {stage4_29[18]}
   );
   gpc1_1 gpc4219 (
      {stage3_29[37]},
      {stage4_29[19]}
   );
   gpc1_1 gpc4220 (
      {stage3_29[38]},
      {stage4_29[20]}
   );
   gpc1_1 gpc4221 (
      {stage3_30[53]},
      {stage4_30[16]}
   );
   gpc1_1 gpc4222 (
      {stage3_30[54]},
      {stage4_30[17]}
   );
   gpc1_1 gpc4223 (
      {stage3_30[55]},
      {stage4_30[18]}
   );
   gpc1_1 gpc4224 (
      {stage3_30[56]},
      {stage4_30[19]}
   );
   gpc1_1 gpc4225 (
      {stage3_30[57]},
      {stage4_30[20]}
   );
   gpc1_1 gpc4226 (
      {stage3_30[58]},
      {stage4_30[21]}
   );
   gpc1_1 gpc4227 (
      {stage3_30[59]},
      {stage4_30[22]}
   );
   gpc1_1 gpc4228 (
      {stage3_32[35]},
      {stage4_32[18]}
   );
   gpc1_1 gpc4229 (
      {stage3_33[39]},
      {stage4_33[13]}
   );
   gpc1_1 gpc4230 (
      {stage3_34[18]},
      {stage4_34[13]}
   );
   gpc1_1 gpc4231 (
      {stage3_34[19]},
      {stage4_34[14]}
   );
   gpc1_1 gpc4232 (
      {stage3_34[20]},
      {stage4_34[15]}
   );
   gpc1_1 gpc4233 (
      {stage3_34[21]},
      {stage4_34[16]}
   );
   gpc1_1 gpc4234 (
      {stage3_35[9]},
      {stage4_35[10]}
   );
   gpc1_1 gpc4235 (
      {stage3_35[10]},
      {stage4_35[11]}
   );
   gpc1_1 gpc4236 (
      {stage3_35[11]},
      {stage4_35[12]}
   );
   gpc1_1 gpc4237 (
      {stage3_35[12]},
      {stage4_35[13]}
   );
   gpc1_1 gpc4238 (
      {stage3_36[1]},
      {stage4_36[4]}
   );
   gpc1_1 gpc4239 (
      {stage3_36[2]},
      {stage4_36[5]}
   );
   gpc1_1 gpc4240 (
      {stage3_36[3]},
      {stage4_36[6]}
   );
   gpc1_1 gpc4241 (
      {stage3_36[4]},
      {stage4_36[7]}
   );
   gpc1_1 gpc4242 (
      {stage3_36[5]},
      {stage4_36[8]}
   );
   gpc1_1 gpc4243 (
      {stage3_36[6]},
      {stage4_36[9]}
   );
   gpc615_5 gpc4244 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4]},
      {stage4_3[0]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc1343_5 gpc4245 (
      {stage4_3[1], stage4_3[2], stage4_3[3]},
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9]},
      {stage4_5[0], stage4_5[1], stage4_5[2]},
      {stage4_6[0]},
      {stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[1],stage5_3[1]}
   );
   gpc606_5 gpc4246 (
      {stage4_4[10], stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15]},
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5], stage4_6[6]},
      {stage5_8[0],stage5_7[1],stage5_6[2],stage5_5[2],stage5_4[2]}
   );
   gpc1415_5 gpc4247 (
      {stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6], stage4_5[7]},
      {stage4_6[7]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3]},
      {stage4_8[0]},
      {stage5_9[0],stage5_8[1],stage5_7[2],stage5_6[3],stage5_5[3]}
   );
   gpc606_5 gpc4248 (
      {stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11], stage4_5[12], stage4_5[13]},
      {stage4_7[4], stage4_7[5], stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9]},
      {stage5_9[1],stage5_8[2],stage5_7[3],stage5_6[4],stage5_5[4]}
   );
   gpc606_5 gpc4249 (
      {stage4_5[14], stage4_5[15], stage4_5[16], stage4_5[17], stage4_5[18], stage4_5[19]},
      {stage4_7[10], stage4_7[11], stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15]},
      {stage5_9[2],stage5_8[3],stage5_7[4],stage5_6[5],stage5_5[5]}
   );
   gpc606_5 gpc4250 (
      {stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11], stage4_6[12], stage4_6[13]},
      {stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5], stage4_8[6]},
      {stage5_10[0],stage5_9[3],stage5_8[4],stage5_7[5],stage5_6[6]}
   );
   gpc615_5 gpc4251 (
      {stage4_6[14], stage4_6[15], stage4_6[16], stage4_6[17], stage4_6[18]},
      {stage4_7[16]},
      {stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11], stage4_8[12]},
      {stage5_10[1],stage5_9[4],stage5_8[5],stage5_7[6],stage5_6[7]}
   );
   gpc1343_5 gpc4252 (
      {stage4_7[17], stage4_7[18], stage4_7[19]},
      {stage4_8[13], stage4_8[14], stage4_8[15], stage4_8[16]},
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[2],stage5_9[5],stage5_8[6],stage5_7[7]}
   );
   gpc615_5 gpc4253 (
      {stage4_7[20], stage4_7[21], stage4_7[22], stage4_7[23], stage4_7[24]},
      {stage4_8[17]},
      {stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6], stage4_9[7], stage4_9[8]},
      {stage5_11[1],stage5_10[3],stage5_9[6],stage5_8[7],stage5_7[8]}
   );
   gpc606_5 gpc4254 (
      {stage4_9[9], stage4_9[10], stage4_9[11], stage4_9[12], stage4_9[13], stage4_9[14]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[0],stage5_11[2],stage5_10[4],stage5_9[7]}
   );
   gpc615_5 gpc4255 (
      {stage4_9[15], stage4_9[16], stage4_9[17], stage4_9[18], stage4_9[19]},
      {stage4_10[1]},
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage5_13[1],stage5_12[1],stage5_11[3],stage5_10[5],stage5_9[8]}
   );
   gpc615_5 gpc4256 (
      {stage4_9[20], stage4_9[21], stage4_9[22], stage4_9[23], stage4_9[24]},
      {stage4_10[2]},
      {stage4_11[12], stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17]},
      {stage5_13[2],stage5_12[2],stage5_11[4],stage5_10[6],stage5_9[9]}
   );
   gpc207_4 gpc4257 (
      {stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[3],stage5_12[3],stage5_11[5],stage5_10[7]}
   );
   gpc615_5 gpc4258 (
      {stage4_10[10], stage4_10[11], stage4_10[12], stage4_10[13], stage4_10[14]},
      {stage4_11[18]},
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7]},
      {stage5_14[0],stage5_13[4],stage5_12[4],stage5_11[6],stage5_10[8]}
   );
   gpc1163_5 gpc4259 (
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage4_15[0]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[1],stage5_13[5]}
   );
   gpc606_5 gpc4260 (
      {stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6], stage4_13[7], stage4_13[8]},
      {stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5], stage4_15[6]},
      {stage5_17[1],stage5_16[1],stage5_15[1],stage5_14[2],stage5_13[6]}
   );
   gpc606_5 gpc4261 (
      {stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12], stage4_13[13], stage4_13[14]},
      {stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11], stage4_15[12]},
      {stage5_17[2],stage5_16[2],stage5_15[2],stage5_14[3],stage5_13[7]}
   );
   gpc606_5 gpc4262 (
      {stage4_13[15], stage4_13[16], stage4_13[17], stage4_13[18], stage4_13[19], stage4_13[20]},
      {stage4_15[13], stage4_15[14], stage4_15[15], stage4_15[16], stage4_15[17], stage4_15[18]},
      {stage5_17[3],stage5_16[3],stage5_15[3],stage5_14[4],stage5_13[8]}
   );
   gpc615_5 gpc4263 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[19]},
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5], stage4_16[6]},
      {stage5_18[0],stage5_17[4],stage5_16[4],stage5_15[4],stage5_14[5]}
   );
   gpc207_4 gpc4264 (
      {stage4_15[20], stage4_15[21], stage4_15[22], stage4_15[23], stage4_15[24], stage4_15[25], stage4_15[26]},
      {stage4_17[0], stage4_17[1]},
      {stage5_18[1],stage5_17[5],stage5_16[5],stage5_15[5]}
   );
   gpc615_5 gpc4265 (
      {stage4_15[27], stage4_15[28], stage4_15[29], stage4_15[30], stage4_15[31]},
      {stage4_16[7]},
      {stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5], stage4_17[6], stage4_17[7]},
      {stage5_19[0],stage5_18[2],stage5_17[6],stage5_16[6],stage5_15[6]}
   );
   gpc615_5 gpc4266 (
      {stage4_15[32], stage4_15[33], stage4_15[34], stage4_15[35], stage4_15[36]},
      {stage4_16[8]},
      {stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11], stage4_17[12], stage4_17[13]},
      {stage5_19[1],stage5_18[3],stage5_17[7],stage5_16[7],stage5_15[7]}
   );
   gpc615_5 gpc4267 (
      {stage4_15[37], stage4_15[38], stage4_15[39], stage4_15[40], stage4_15[41]},
      {stage4_16[9]},
      {stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17], stage4_17[18], stage4_17[19]},
      {stage5_19[2],stage5_18[4],stage5_17[8],stage5_16[8],stage5_15[8]}
   );
   gpc615_5 gpc4268 (
      {stage4_15[42], stage4_15[43], stage4_15[44], stage4_15[45], stage4_15[46]},
      {stage4_16[10]},
      {stage4_17[20], stage4_17[21], stage4_17[22], stage4_17[23], stage4_17[24], stage4_17[25]},
      {stage5_19[3],stage5_18[5],stage5_17[9],stage5_16[9],stage5_15[9]}
   );
   gpc207_4 gpc4269 (
      {stage4_16[11], stage4_16[12], stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17]},
      {stage4_18[0], stage4_18[1]},
      {stage5_19[4],stage5_18[6],stage5_17[10],stage5_16[10]}
   );
   gpc606_5 gpc4270 (
      {stage4_17[26], stage4_17[27], stage4_17[28], stage4_17[29], stage4_17[30], stage4_17[31]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[0],stage5_19[5],stage5_18[7],stage5_17[11]}
   );
   gpc615_5 gpc4271 (
      {stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6]},
      {stage4_19[6]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[1],stage5_20[1],stage5_19[6],stage5_18[8]}
   );
   gpc615_5 gpc4272 (
      {stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11]},
      {stage4_19[7]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], stage4_20[11]},
      {stage5_22[1],stage5_21[2],stage5_20[2],stage5_19[7],stage5_18[9]}
   );
   gpc615_5 gpc4273 (
      {stage4_18[12], stage4_18[13], stage4_18[14], stage4_18[15], stage4_18[16]},
      {stage4_19[8]},
      {stage4_20[12], stage4_20[13], stage4_20[14], stage4_20[15], stage4_20[16], stage4_20[17]},
      {stage5_22[2],stage5_21[3],stage5_20[3],stage5_19[8],stage5_18[10]}
   );
   gpc2135_5 gpc4274 (
      {stage4_19[9], stage4_19[10], stage4_19[11], stage4_19[12], stage4_19[13]},
      {stage4_20[18], stage4_20[19], stage4_20[20]},
      {stage4_21[0]},
      {stage4_22[0], stage4_22[1]},
      {stage5_23[0],stage5_22[3],stage5_21[4],stage5_20[4],stage5_19[9]}
   );
   gpc615_5 gpc4275 (
      {stage4_19[14], stage4_19[15], stage4_19[16], stage4_19[17], stage4_19[18]},
      {stage4_20[21]},
      {stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5], stage4_21[6]},
      {stage5_23[1],stage5_22[4],stage5_21[5],stage5_20[5],stage5_19[10]}
   );
   gpc615_5 gpc4276 (
      {stage4_19[19], stage4_19[20], stage4_19[21], stage4_19[22], stage4_19[23]},
      {stage4_20[22]},
      {stage4_21[7], stage4_21[8], stage4_21[9], stage4_21[10], stage4_21[11], stage4_21[12]},
      {stage5_23[2],stage5_22[5],stage5_21[6],stage5_20[6],stage5_19[11]}
   );
   gpc615_5 gpc4277 (
      {stage4_19[24], stage4_19[25], stage4_19[26], stage4_19[27], stage4_19[28]},
      {stage4_20[23]},
      {stage4_21[13], stage4_21[14], stage4_21[15], stage4_21[16], stage4_21[17], stage4_21[18]},
      {stage5_23[3],stage5_22[6],stage5_21[7],stage5_20[7],stage5_19[12]}
   );
   gpc615_5 gpc4278 (
      {stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5], stage4_22[6]},
      {stage4_23[0]},
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage5_26[0],stage5_25[0],stage5_24[0],stage5_23[4],stage5_22[7]}
   );
   gpc615_5 gpc4279 (
      {stage4_22[7], stage4_22[8], stage4_22[9], stage4_22[10], stage4_22[11]},
      {stage4_23[1]},
      {stage4_24[6], stage4_24[7], stage4_24[8], stage4_24[9], stage4_24[10], stage4_24[11]},
      {stage5_26[1],stage5_25[1],stage5_24[1],stage5_23[5],stage5_22[8]}
   );
   gpc615_5 gpc4280 (
      {stage4_22[12], stage4_22[13], stage4_22[14], stage4_22[15], stage4_22[16]},
      {stage4_23[2]},
      {stage4_24[12], stage4_24[13], stage4_24[14], stage4_24[15], stage4_24[16], stage4_24[17]},
      {stage5_26[2],stage5_25[2],stage5_24[2],stage5_23[6],stage5_22[9]}
   );
   gpc615_5 gpc4281 (
      {stage4_22[17], stage4_22[18], stage4_22[19], stage4_22[20], stage4_22[21]},
      {stage4_23[3]},
      {stage4_24[18], stage4_24[19], stage4_24[20], stage4_24[21], stage4_24[22], stage4_24[23]},
      {stage5_26[3],stage5_25[3],stage5_24[3],stage5_23[7],stage5_22[10]}
   );
   gpc615_5 gpc4282 (
      {stage4_23[4], stage4_23[5], stage4_23[6], stage4_23[7], stage4_23[8]},
      {stage4_24[24]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[4],stage5_25[4],stage5_24[4],stage5_23[8]}
   );
   gpc615_5 gpc4283 (
      {stage4_23[9], stage4_23[10], stage4_23[11], stage4_23[12], stage4_23[13]},
      {stage4_24[25]},
      {stage4_25[6], stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11]},
      {stage5_27[1],stage5_26[5],stage5_25[5],stage5_24[5],stage5_23[9]}
   );
   gpc615_5 gpc4284 (
      {stage4_23[14], stage4_23[15], stage4_23[16], stage4_23[17], stage4_23[18]},
      {stage4_24[26]},
      {stage4_25[12], stage4_25[13], stage4_25[14], stage4_25[15], stage4_25[16], 1'b0},
      {stage5_27[2],stage5_26[6],stage5_25[6],stage5_24[6],stage5_23[10]}
   );
   gpc606_5 gpc4285 (
      {stage4_24[27], stage4_24[28], stage4_24[29], stage4_24[30], 1'b0, 1'b0},
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5]},
      {stage5_28[0],stage5_27[3],stage5_26[7],stage5_25[7],stage5_24[7]}
   );
   gpc615_5 gpc4286 (
      {stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10]},
      {stage4_27[0]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[4],stage5_26[8]}
   );
   gpc615_5 gpc4287 (
      {stage4_26[11], stage4_26[12], stage4_26[13], stage4_26[14], stage4_26[15]},
      {stage4_27[1]},
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11]},
      {stage5_30[1],stage5_29[1],stage5_28[2],stage5_27[5],stage5_26[9]}
   );
   gpc615_5 gpc4288 (
      {stage4_26[16], stage4_26[17], stage4_26[18], stage4_26[19], stage4_26[20]},
      {stage4_27[2]},
      {stage4_28[12], stage4_28[13], stage4_28[14], stage4_28[15], stage4_28[16], stage4_28[17]},
      {stage5_30[2],stage5_29[2],stage5_28[3],stage5_27[6],stage5_26[10]}
   );
   gpc207_4 gpc4289 (
      {stage4_27[3], stage4_27[4], stage4_27[5], stage4_27[6], stage4_27[7], stage4_27[8], stage4_27[9]},
      {stage4_29[0], stage4_29[1]},
      {stage5_30[3],stage5_29[3],stage5_28[4],stage5_27[7]}
   );
   gpc207_4 gpc4290 (
      {stage4_27[10], stage4_27[11], stage4_27[12], stage4_27[13], stage4_27[14], stage4_27[15], stage4_27[16]},
      {stage4_29[2], stage4_29[3]},
      {stage5_30[4],stage5_29[4],stage5_28[5],stage5_27[8]}
   );
   gpc207_4 gpc4291 (
      {stage4_27[17], stage4_27[18], stage4_27[19], stage4_27[20], stage4_27[21], stage4_27[22], stage4_27[23]},
      {stage4_29[4], stage4_29[5]},
      {stage5_30[5],stage5_29[5],stage5_28[6],stage5_27[9]}
   );
   gpc615_5 gpc4292 (
      {stage4_29[6], stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10]},
      {stage4_30[0]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[6],stage5_29[6]}
   );
   gpc615_5 gpc4293 (
      {stage4_29[11], stage4_29[12], stage4_29[13], stage4_29[14], stage4_29[15]},
      {stage4_30[1]},
      {stage4_31[6], stage4_31[7], stage4_31[8], stage4_31[9], stage4_31[10], stage4_31[11]},
      {stage5_33[1],stage5_32[1],stage5_31[1],stage5_30[7],stage5_29[7]}
   );
   gpc117_4 gpc4294 (
      {stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5], stage4_30[6], stage4_30[7], stage4_30[8]},
      {stage4_31[12]},
      {stage4_32[0]},
      {stage5_33[2],stage5_32[2],stage5_31[2],stage5_30[8]}
   );
   gpc117_4 gpc4295 (
      {stage4_30[9], stage4_30[10], stage4_30[11], stage4_30[12], stage4_30[13], stage4_30[14], stage4_30[15]},
      {stage4_31[13]},
      {stage4_32[1]},
      {stage5_33[3],stage5_32[3],stage5_31[3],stage5_30[9]}
   );
   gpc615_5 gpc4296 (
      {stage4_30[16], stage4_30[17], stage4_30[18], stage4_30[19], stage4_30[20]},
      {stage4_31[14]},
      {stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5], stage4_32[6], stage4_32[7]},
      {stage5_34[0],stage5_33[4],stage5_32[4],stage5_31[4],stage5_30[10]}
   );
   gpc615_5 gpc4297 (
      {stage4_30[21], stage4_30[22], 1'b0, 1'b0, 1'b0},
      {stage4_31[15]},
      {stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11], stage4_32[12], stage4_32[13]},
      {stage5_34[1],stage5_33[5],stage5_32[5],stage5_31[5],stage5_30[11]}
   );
   gpc2135_5 gpc4298 (
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4]},
      {stage4_34[0], stage4_34[1], stage4_34[2]},
      {stage4_35[0]},
      {stage4_36[0], stage4_36[1]},
      {stage5_37[0],stage5_36[0],stage5_35[0],stage5_34[2],stage5_33[6]}
   );
   gpc2135_5 gpc4299 (
      {stage4_33[5], stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9]},
      {stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage4_35[1]},
      {stage4_36[2], stage4_36[3]},
      {stage5_37[1],stage5_36[1],stage5_35[1],stage5_34[3],stage5_33[7]}
   );
   gpc2135_5 gpc4300 (
      {stage4_33[10], stage4_33[11], stage4_33[12], stage4_33[13], 1'b0},
      {stage4_34[6], stage4_34[7], stage4_34[8]},
      {stage4_35[2]},
      {stage4_36[4], stage4_36[5]},
      {stage5_37[2],stage5_36[2],stage5_35[2],stage5_34[4],stage5_33[8]}
   );
   gpc606_5 gpc4301 (
      {stage4_34[9], stage4_34[10], stage4_34[11], stage4_34[12], stage4_34[13], stage4_34[14]},
      {stage4_36[6], stage4_36[7], stage4_36[8], stage4_36[9], 1'b0, 1'b0},
      {stage5_38[0],stage5_37[3],stage5_36[3],stage5_35[3],stage5_34[5]}
   );
   gpc1_1 gpc4302 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc4303 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc4304 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc4305 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc4306 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc4307 (
      {stage4_1[2]},
      {stage5_1[2]}
   );
   gpc1_1 gpc4308 (
      {stage4_1[3]},
      {stage5_1[3]}
   );
   gpc1_1 gpc4309 (
      {stage4_1[4]},
      {stage5_1[4]}
   );
   gpc1_1 gpc4310 (
      {stage4_1[5]},
      {stage5_1[5]}
   );
   gpc1_1 gpc4311 (
      {stage4_1[6]},
      {stage5_1[6]}
   );
   gpc1_1 gpc4312 (
      {stage4_1[7]},
      {stage5_1[7]}
   );
   gpc1_1 gpc4313 (
      {stage4_1[8]},
      {stage5_1[8]}
   );
   gpc1_1 gpc4314 (
      {stage4_2[5]},
      {stage5_2[1]}
   );
   gpc1_1 gpc4315 (
      {stage4_2[6]},
      {stage5_2[2]}
   );
   gpc1_1 gpc4316 (
      {stage4_2[7]},
      {stage5_2[3]}
   );
   gpc1_1 gpc4317 (
      {stage4_2[8]},
      {stage5_2[4]}
   );
   gpc1_1 gpc4318 (
      {stage4_3[4]},
      {stage5_3[2]}
   );
   gpc1_1 gpc4319 (
      {stage4_3[5]},
      {stage5_3[3]}
   );
   gpc1_1 gpc4320 (
      {stage4_3[6]},
      {stage5_3[4]}
   );
   gpc1_1 gpc4321 (
      {stage4_3[7]},
      {stage5_3[5]}
   );
   gpc1_1 gpc4322 (
      {stage4_3[8]},
      {stage5_3[6]}
   );
   gpc1_1 gpc4323 (
      {stage4_3[9]},
      {stage5_3[7]}
   );
   gpc1_1 gpc4324 (
      {stage4_4[16]},
      {stage5_4[3]}
   );
   gpc1_1 gpc4325 (
      {stage4_5[20]},
      {stage5_5[6]}
   );
   gpc1_1 gpc4326 (
      {stage4_5[21]},
      {stage5_5[7]}
   );
   gpc1_1 gpc4327 (
      {stage4_5[22]},
      {stage5_5[8]}
   );
   gpc1_1 gpc4328 (
      {stage4_6[19]},
      {stage5_6[8]}
   );
   gpc1_1 gpc4329 (
      {stage4_6[20]},
      {stage5_6[9]}
   );
   gpc1_1 gpc4330 (
      {stage4_7[25]},
      {stage5_7[9]}
   );
   gpc1_1 gpc4331 (
      {stage4_7[26]},
      {stage5_7[10]}
   );
   gpc1_1 gpc4332 (
      {stage4_8[18]},
      {stage5_8[8]}
   );
   gpc1_1 gpc4333 (
      {stage4_8[19]},
      {stage5_8[9]}
   );
   gpc1_1 gpc4334 (
      {stage4_8[20]},
      {stage5_8[10]}
   );
   gpc1_1 gpc4335 (
      {stage4_8[21]},
      {stage5_8[11]}
   );
   gpc1_1 gpc4336 (
      {stage4_8[22]},
      {stage5_8[12]}
   );
   gpc1_1 gpc4337 (
      {stage4_9[25]},
      {stage5_9[10]}
   );
   gpc1_1 gpc4338 (
      {stage4_9[26]},
      {stage5_9[11]}
   );
   gpc1_1 gpc4339 (
      {stage4_10[15]},
      {stage5_10[9]}
   );
   gpc1_1 gpc4340 (
      {stage4_10[16]},
      {stage5_10[10]}
   );
   gpc1_1 gpc4341 (
      {stage4_10[17]},
      {stage5_10[11]}
   );
   gpc1_1 gpc4342 (
      {stage4_10[18]},
      {stage5_10[12]}
   );
   gpc1_1 gpc4343 (
      {stage4_10[19]},
      {stage5_10[13]}
   );
   gpc1_1 gpc4344 (
      {stage4_10[20]},
      {stage5_10[14]}
   );
   gpc1_1 gpc4345 (
      {stage4_10[21]},
      {stage5_10[15]}
   );
   gpc1_1 gpc4346 (
      {stage4_10[22]},
      {stage5_10[16]}
   );
   gpc1_1 gpc4347 (
      {stage4_10[23]},
      {stage5_10[17]}
   );
   gpc1_1 gpc4348 (
      {stage4_10[24]},
      {stage5_10[18]}
   );
   gpc1_1 gpc4349 (
      {stage4_10[25]},
      {stage5_10[19]}
   );
   gpc1_1 gpc4350 (
      {stage4_10[26]},
      {stage5_10[20]}
   );
   gpc1_1 gpc4351 (
      {stage4_10[27]},
      {stage5_10[21]}
   );
   gpc1_1 gpc4352 (
      {stage4_10[28]},
      {stage5_10[22]}
   );
   gpc1_1 gpc4353 (
      {stage4_11[19]},
      {stage5_11[7]}
   );
   gpc1_1 gpc4354 (
      {stage4_11[20]},
      {stage5_11[8]}
   );
   gpc1_1 gpc4355 (
      {stage4_12[8]},
      {stage5_12[5]}
   );
   gpc1_1 gpc4356 (
      {stage4_12[9]},
      {stage5_12[6]}
   );
   gpc1_1 gpc4357 (
      {stage4_12[10]},
      {stage5_12[7]}
   );
   gpc1_1 gpc4358 (
      {stage4_12[11]},
      {stage5_12[8]}
   );
   gpc1_1 gpc4359 (
      {stage4_12[12]},
      {stage5_12[9]}
   );
   gpc1_1 gpc4360 (
      {stage4_12[13]},
      {stage5_12[10]}
   );
   gpc1_1 gpc4361 (
      {stage4_13[21]},
      {stage5_13[9]}
   );
   gpc1_1 gpc4362 (
      {stage4_13[22]},
      {stage5_13[10]}
   );
   gpc1_1 gpc4363 (
      {stage4_13[23]},
      {stage5_13[11]}
   );
   gpc1_1 gpc4364 (
      {stage4_13[24]},
      {stage5_13[12]}
   );
   gpc1_1 gpc4365 (
      {stage4_13[25]},
      {stage5_13[13]}
   );
   gpc1_1 gpc4366 (
      {stage4_13[26]},
      {stage5_13[14]}
   );
   gpc1_1 gpc4367 (
      {stage4_13[27]},
      {stage5_13[15]}
   );
   gpc1_1 gpc4368 (
      {stage4_14[11]},
      {stage5_14[6]}
   );
   gpc1_1 gpc4369 (
      {stage4_14[12]},
      {stage5_14[7]}
   );
   gpc1_1 gpc4370 (
      {stage4_15[47]},
      {stage5_15[10]}
   );
   gpc1_1 gpc4371 (
      {stage4_16[18]},
      {stage5_16[11]}
   );
   gpc1_1 gpc4372 (
      {stage4_16[19]},
      {stage5_16[12]}
   );
   gpc1_1 gpc4373 (
      {stage4_16[20]},
      {stage5_16[13]}
   );
   gpc1_1 gpc4374 (
      {stage4_16[21]},
      {stage5_16[14]}
   );
   gpc1_1 gpc4375 (
      {stage4_16[22]},
      {stage5_16[15]}
   );
   gpc1_1 gpc4376 (
      {stage4_16[23]},
      {stage5_16[16]}
   );
   gpc1_1 gpc4377 (
      {stage4_16[24]},
      {stage5_16[17]}
   );
   gpc1_1 gpc4378 (
      {stage4_16[25]},
      {stage5_16[18]}
   );
   gpc1_1 gpc4379 (
      {stage4_16[26]},
      {stage5_16[19]}
   );
   gpc1_1 gpc4380 (
      {stage4_16[27]},
      {stage5_16[20]}
   );
   gpc1_1 gpc4381 (
      {stage4_16[28]},
      {stage5_16[21]}
   );
   gpc1_1 gpc4382 (
      {stage4_17[32]},
      {stage5_17[12]}
   );
   gpc1_1 gpc4383 (
      {stage4_17[33]},
      {stage5_17[13]}
   );
   gpc1_1 gpc4384 (
      {stage4_17[34]},
      {stage5_17[14]}
   );
   gpc1_1 gpc4385 (
      {stage4_18[17]},
      {stage5_18[11]}
   );
   gpc1_1 gpc4386 (
      {stage4_18[18]},
      {stage5_18[12]}
   );
   gpc1_1 gpc4387 (
      {stage4_20[24]},
      {stage5_20[8]}
   );
   gpc1_1 gpc4388 (
      {stage4_20[25]},
      {stage5_20[9]}
   );
   gpc1_1 gpc4389 (
      {stage4_21[19]},
      {stage5_21[8]}
   );
   gpc1_1 gpc4390 (
      {stage4_21[20]},
      {stage5_21[9]}
   );
   gpc1_1 gpc4391 (
      {stage4_21[21]},
      {stage5_21[10]}
   );
   gpc1_1 gpc4392 (
      {stage4_22[22]},
      {stage5_22[11]}
   );
   gpc1_1 gpc4393 (
      {stage4_23[19]},
      {stage5_23[11]}
   );
   gpc1_1 gpc4394 (
      {stage4_23[20]},
      {stage5_23[12]}
   );
   gpc1_1 gpc4395 (
      {stage4_23[21]},
      {stage5_23[13]}
   );
   gpc1_1 gpc4396 (
      {stage4_26[21]},
      {stage5_26[11]}
   );
   gpc1_1 gpc4397 (
      {stage4_26[22]},
      {stage5_26[12]}
   );
   gpc1_1 gpc4398 (
      {stage4_26[23]},
      {stage5_26[13]}
   );
   gpc1_1 gpc4399 (
      {stage4_27[24]},
      {stage5_27[10]}
   );
   gpc1_1 gpc4400 (
      {stage4_27[25]},
      {stage5_27[11]}
   );
   gpc1_1 gpc4401 (
      {stage4_27[26]},
      {stage5_27[12]}
   );
   gpc1_1 gpc4402 (
      {stage4_27[27]},
      {stage5_27[13]}
   );
   gpc1_1 gpc4403 (
      {stage4_29[16]},
      {stage5_29[8]}
   );
   gpc1_1 gpc4404 (
      {stage4_29[17]},
      {stage5_29[9]}
   );
   gpc1_1 gpc4405 (
      {stage4_29[18]},
      {stage5_29[10]}
   );
   gpc1_1 gpc4406 (
      {stage4_29[19]},
      {stage5_29[11]}
   );
   gpc1_1 gpc4407 (
      {stage4_29[20]},
      {stage5_29[12]}
   );
   gpc1_1 gpc4408 (
      {stage4_31[16]},
      {stage5_31[6]}
   );
   gpc1_1 gpc4409 (
      {stage4_31[17]},
      {stage5_31[7]}
   );
   gpc1_1 gpc4410 (
      {stage4_31[18]},
      {stage5_31[8]}
   );
   gpc1_1 gpc4411 (
      {stage4_31[19]},
      {stage5_31[9]}
   );
   gpc1_1 gpc4412 (
      {stage4_31[20]},
      {stage5_31[10]}
   );
   gpc1_1 gpc4413 (
      {stage4_32[14]},
      {stage5_32[6]}
   );
   gpc1_1 gpc4414 (
      {stage4_32[15]},
      {stage5_32[7]}
   );
   gpc1_1 gpc4415 (
      {stage4_32[16]},
      {stage5_32[8]}
   );
   gpc1_1 gpc4416 (
      {stage4_32[17]},
      {stage5_32[9]}
   );
   gpc1_1 gpc4417 (
      {stage4_32[18]},
      {stage5_32[10]}
   );
   gpc1_1 gpc4418 (
      {stage4_34[15]},
      {stage5_34[6]}
   );
   gpc1_1 gpc4419 (
      {stage4_34[16]},
      {stage5_34[7]}
   );
   gpc1_1 gpc4420 (
      {stage4_35[3]},
      {stage5_35[4]}
   );
   gpc1_1 gpc4421 (
      {stage4_35[4]},
      {stage5_35[5]}
   );
   gpc1_1 gpc4422 (
      {stage4_35[5]},
      {stage5_35[6]}
   );
   gpc1_1 gpc4423 (
      {stage4_35[6]},
      {stage5_35[7]}
   );
   gpc1_1 gpc4424 (
      {stage4_35[7]},
      {stage5_35[8]}
   );
   gpc1_1 gpc4425 (
      {stage4_35[8]},
      {stage5_35[9]}
   );
   gpc1_1 gpc4426 (
      {stage4_35[9]},
      {stage5_35[10]}
   );
   gpc1_1 gpc4427 (
      {stage4_35[10]},
      {stage5_35[11]}
   );
   gpc1_1 gpc4428 (
      {stage4_35[11]},
      {stage5_35[12]}
   );
   gpc1_1 gpc4429 (
      {stage4_35[12]},
      {stage5_35[13]}
   );
   gpc1_1 gpc4430 (
      {stage4_35[13]},
      {stage5_35[14]}
   );
   gpc1_1 gpc4431 (
      {stage4_37[0]},
      {stage5_37[4]}
   );
   gpc1_1 gpc4432 (
      {stage4_37[1]},
      {stage5_37[5]}
   );
   gpc1_1 gpc4433 (
      {stage4_38[0]},
      {stage5_38[1]}
   );
   gpc1163_5 gpc4434 (
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4], 1'b0},
      {stage5_3[0]},
      {stage5_4[0]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0]}
   );
   gpc135_4 gpc4435 (
      {stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5]},
      {stage5_4[1], stage5_4[2], stage5_4[3]},
      {stage5_5[0]},
      {stage6_6[0],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc1343_5 gpc4436 (
      {stage5_5[1], stage5_5[2], stage5_5[3]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3]},
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0]},
      {stage6_9[0],stage6_8[0],stage6_7[0],stage6_6[1],stage6_5[2]}
   );
   gpc1343_5 gpc4437 (
      {stage5_5[4], stage5_5[5], stage5_5[6]},
      {stage5_6[4], stage5_6[5], stage5_6[6], stage5_6[7]},
      {stage5_7[3], stage5_7[4], stage5_7[5]},
      {stage5_8[1]},
      {stage6_9[1],stage6_8[1],stage6_7[1],stage6_6[2],stage6_5[3]}
   );
   gpc615_5 gpc4438 (
      {stage5_7[6], stage5_7[7], stage5_7[8], stage5_7[9], stage5_7[10]},
      {stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[0],stage6_9[2],stage6_8[2],stage6_7[2]}
   );
   gpc1163_5 gpc4439 (
      {stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage5_9[6], stage5_9[7], stage5_9[8], stage5_9[9], stage5_9[10], stage5_9[11]},
      {stage5_10[0]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[1],stage6_10[1],stage6_9[3],stage6_8[3]}
   );
   gpc606_5 gpc4440 (
      {stage5_8[6], stage5_8[7], stage5_8[8], stage5_8[9], stage5_8[10], stage5_8[11]},
      {stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5], stage5_10[6]},
      {stage6_12[1],stage6_11[2],stage6_10[2],stage6_9[4],stage6_8[4]}
   );
   gpc117_4 gpc4441 (
      {stage5_10[7], stage5_10[8], stage5_10[9], stage5_10[10], stage5_10[11], stage5_10[12], stage5_10[13]},
      {stage5_11[1]},
      {stage5_12[0]},
      {stage6_13[0],stage6_12[2],stage6_11[3],stage6_10[3]}
   );
   gpc117_4 gpc4442 (
      {stage5_10[14], stage5_10[15], stage5_10[16], stage5_10[17], stage5_10[18], stage5_10[19], stage5_10[20]},
      {stage5_11[2]},
      {stage5_12[1]},
      {stage6_13[1],stage6_12[3],stage6_11[4],stage6_10[4]}
   );
   gpc117_4 gpc4443 (
      {stage5_11[3], stage5_11[4], stage5_11[5], stage5_11[6], stage5_11[7], stage5_11[8], 1'b0},
      {stage5_12[2]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[2],stage6_12[4],stage6_11[5]}
   );
   gpc207_4 gpc4444 (
      {stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6], stage5_12[7], stage5_12[8], stage5_12[9]},
      {stage5_14[0], stage5_14[1]},
      {stage6_15[0],stage6_14[1],stage6_13[3],stage6_12[5]}
   );
   gpc1406_5 gpc4445 (
      {stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5], stage5_13[6]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[1],stage6_14[2],stage6_13[4]}
   );
   gpc1406_5 gpc4446 (
      {stage5_13[7], stage5_13[8], stage5_13[9], stage5_13[10], stage5_13[11], stage5_13[12]},
      {stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7]},
      {stage5_16[1]},
      {stage6_17[1],stage6_16[1],stage6_15[2],stage6_14[3],stage6_13[5]}
   );
   gpc615_5 gpc4447 (
      {stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5], stage5_14[6]},
      {stage5_15[8]},
      {stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5], stage5_16[6], stage5_16[7]},
      {stage6_18[0],stage6_17[2],stage6_16[2],stage6_15[3],stage6_14[4]}
   );
   gpc117_4 gpc4448 (
      {stage5_16[8], stage5_16[9], stage5_16[10], stage5_16[11], stage5_16[12], stage5_16[13], stage5_16[14]},
      {stage5_17[0]},
      {stage5_18[0]},
      {stage6_19[0],stage6_18[1],stage6_17[3],stage6_16[3]}
   );
   gpc7_3 gpc4449 (
      {stage5_16[15], stage5_16[16], stage5_16[17], stage5_16[18], stage5_16[19], stage5_16[20], stage5_16[21]},
      {stage6_18[2],stage6_17[4],stage6_16[4]}
   );
   gpc1163_5 gpc4450 (
      {stage5_17[1], stage5_17[2], stage5_17[3]},
      {stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5], stage5_18[6]},
      {stage5_19[0]},
      {stage5_20[0]},
      {stage6_21[0],stage6_20[0],stage6_19[1],stage6_18[3],stage6_17[5]}
   );
   gpc1163_5 gpc4451 (
      {stage5_17[4], stage5_17[5], stage5_17[6]},
      {stage5_18[7], stage5_18[8], stage5_18[9], stage5_18[10], stage5_18[11], stage5_18[12]},
      {stage5_19[1]},
      {stage5_20[1]},
      {stage6_21[1],stage6_20[1],stage6_19[2],stage6_18[4],stage6_17[6]}
   );
   gpc606_5 gpc4452 (
      {stage5_17[7], stage5_17[8], stage5_17[9], stage5_17[10], stage5_17[11], stage5_17[12]},
      {stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5], stage5_19[6], stage5_19[7]},
      {stage6_21[2],stage6_20[2],stage6_19[3],stage6_18[5],stage6_17[7]}
   );
   gpc615_5 gpc4453 (
      {stage5_19[8], stage5_19[9], stage5_19[10], stage5_19[11], stage5_19[12]},
      {stage5_20[2]},
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage6_23[0],stage6_22[0],stage6_21[3],stage6_20[3],stage6_19[4]}
   );
   gpc606_5 gpc4454 (
      {stage5_20[3], stage5_20[4], stage5_20[5], stage5_20[6], stage5_20[7], stage5_20[8]},
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4], stage5_22[5]},
      {stage6_24[0],stage6_23[1],stage6_22[1],stage6_21[4],stage6_20[4]}
   );
   gpc1406_5 gpc4455 (
      {stage5_21[6], stage5_21[7], stage5_21[8], stage5_21[9], stage5_21[10], 1'b0},
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3]},
      {stage5_24[0]},
      {stage6_25[0],stage6_24[1],stage6_23[2],stage6_22[2],stage6_21[5]}
   );
   gpc615_5 gpc4456 (
      {stage5_22[6], stage5_22[7], stage5_22[8], stage5_22[9], stage5_22[10]},
      {stage5_23[4]},
      {stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], stage5_24[6]},
      {stage6_26[0],stage6_25[1],stage6_24[2],stage6_23[3],stage6_22[3]}
   );
   gpc615_5 gpc4457 (
      {stage5_23[5], stage5_23[6], stage5_23[7], stage5_23[8], stage5_23[9]},
      {stage5_24[7]},
      {stage5_25[0], stage5_25[1], stage5_25[2], stage5_25[3], stage5_25[4], stage5_25[5]},
      {stage6_27[0],stage6_26[1],stage6_25[2],stage6_24[3],stage6_23[4]}
   );
   gpc135_4 gpc4458 (
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4]},
      {stage5_27[0], stage5_27[1], stage5_27[2]},
      {stage5_28[0]},
      {stage6_29[0],stage6_28[0],stage6_27[1],stage6_26[2]}
   );
   gpc615_5 gpc4459 (
      {stage5_27[3], stage5_27[4], stage5_27[5], stage5_27[6], stage5_27[7]},
      {stage5_28[1]},
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage6_31[0],stage6_30[0],stage6_29[1],stage6_28[1],stage6_27[2]}
   );
   gpc606_5 gpc4460 (
      {stage5_29[6], stage5_29[7], stage5_29[8], stage5_29[9], stage5_29[10], stage5_29[11]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[0],stage6_31[1],stage6_30[1],stage6_29[2]}
   );
   gpc1406_5 gpc4461 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5]},
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3]},
      {stage5_33[0]},
      {stage6_34[0],stage6_33[1],stage6_32[1],stage6_31[2],stage6_30[2]}
   );
   gpc615_5 gpc4462 (
      {stage5_30[6], stage5_30[7], stage5_30[8], stage5_30[9], stage5_30[10]},
      {stage5_31[6]},
      {stage5_32[4], stage5_32[5], stage5_32[6], stage5_32[7], stage5_32[8], stage5_32[9]},
      {stage6_34[1],stage6_33[2],stage6_32[2],stage6_31[3],stage6_30[3]}
   );
   gpc606_5 gpc4463 (
      {stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4], stage5_33[5], stage5_33[6]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], stage5_35[4], stage5_35[5]},
      {stage6_37[0],stage6_36[0],stage6_35[0],stage6_34[2],stage6_33[3]}
   );
   gpc606_5 gpc4464 (
      {stage5_35[6], stage5_35[7], stage5_35[8], stage5_35[9], stage5_35[10], stage5_35[11]},
      {stage5_37[0], stage5_37[1], stage5_37[2], stage5_37[3], stage5_37[4], stage5_37[5]},
      {stage6_39[0],stage6_38[0],stage6_37[1],stage6_36[1],stage6_35[1]}
   );
   gpc1_1 gpc4465 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc4466 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc4467 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc4468 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc4469 (
      {stage5_1[4]},
      {stage6_1[2]}
   );
   gpc1_1 gpc4470 (
      {stage5_1[5]},
      {stage6_1[3]}
   );
   gpc1_1 gpc4471 (
      {stage5_1[6]},
      {stage6_1[4]}
   );
   gpc1_1 gpc4472 (
      {stage5_1[7]},
      {stage6_1[5]}
   );
   gpc1_1 gpc4473 (
      {stage5_1[8]},
      {stage6_1[6]}
   );
   gpc1_1 gpc4474 (
      {stage5_3[6]},
      {stage6_3[2]}
   );
   gpc1_1 gpc4475 (
      {stage5_3[7]},
      {stage6_3[3]}
   );
   gpc1_1 gpc4476 (
      {stage5_5[7]},
      {stage6_5[4]}
   );
   gpc1_1 gpc4477 (
      {stage5_5[8]},
      {stage6_5[5]}
   );
   gpc1_1 gpc4478 (
      {stage5_6[8]},
      {stage6_6[3]}
   );
   gpc1_1 gpc4479 (
      {stage5_6[9]},
      {stage6_6[4]}
   );
   gpc1_1 gpc4480 (
      {stage5_8[12]},
      {stage6_8[5]}
   );
   gpc1_1 gpc4481 (
      {stage5_10[21]},
      {stage6_10[5]}
   );
   gpc1_1 gpc4482 (
      {stage5_10[22]},
      {stage6_10[6]}
   );
   gpc1_1 gpc4483 (
      {stage5_12[10]},
      {stage6_12[6]}
   );
   gpc1_1 gpc4484 (
      {stage5_13[13]},
      {stage6_13[6]}
   );
   gpc1_1 gpc4485 (
      {stage5_13[14]},
      {stage6_13[7]}
   );
   gpc1_1 gpc4486 (
      {stage5_13[15]},
      {stage6_13[8]}
   );
   gpc1_1 gpc4487 (
      {stage5_14[7]},
      {stage6_14[5]}
   );
   gpc1_1 gpc4488 (
      {stage5_15[9]},
      {stage6_15[4]}
   );
   gpc1_1 gpc4489 (
      {stage5_15[10]},
      {stage6_15[5]}
   );
   gpc1_1 gpc4490 (
      {stage5_17[13]},
      {stage6_17[8]}
   );
   gpc1_1 gpc4491 (
      {stage5_17[14]},
      {stage6_17[9]}
   );
   gpc1_1 gpc4492 (
      {stage5_20[9]},
      {stage6_20[5]}
   );
   gpc1_1 gpc4493 (
      {stage5_22[11]},
      {stage6_22[4]}
   );
   gpc1_1 gpc4494 (
      {stage5_23[10]},
      {stage6_23[5]}
   );
   gpc1_1 gpc4495 (
      {stage5_23[11]},
      {stage6_23[6]}
   );
   gpc1_1 gpc4496 (
      {stage5_23[12]},
      {stage6_23[7]}
   );
   gpc1_1 gpc4497 (
      {stage5_23[13]},
      {stage6_23[8]}
   );
   gpc1_1 gpc4498 (
      {stage5_25[6]},
      {stage6_25[3]}
   );
   gpc1_1 gpc4499 (
      {stage5_25[7]},
      {stage6_25[4]}
   );
   gpc1_1 gpc4500 (
      {stage5_26[5]},
      {stage6_26[3]}
   );
   gpc1_1 gpc4501 (
      {stage5_26[6]},
      {stage6_26[4]}
   );
   gpc1_1 gpc4502 (
      {stage5_26[7]},
      {stage6_26[5]}
   );
   gpc1_1 gpc4503 (
      {stage5_26[8]},
      {stage6_26[6]}
   );
   gpc1_1 gpc4504 (
      {stage5_26[9]},
      {stage6_26[7]}
   );
   gpc1_1 gpc4505 (
      {stage5_26[10]},
      {stage6_26[8]}
   );
   gpc1_1 gpc4506 (
      {stage5_26[11]},
      {stage6_26[9]}
   );
   gpc1_1 gpc4507 (
      {stage5_26[12]},
      {stage6_26[10]}
   );
   gpc1_1 gpc4508 (
      {stage5_26[13]},
      {stage6_26[11]}
   );
   gpc1_1 gpc4509 (
      {stage5_27[8]},
      {stage6_27[3]}
   );
   gpc1_1 gpc4510 (
      {stage5_27[9]},
      {stage6_27[4]}
   );
   gpc1_1 gpc4511 (
      {stage5_27[10]},
      {stage6_27[5]}
   );
   gpc1_1 gpc4512 (
      {stage5_27[11]},
      {stage6_27[6]}
   );
   gpc1_1 gpc4513 (
      {stage5_27[12]},
      {stage6_27[7]}
   );
   gpc1_1 gpc4514 (
      {stage5_27[13]},
      {stage6_27[8]}
   );
   gpc1_1 gpc4515 (
      {stage5_28[2]},
      {stage6_28[2]}
   );
   gpc1_1 gpc4516 (
      {stage5_28[3]},
      {stage6_28[3]}
   );
   gpc1_1 gpc4517 (
      {stage5_28[4]},
      {stage6_28[4]}
   );
   gpc1_1 gpc4518 (
      {stage5_28[5]},
      {stage6_28[5]}
   );
   gpc1_1 gpc4519 (
      {stage5_28[6]},
      {stage6_28[6]}
   );
   gpc1_1 gpc4520 (
      {stage5_29[12]},
      {stage6_29[3]}
   );
   gpc1_1 gpc4521 (
      {stage5_30[11]},
      {stage6_30[4]}
   );
   gpc1_1 gpc4522 (
      {stage5_31[7]},
      {stage6_31[4]}
   );
   gpc1_1 gpc4523 (
      {stage5_31[8]},
      {stage6_31[5]}
   );
   gpc1_1 gpc4524 (
      {stage5_31[9]},
      {stage6_31[6]}
   );
   gpc1_1 gpc4525 (
      {stage5_31[10]},
      {stage6_31[7]}
   );
   gpc1_1 gpc4526 (
      {stage5_32[10]},
      {stage6_32[3]}
   );
   gpc1_1 gpc4527 (
      {stage5_33[7]},
      {stage6_33[4]}
   );
   gpc1_1 gpc4528 (
      {stage5_33[8]},
      {stage6_33[5]}
   );
   gpc1_1 gpc4529 (
      {stage5_34[0]},
      {stage6_34[3]}
   );
   gpc1_1 gpc4530 (
      {stage5_34[1]},
      {stage6_34[4]}
   );
   gpc1_1 gpc4531 (
      {stage5_34[2]},
      {stage6_34[5]}
   );
   gpc1_1 gpc4532 (
      {stage5_34[3]},
      {stage6_34[6]}
   );
   gpc1_1 gpc4533 (
      {stage5_34[4]},
      {stage6_34[7]}
   );
   gpc1_1 gpc4534 (
      {stage5_34[5]},
      {stage6_34[8]}
   );
   gpc1_1 gpc4535 (
      {stage5_34[6]},
      {stage6_34[9]}
   );
   gpc1_1 gpc4536 (
      {stage5_34[7]},
      {stage6_34[10]}
   );
   gpc1_1 gpc4537 (
      {stage5_35[12]},
      {stage6_35[2]}
   );
   gpc1_1 gpc4538 (
      {stage5_35[13]},
      {stage6_35[3]}
   );
   gpc1_1 gpc4539 (
      {stage5_35[14]},
      {stage6_35[4]}
   );
   gpc1_1 gpc4540 (
      {stage5_36[0]},
      {stage6_36[2]}
   );
   gpc1_1 gpc4541 (
      {stage5_36[1]},
      {stage6_36[3]}
   );
   gpc1_1 gpc4542 (
      {stage5_36[2]},
      {stage6_36[4]}
   );
   gpc1_1 gpc4543 (
      {stage5_36[3]},
      {stage6_36[5]}
   );
   gpc1_1 gpc4544 (
      {stage5_38[0]},
      {stage6_38[1]}
   );
   gpc1_1 gpc4545 (
      {stage5_38[1]},
      {stage6_38[2]}
   );
   gpc223_4 gpc4546 (
      {stage6_5[0], stage6_5[1], stage6_5[2]},
      {stage6_6[0], stage6_6[1]},
      {stage6_7[0], stage6_7[1]},
      {stage7_8[0],stage7_7[0],stage7_6[0],stage7_5[0]}
   );
   gpc135_4 gpc4547 (
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4]},
      {stage6_10[0], stage6_10[1], stage6_10[2]},
      {stage6_11[0]},
      {stage7_12[0],stage7_11[0],stage7_10[0],stage7_9[0]}
   );
   gpc615_5 gpc4548 (
      {stage6_11[1], stage6_11[2], stage6_11[3], stage6_11[4], stage6_11[5]},
      {stage6_12[0]},
      {stage6_13[0], stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5]},
      {stage7_15[0],stage7_14[0],stage7_13[0],stage7_12[1],stage7_11[1]}
   );
   gpc2135_5 gpc4549 (
      {stage6_12[1], stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage6_13[6], stage6_13[7], stage6_13[8]},
      {stage6_14[0]},
      {stage6_15[0], stage6_15[1]},
      {stage7_16[0],stage7_15[1],stage7_14[1],stage7_13[1],stage7_12[2]}
   );
   gpc615_5 gpc4550 (
      {stage6_16[0], stage6_16[1], stage6_16[2], stage6_16[3], stage6_16[4]},
      {stage6_17[0]},
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage7_20[0],stage7_19[0],stage7_18[0],stage7_17[0],stage7_16[1]}
   );
   gpc7_3 gpc4551 (
      {stage6_17[1], stage6_17[2], stage6_17[3], stage6_17[4], stage6_17[5], stage6_17[6], stage6_17[7]},
      {stage7_19[1],stage7_18[1],stage7_17[1]}
   );
   gpc615_5 gpc4552 (
      {stage6_19[0], stage6_19[1], stage6_19[2], stage6_19[3], stage6_19[4]},
      {stage6_20[0]},
      {stage6_21[0], stage6_21[1], stage6_21[2], stage6_21[3], stage6_21[4], stage6_21[5]},
      {stage7_23[0],stage7_22[0],stage7_21[0],stage7_20[1],stage7_19[2]}
   );
   gpc615_5 gpc4553 (
      {stage6_23[0], stage6_23[1], stage6_23[2], stage6_23[3], stage6_23[4]},
      {stage6_24[0]},
      {stage6_25[0], stage6_25[1], stage6_25[2], stage6_25[3], stage6_25[4], 1'b0},
      {stage7_27[0],stage7_26[0],stage7_25[0],stage7_24[0],stage7_23[1]}
   );
   gpc7_3 gpc4554 (
      {stage6_26[0], stage6_26[1], stage6_26[2], stage6_26[3], stage6_26[4], stage6_26[5], stage6_26[6]},
      {stage7_28[0],stage7_27[1],stage7_26[1]}
   );
   gpc7_3 gpc4555 (
      {stage6_26[7], stage6_26[8], stage6_26[9], stage6_26[10], stage6_26[11], 1'b0, 1'b0},
      {stage7_28[1],stage7_27[2],stage7_26[2]}
   );
   gpc7_3 gpc4556 (
      {stage6_27[0], stage6_27[1], stage6_27[2], stage6_27[3], stage6_27[4], stage6_27[5], stage6_27[6]},
      {stage7_29[0],stage7_28[2],stage7_27[3]}
   );
   gpc1325_5 gpc4557 (
      {stage6_28[0], stage6_28[1], stage6_28[2], stage6_28[3], stage6_28[4]},
      {stage6_29[0], stage6_29[1]},
      {stage6_30[0], stage6_30[1], stage6_30[2]},
      {stage6_31[0]},
      {stage7_32[0],stage7_31[0],stage7_30[0],stage7_29[1],stage7_28[3]}
   );
   gpc7_3 gpc4558 (
      {stage6_31[1], stage6_31[2], stage6_31[3], stage6_31[4], stage6_31[5], stage6_31[6], stage6_31[7]},
      {stage7_33[0],stage7_32[1],stage7_31[1]}
   );
   gpc606_5 gpc4559 (
      {stage6_33[0], stage6_33[1], stage6_33[2], stage6_33[3], stage6_33[4], stage6_33[5]},
      {stage6_35[0], stage6_35[1], stage6_35[2], stage6_35[3], stage6_35[4], 1'b0},
      {stage7_37[0],stage7_36[0],stage7_35[0],stage7_34[0],stage7_33[1]}
   );
   gpc606_5 gpc4560 (
      {stage6_34[0], stage6_34[1], stage6_34[2], stage6_34[3], stage6_34[4], stage6_34[5]},
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3], stage6_36[4], stage6_36[5]},
      {stage7_38[0],stage7_37[1],stage7_36[1],stage7_35[1],stage7_34[1]}
   );
   gpc1_1 gpc4561 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc4562 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc4563 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc4564 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc4565 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc4566 (
      {stage6_1[2]},
      {stage7_1[2]}
   );
   gpc1_1 gpc4567 (
      {stage6_1[3]},
      {stage7_1[3]}
   );
   gpc1_1 gpc4568 (
      {stage6_1[4]},
      {stage7_1[4]}
   );
   gpc1_1 gpc4569 (
      {stage6_1[5]},
      {stage7_1[5]}
   );
   gpc1_1 gpc4570 (
      {stage6_1[6]},
      {stage7_1[6]}
   );
   gpc1_1 gpc4571 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc4572 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc4573 (
      {stage6_3[1]},
      {stage7_3[1]}
   );
   gpc1_1 gpc4574 (
      {stage6_3[2]},
      {stage7_3[2]}
   );
   gpc1_1 gpc4575 (
      {stage6_3[3]},
      {stage7_3[3]}
   );
   gpc1_1 gpc4576 (
      {stage6_4[0]},
      {stage7_4[0]}
   );
   gpc1_1 gpc4577 (
      {stage6_4[1]},
      {stage7_4[1]}
   );
   gpc1_1 gpc4578 (
      {stage6_5[3]},
      {stage7_5[1]}
   );
   gpc1_1 gpc4579 (
      {stage6_5[4]},
      {stage7_5[2]}
   );
   gpc1_1 gpc4580 (
      {stage6_5[5]},
      {stage7_5[3]}
   );
   gpc1_1 gpc4581 (
      {stage6_6[2]},
      {stage7_6[1]}
   );
   gpc1_1 gpc4582 (
      {stage6_6[3]},
      {stage7_6[2]}
   );
   gpc1_1 gpc4583 (
      {stage6_6[4]},
      {stage7_6[3]}
   );
   gpc1_1 gpc4584 (
      {stage6_7[2]},
      {stage7_7[1]}
   );
   gpc1_1 gpc4585 (
      {stage6_8[0]},
      {stage7_8[1]}
   );
   gpc1_1 gpc4586 (
      {stage6_8[1]},
      {stage7_8[2]}
   );
   gpc1_1 gpc4587 (
      {stage6_8[2]},
      {stage7_8[3]}
   );
   gpc1_1 gpc4588 (
      {stage6_8[3]},
      {stage7_8[4]}
   );
   gpc1_1 gpc4589 (
      {stage6_8[4]},
      {stage7_8[5]}
   );
   gpc1_1 gpc4590 (
      {stage6_8[5]},
      {stage7_8[6]}
   );
   gpc1_1 gpc4591 (
      {stage6_10[3]},
      {stage7_10[1]}
   );
   gpc1_1 gpc4592 (
      {stage6_10[4]},
      {stage7_10[2]}
   );
   gpc1_1 gpc4593 (
      {stage6_10[5]},
      {stage7_10[3]}
   );
   gpc1_1 gpc4594 (
      {stage6_10[6]},
      {stage7_10[4]}
   );
   gpc1_1 gpc4595 (
      {stage6_12[6]},
      {stage7_12[3]}
   );
   gpc1_1 gpc4596 (
      {stage6_14[1]},
      {stage7_14[2]}
   );
   gpc1_1 gpc4597 (
      {stage6_14[2]},
      {stage7_14[3]}
   );
   gpc1_1 gpc4598 (
      {stage6_14[3]},
      {stage7_14[4]}
   );
   gpc1_1 gpc4599 (
      {stage6_14[4]},
      {stage7_14[5]}
   );
   gpc1_1 gpc4600 (
      {stage6_14[5]},
      {stage7_14[6]}
   );
   gpc1_1 gpc4601 (
      {stage6_15[2]},
      {stage7_15[2]}
   );
   gpc1_1 gpc4602 (
      {stage6_15[3]},
      {stage7_15[3]}
   );
   gpc1_1 gpc4603 (
      {stage6_15[4]},
      {stage7_15[4]}
   );
   gpc1_1 gpc4604 (
      {stage6_15[5]},
      {stage7_15[5]}
   );
   gpc1_1 gpc4605 (
      {stage6_17[8]},
      {stage7_17[2]}
   );
   gpc1_1 gpc4606 (
      {stage6_17[9]},
      {stage7_17[3]}
   );
   gpc1_1 gpc4607 (
      {stage6_20[1]},
      {stage7_20[2]}
   );
   gpc1_1 gpc4608 (
      {stage6_20[2]},
      {stage7_20[3]}
   );
   gpc1_1 gpc4609 (
      {stage6_20[3]},
      {stage7_20[4]}
   );
   gpc1_1 gpc4610 (
      {stage6_20[4]},
      {stage7_20[5]}
   );
   gpc1_1 gpc4611 (
      {stage6_20[5]},
      {stage7_20[6]}
   );
   gpc1_1 gpc4612 (
      {stage6_22[0]},
      {stage7_22[1]}
   );
   gpc1_1 gpc4613 (
      {stage6_22[1]},
      {stage7_22[2]}
   );
   gpc1_1 gpc4614 (
      {stage6_22[2]},
      {stage7_22[3]}
   );
   gpc1_1 gpc4615 (
      {stage6_22[3]},
      {stage7_22[4]}
   );
   gpc1_1 gpc4616 (
      {stage6_22[4]},
      {stage7_22[5]}
   );
   gpc1_1 gpc4617 (
      {stage6_23[5]},
      {stage7_23[2]}
   );
   gpc1_1 gpc4618 (
      {stage6_23[6]},
      {stage7_23[3]}
   );
   gpc1_1 gpc4619 (
      {stage6_23[7]},
      {stage7_23[4]}
   );
   gpc1_1 gpc4620 (
      {stage6_23[8]},
      {stage7_23[5]}
   );
   gpc1_1 gpc4621 (
      {stage6_24[1]},
      {stage7_24[1]}
   );
   gpc1_1 gpc4622 (
      {stage6_24[2]},
      {stage7_24[2]}
   );
   gpc1_1 gpc4623 (
      {stage6_24[3]},
      {stage7_24[3]}
   );
   gpc1_1 gpc4624 (
      {stage6_27[7]},
      {stage7_27[4]}
   );
   gpc1_1 gpc4625 (
      {stage6_27[8]},
      {stage7_27[5]}
   );
   gpc1_1 gpc4626 (
      {stage6_28[5]},
      {stage7_28[4]}
   );
   gpc1_1 gpc4627 (
      {stage6_28[6]},
      {stage7_28[5]}
   );
   gpc1_1 gpc4628 (
      {stage6_29[2]},
      {stage7_29[2]}
   );
   gpc1_1 gpc4629 (
      {stage6_29[3]},
      {stage7_29[3]}
   );
   gpc1_1 gpc4630 (
      {stage6_30[3]},
      {stage7_30[1]}
   );
   gpc1_1 gpc4631 (
      {stage6_30[4]},
      {stage7_30[2]}
   );
   gpc1_1 gpc4632 (
      {stage6_32[0]},
      {stage7_32[2]}
   );
   gpc1_1 gpc4633 (
      {stage6_32[1]},
      {stage7_32[3]}
   );
   gpc1_1 gpc4634 (
      {stage6_32[2]},
      {stage7_32[4]}
   );
   gpc1_1 gpc4635 (
      {stage6_32[3]},
      {stage7_32[5]}
   );
   gpc1_1 gpc4636 (
      {stage6_34[6]},
      {stage7_34[2]}
   );
   gpc1_1 gpc4637 (
      {stage6_34[7]},
      {stage7_34[3]}
   );
   gpc1_1 gpc4638 (
      {stage6_34[8]},
      {stage7_34[4]}
   );
   gpc1_1 gpc4639 (
      {stage6_34[9]},
      {stage7_34[5]}
   );
   gpc1_1 gpc4640 (
      {stage6_34[10]},
      {stage7_34[6]}
   );
   gpc1_1 gpc4641 (
      {stage6_37[0]},
      {stage7_37[2]}
   );
   gpc1_1 gpc4642 (
      {stage6_37[1]},
      {stage7_37[3]}
   );
   gpc1_1 gpc4643 (
      {stage6_38[0]},
      {stage7_38[1]}
   );
   gpc1_1 gpc4644 (
      {stage6_38[1]},
      {stage7_38[2]}
   );
   gpc1_1 gpc4645 (
      {stage6_38[2]},
      {stage7_38[3]}
   );
   gpc1_1 gpc4646 (
      {stage6_39[0]},
      {stage7_39[0]}
   );
   gpc1163_5 gpc4647 (
      {stage7_0[0], stage7_0[1], stage7_0[2]},
      {stage7_1[0], stage7_1[1], stage7_1[2], stage7_1[3], stage7_1[4], stage7_1[5]},
      {stage7_2[0]},
      {stage7_3[0]},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc1423_5 gpc4648 (
      {stage7_3[1], stage7_3[2], stage7_3[3]},
      {stage7_4[0], stage7_4[1]},
      {stage7_5[0], stage7_5[1], stage7_5[2], stage7_5[3]},
      {stage7_6[0]},
      {stage8_7[0],stage8_6[0],stage8_5[0],stage8_4[1],stage8_3[1]}
   );
   gpc623_5 gpc4649 (
      {stage7_6[1], stage7_6[2], stage7_6[3]},
      {stage7_7[0], stage7_7[1]},
      {stage7_8[0], stage7_8[1], stage7_8[2], stage7_8[3], stage7_8[4], stage7_8[5]},
      {stage8_10[0],stage8_9[0],stage8_8[0],stage8_7[1],stage8_6[1]}
   );
   gpc1325_5 gpc4650 (
      {stage7_10[0], stage7_10[1], stage7_10[2], stage7_10[3], stage7_10[4]},
      {stage7_11[0], stage7_11[1]},
      {stage7_12[0], stage7_12[1], stage7_12[2]},
      {stage7_13[0]},
      {stage8_14[0],stage8_13[0],stage8_12[0],stage8_11[0],stage8_10[1]}
   );
   gpc117_4 gpc4651 (
      {stage7_14[0], stage7_14[1], stage7_14[2], stage7_14[3], stage7_14[4], stage7_14[5], stage7_14[6]},
      {stage7_15[0]},
      {stage7_16[0]},
      {stage8_17[0],stage8_16[0],stage8_15[0],stage8_14[1]}
   );
   gpc1415_5 gpc4652 (
      {stage7_15[1], stage7_15[2], stage7_15[3], stage7_15[4], stage7_15[5]},
      {stage7_16[1]},
      {stage7_17[0], stage7_17[1], stage7_17[2], stage7_17[3]},
      {stage7_18[0]},
      {stage8_19[0],stage8_18[0],stage8_17[1],stage8_16[1],stage8_15[1]}
   );
   gpc3_2 gpc4653 (
      {stage7_19[0], stage7_19[1], stage7_19[2]},
      {stage8_20[0],stage8_19[1]}
   );
   gpc7_3 gpc4654 (
      {stage7_20[0], stage7_20[1], stage7_20[2], stage7_20[3], stage7_20[4], stage7_20[5], stage7_20[6]},
      {stage8_22[0],stage8_21[0],stage8_20[1]}
   );
   gpc117_4 gpc4655 (
      {stage7_22[0], stage7_22[1], stage7_22[2], stage7_22[3], stage7_22[4], stage7_22[5], 1'b0},
      {stage7_23[0]},
      {stage7_24[0]},
      {stage8_25[0],stage8_24[0],stage8_23[0],stage8_22[1]}
   );
   gpc2135_5 gpc4656 (
      {stage7_23[1], stage7_23[2], stage7_23[3], stage7_23[4], stage7_23[5]},
      {stage7_24[1], stage7_24[2], stage7_24[3]},
      {stage7_25[0]},
      {stage7_26[0], stage7_26[1]},
      {stage8_27[0],stage8_26[0],stage8_25[1],stage8_24[1],stage8_23[1]}
   );
   gpc2116_5 gpc4657 (
      {stage7_27[0], stage7_27[1], stage7_27[2], stage7_27[3], stage7_27[4], stage7_27[5]},
      {stage7_28[0]},
      {stage7_29[0]},
      {stage7_30[0], stage7_30[1]},
      {stage8_31[0],stage8_30[0],stage8_29[0],stage8_28[0],stage8_27[1]}
   );
   gpc2135_5 gpc4658 (
      {stage7_28[1], stage7_28[2], stage7_28[3], stage7_28[4], stage7_28[5]},
      {stage7_29[1], stage7_29[2], stage7_29[3]},
      {stage7_30[2]},
      {stage7_31[0], stage7_31[1]},
      {stage8_32[0],stage8_31[1],stage8_30[1],stage8_29[1],stage8_28[1]}
   );
   gpc2116_5 gpc4659 (
      {stage7_32[0], stage7_32[1], stage7_32[2], stage7_32[3], stage7_32[4], stage7_32[5]},
      {stage7_33[0]},
      {stage7_34[0]},
      {stage7_35[0], stage7_35[1]},
      {stage8_36[0],stage8_35[0],stage8_34[0],stage8_33[0],stage8_32[1]}
   );
   gpc207_4 gpc4660 (
      {stage7_34[1], stage7_34[2], stage7_34[3], stage7_34[4], stage7_34[5], stage7_34[6], 1'b0},
      {stage7_36[0], stage7_36[1]},
      {stage8_37[0],stage8_36[1],stage8_35[1],stage8_34[1]}
   );
   gpc135_4 gpc4661 (
      {stage7_37[0], stage7_37[1], stage7_37[2], stage7_37[3], 1'b0},
      {stage7_38[0], stage7_38[1], stage7_38[2]},
      {stage7_39[0]},
      {stage8_40[0],stage8_39[0],stage8_38[0],stage8_37[1]}
   );
   gpc1_1 gpc4662 (
      {stage7_1[6]},
      {stage8_1[1]}
   );
   gpc1_1 gpc4663 (
      {stage7_8[6]},
      {stage8_8[1]}
   );
   gpc1_1 gpc4664 (
      {stage7_9[0]},
      {stage8_9[1]}
   );
   gpc1_1 gpc4665 (
      {stage7_12[3]},
      {stage8_12[1]}
   );
   gpc1_1 gpc4666 (
      {stage7_13[1]},
      {stage8_13[1]}
   );
   gpc1_1 gpc4667 (
      {stage7_18[1]},
      {stage8_18[1]}
   );
   gpc1_1 gpc4668 (
      {stage7_21[0]},
      {stage8_21[1]}
   );
   gpc1_1 gpc4669 (
      {stage7_26[2]},
      {stage8_26[1]}
   );
   gpc1_1 gpc4670 (
      {stage7_33[1]},
      {stage8_33[1]}
   );
   gpc1_1 gpc4671 (
      {stage7_38[3]},
      {stage8_38[1]}
   );
endmodule

module testbench();
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    reg [485:0] src16;
    reg [485:0] src17;
    reg [485:0] src18;
    reg [485:0] src19;
    reg [485:0] src20;
    reg [485:0] src21;
    reg [485:0] src22;
    reg [485:0] src23;
    reg [485:0] src24;
    reg [485:0] src25;
    reg [485:0] src26;
    reg [485:0] src27;
    reg [485:0] src28;
    reg [485:0] src29;
    reg [485:0] src30;
    reg [485:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [40:0] srcsum;
    wire [40:0] dstsum;
    wire test;
    compressor_CLA486_32 compressor_CLA486_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255] + src16[256] + src16[257] + src16[258] + src16[259] + src16[260] + src16[261] + src16[262] + src16[263] + src16[264] + src16[265] + src16[266] + src16[267] + src16[268] + src16[269] + src16[270] + src16[271] + src16[272] + src16[273] + src16[274] + src16[275] + src16[276] + src16[277] + src16[278] + src16[279] + src16[280] + src16[281] + src16[282] + src16[283] + src16[284] + src16[285] + src16[286] + src16[287] + src16[288] + src16[289] + src16[290] + src16[291] + src16[292] + src16[293] + src16[294] + src16[295] + src16[296] + src16[297] + src16[298] + src16[299] + src16[300] + src16[301] + src16[302] + src16[303] + src16[304] + src16[305] + src16[306] + src16[307] + src16[308] + src16[309] + src16[310] + src16[311] + src16[312] + src16[313] + src16[314] + src16[315] + src16[316] + src16[317] + src16[318] + src16[319] + src16[320] + src16[321] + src16[322] + src16[323] + src16[324] + src16[325] + src16[326] + src16[327] + src16[328] + src16[329] + src16[330] + src16[331] + src16[332] + src16[333] + src16[334] + src16[335] + src16[336] + src16[337] + src16[338] + src16[339] + src16[340] + src16[341] + src16[342] + src16[343] + src16[344] + src16[345] + src16[346] + src16[347] + src16[348] + src16[349] + src16[350] + src16[351] + src16[352] + src16[353] + src16[354] + src16[355] + src16[356] + src16[357] + src16[358] + src16[359] + src16[360] + src16[361] + src16[362] + src16[363] + src16[364] + src16[365] + src16[366] + src16[367] + src16[368] + src16[369] + src16[370] + src16[371] + src16[372] + src16[373] + src16[374] + src16[375] + src16[376] + src16[377] + src16[378] + src16[379] + src16[380] + src16[381] + src16[382] + src16[383] + src16[384] + src16[385] + src16[386] + src16[387] + src16[388] + src16[389] + src16[390] + src16[391] + src16[392] + src16[393] + src16[394] + src16[395] + src16[396] + src16[397] + src16[398] + src16[399] + src16[400] + src16[401] + src16[402] + src16[403] + src16[404] + src16[405] + src16[406] + src16[407] + src16[408] + src16[409] + src16[410] + src16[411] + src16[412] + src16[413] + src16[414] + src16[415] + src16[416] + src16[417] + src16[418] + src16[419] + src16[420] + src16[421] + src16[422] + src16[423] + src16[424] + src16[425] + src16[426] + src16[427] + src16[428] + src16[429] + src16[430] + src16[431] + src16[432] + src16[433] + src16[434] + src16[435] + src16[436] + src16[437] + src16[438] + src16[439] + src16[440] + src16[441] + src16[442] + src16[443] + src16[444] + src16[445] + src16[446] + src16[447] + src16[448] + src16[449] + src16[450] + src16[451] + src16[452] + src16[453] + src16[454] + src16[455] + src16[456] + src16[457] + src16[458] + src16[459] + src16[460] + src16[461] + src16[462] + src16[463] + src16[464] + src16[465] + src16[466] + src16[467] + src16[468] + src16[469] + src16[470] + src16[471] + src16[472] + src16[473] + src16[474] + src16[475] + src16[476] + src16[477] + src16[478] + src16[479] + src16[480] + src16[481] + src16[482] + src16[483] + src16[484] + src16[485])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255] + src17[256] + src17[257] + src17[258] + src17[259] + src17[260] + src17[261] + src17[262] + src17[263] + src17[264] + src17[265] + src17[266] + src17[267] + src17[268] + src17[269] + src17[270] + src17[271] + src17[272] + src17[273] + src17[274] + src17[275] + src17[276] + src17[277] + src17[278] + src17[279] + src17[280] + src17[281] + src17[282] + src17[283] + src17[284] + src17[285] + src17[286] + src17[287] + src17[288] + src17[289] + src17[290] + src17[291] + src17[292] + src17[293] + src17[294] + src17[295] + src17[296] + src17[297] + src17[298] + src17[299] + src17[300] + src17[301] + src17[302] + src17[303] + src17[304] + src17[305] + src17[306] + src17[307] + src17[308] + src17[309] + src17[310] + src17[311] + src17[312] + src17[313] + src17[314] + src17[315] + src17[316] + src17[317] + src17[318] + src17[319] + src17[320] + src17[321] + src17[322] + src17[323] + src17[324] + src17[325] + src17[326] + src17[327] + src17[328] + src17[329] + src17[330] + src17[331] + src17[332] + src17[333] + src17[334] + src17[335] + src17[336] + src17[337] + src17[338] + src17[339] + src17[340] + src17[341] + src17[342] + src17[343] + src17[344] + src17[345] + src17[346] + src17[347] + src17[348] + src17[349] + src17[350] + src17[351] + src17[352] + src17[353] + src17[354] + src17[355] + src17[356] + src17[357] + src17[358] + src17[359] + src17[360] + src17[361] + src17[362] + src17[363] + src17[364] + src17[365] + src17[366] + src17[367] + src17[368] + src17[369] + src17[370] + src17[371] + src17[372] + src17[373] + src17[374] + src17[375] + src17[376] + src17[377] + src17[378] + src17[379] + src17[380] + src17[381] + src17[382] + src17[383] + src17[384] + src17[385] + src17[386] + src17[387] + src17[388] + src17[389] + src17[390] + src17[391] + src17[392] + src17[393] + src17[394] + src17[395] + src17[396] + src17[397] + src17[398] + src17[399] + src17[400] + src17[401] + src17[402] + src17[403] + src17[404] + src17[405] + src17[406] + src17[407] + src17[408] + src17[409] + src17[410] + src17[411] + src17[412] + src17[413] + src17[414] + src17[415] + src17[416] + src17[417] + src17[418] + src17[419] + src17[420] + src17[421] + src17[422] + src17[423] + src17[424] + src17[425] + src17[426] + src17[427] + src17[428] + src17[429] + src17[430] + src17[431] + src17[432] + src17[433] + src17[434] + src17[435] + src17[436] + src17[437] + src17[438] + src17[439] + src17[440] + src17[441] + src17[442] + src17[443] + src17[444] + src17[445] + src17[446] + src17[447] + src17[448] + src17[449] + src17[450] + src17[451] + src17[452] + src17[453] + src17[454] + src17[455] + src17[456] + src17[457] + src17[458] + src17[459] + src17[460] + src17[461] + src17[462] + src17[463] + src17[464] + src17[465] + src17[466] + src17[467] + src17[468] + src17[469] + src17[470] + src17[471] + src17[472] + src17[473] + src17[474] + src17[475] + src17[476] + src17[477] + src17[478] + src17[479] + src17[480] + src17[481] + src17[482] + src17[483] + src17[484] + src17[485])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255] + src18[256] + src18[257] + src18[258] + src18[259] + src18[260] + src18[261] + src18[262] + src18[263] + src18[264] + src18[265] + src18[266] + src18[267] + src18[268] + src18[269] + src18[270] + src18[271] + src18[272] + src18[273] + src18[274] + src18[275] + src18[276] + src18[277] + src18[278] + src18[279] + src18[280] + src18[281] + src18[282] + src18[283] + src18[284] + src18[285] + src18[286] + src18[287] + src18[288] + src18[289] + src18[290] + src18[291] + src18[292] + src18[293] + src18[294] + src18[295] + src18[296] + src18[297] + src18[298] + src18[299] + src18[300] + src18[301] + src18[302] + src18[303] + src18[304] + src18[305] + src18[306] + src18[307] + src18[308] + src18[309] + src18[310] + src18[311] + src18[312] + src18[313] + src18[314] + src18[315] + src18[316] + src18[317] + src18[318] + src18[319] + src18[320] + src18[321] + src18[322] + src18[323] + src18[324] + src18[325] + src18[326] + src18[327] + src18[328] + src18[329] + src18[330] + src18[331] + src18[332] + src18[333] + src18[334] + src18[335] + src18[336] + src18[337] + src18[338] + src18[339] + src18[340] + src18[341] + src18[342] + src18[343] + src18[344] + src18[345] + src18[346] + src18[347] + src18[348] + src18[349] + src18[350] + src18[351] + src18[352] + src18[353] + src18[354] + src18[355] + src18[356] + src18[357] + src18[358] + src18[359] + src18[360] + src18[361] + src18[362] + src18[363] + src18[364] + src18[365] + src18[366] + src18[367] + src18[368] + src18[369] + src18[370] + src18[371] + src18[372] + src18[373] + src18[374] + src18[375] + src18[376] + src18[377] + src18[378] + src18[379] + src18[380] + src18[381] + src18[382] + src18[383] + src18[384] + src18[385] + src18[386] + src18[387] + src18[388] + src18[389] + src18[390] + src18[391] + src18[392] + src18[393] + src18[394] + src18[395] + src18[396] + src18[397] + src18[398] + src18[399] + src18[400] + src18[401] + src18[402] + src18[403] + src18[404] + src18[405] + src18[406] + src18[407] + src18[408] + src18[409] + src18[410] + src18[411] + src18[412] + src18[413] + src18[414] + src18[415] + src18[416] + src18[417] + src18[418] + src18[419] + src18[420] + src18[421] + src18[422] + src18[423] + src18[424] + src18[425] + src18[426] + src18[427] + src18[428] + src18[429] + src18[430] + src18[431] + src18[432] + src18[433] + src18[434] + src18[435] + src18[436] + src18[437] + src18[438] + src18[439] + src18[440] + src18[441] + src18[442] + src18[443] + src18[444] + src18[445] + src18[446] + src18[447] + src18[448] + src18[449] + src18[450] + src18[451] + src18[452] + src18[453] + src18[454] + src18[455] + src18[456] + src18[457] + src18[458] + src18[459] + src18[460] + src18[461] + src18[462] + src18[463] + src18[464] + src18[465] + src18[466] + src18[467] + src18[468] + src18[469] + src18[470] + src18[471] + src18[472] + src18[473] + src18[474] + src18[475] + src18[476] + src18[477] + src18[478] + src18[479] + src18[480] + src18[481] + src18[482] + src18[483] + src18[484] + src18[485])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255] + src19[256] + src19[257] + src19[258] + src19[259] + src19[260] + src19[261] + src19[262] + src19[263] + src19[264] + src19[265] + src19[266] + src19[267] + src19[268] + src19[269] + src19[270] + src19[271] + src19[272] + src19[273] + src19[274] + src19[275] + src19[276] + src19[277] + src19[278] + src19[279] + src19[280] + src19[281] + src19[282] + src19[283] + src19[284] + src19[285] + src19[286] + src19[287] + src19[288] + src19[289] + src19[290] + src19[291] + src19[292] + src19[293] + src19[294] + src19[295] + src19[296] + src19[297] + src19[298] + src19[299] + src19[300] + src19[301] + src19[302] + src19[303] + src19[304] + src19[305] + src19[306] + src19[307] + src19[308] + src19[309] + src19[310] + src19[311] + src19[312] + src19[313] + src19[314] + src19[315] + src19[316] + src19[317] + src19[318] + src19[319] + src19[320] + src19[321] + src19[322] + src19[323] + src19[324] + src19[325] + src19[326] + src19[327] + src19[328] + src19[329] + src19[330] + src19[331] + src19[332] + src19[333] + src19[334] + src19[335] + src19[336] + src19[337] + src19[338] + src19[339] + src19[340] + src19[341] + src19[342] + src19[343] + src19[344] + src19[345] + src19[346] + src19[347] + src19[348] + src19[349] + src19[350] + src19[351] + src19[352] + src19[353] + src19[354] + src19[355] + src19[356] + src19[357] + src19[358] + src19[359] + src19[360] + src19[361] + src19[362] + src19[363] + src19[364] + src19[365] + src19[366] + src19[367] + src19[368] + src19[369] + src19[370] + src19[371] + src19[372] + src19[373] + src19[374] + src19[375] + src19[376] + src19[377] + src19[378] + src19[379] + src19[380] + src19[381] + src19[382] + src19[383] + src19[384] + src19[385] + src19[386] + src19[387] + src19[388] + src19[389] + src19[390] + src19[391] + src19[392] + src19[393] + src19[394] + src19[395] + src19[396] + src19[397] + src19[398] + src19[399] + src19[400] + src19[401] + src19[402] + src19[403] + src19[404] + src19[405] + src19[406] + src19[407] + src19[408] + src19[409] + src19[410] + src19[411] + src19[412] + src19[413] + src19[414] + src19[415] + src19[416] + src19[417] + src19[418] + src19[419] + src19[420] + src19[421] + src19[422] + src19[423] + src19[424] + src19[425] + src19[426] + src19[427] + src19[428] + src19[429] + src19[430] + src19[431] + src19[432] + src19[433] + src19[434] + src19[435] + src19[436] + src19[437] + src19[438] + src19[439] + src19[440] + src19[441] + src19[442] + src19[443] + src19[444] + src19[445] + src19[446] + src19[447] + src19[448] + src19[449] + src19[450] + src19[451] + src19[452] + src19[453] + src19[454] + src19[455] + src19[456] + src19[457] + src19[458] + src19[459] + src19[460] + src19[461] + src19[462] + src19[463] + src19[464] + src19[465] + src19[466] + src19[467] + src19[468] + src19[469] + src19[470] + src19[471] + src19[472] + src19[473] + src19[474] + src19[475] + src19[476] + src19[477] + src19[478] + src19[479] + src19[480] + src19[481] + src19[482] + src19[483] + src19[484] + src19[485])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255] + src20[256] + src20[257] + src20[258] + src20[259] + src20[260] + src20[261] + src20[262] + src20[263] + src20[264] + src20[265] + src20[266] + src20[267] + src20[268] + src20[269] + src20[270] + src20[271] + src20[272] + src20[273] + src20[274] + src20[275] + src20[276] + src20[277] + src20[278] + src20[279] + src20[280] + src20[281] + src20[282] + src20[283] + src20[284] + src20[285] + src20[286] + src20[287] + src20[288] + src20[289] + src20[290] + src20[291] + src20[292] + src20[293] + src20[294] + src20[295] + src20[296] + src20[297] + src20[298] + src20[299] + src20[300] + src20[301] + src20[302] + src20[303] + src20[304] + src20[305] + src20[306] + src20[307] + src20[308] + src20[309] + src20[310] + src20[311] + src20[312] + src20[313] + src20[314] + src20[315] + src20[316] + src20[317] + src20[318] + src20[319] + src20[320] + src20[321] + src20[322] + src20[323] + src20[324] + src20[325] + src20[326] + src20[327] + src20[328] + src20[329] + src20[330] + src20[331] + src20[332] + src20[333] + src20[334] + src20[335] + src20[336] + src20[337] + src20[338] + src20[339] + src20[340] + src20[341] + src20[342] + src20[343] + src20[344] + src20[345] + src20[346] + src20[347] + src20[348] + src20[349] + src20[350] + src20[351] + src20[352] + src20[353] + src20[354] + src20[355] + src20[356] + src20[357] + src20[358] + src20[359] + src20[360] + src20[361] + src20[362] + src20[363] + src20[364] + src20[365] + src20[366] + src20[367] + src20[368] + src20[369] + src20[370] + src20[371] + src20[372] + src20[373] + src20[374] + src20[375] + src20[376] + src20[377] + src20[378] + src20[379] + src20[380] + src20[381] + src20[382] + src20[383] + src20[384] + src20[385] + src20[386] + src20[387] + src20[388] + src20[389] + src20[390] + src20[391] + src20[392] + src20[393] + src20[394] + src20[395] + src20[396] + src20[397] + src20[398] + src20[399] + src20[400] + src20[401] + src20[402] + src20[403] + src20[404] + src20[405] + src20[406] + src20[407] + src20[408] + src20[409] + src20[410] + src20[411] + src20[412] + src20[413] + src20[414] + src20[415] + src20[416] + src20[417] + src20[418] + src20[419] + src20[420] + src20[421] + src20[422] + src20[423] + src20[424] + src20[425] + src20[426] + src20[427] + src20[428] + src20[429] + src20[430] + src20[431] + src20[432] + src20[433] + src20[434] + src20[435] + src20[436] + src20[437] + src20[438] + src20[439] + src20[440] + src20[441] + src20[442] + src20[443] + src20[444] + src20[445] + src20[446] + src20[447] + src20[448] + src20[449] + src20[450] + src20[451] + src20[452] + src20[453] + src20[454] + src20[455] + src20[456] + src20[457] + src20[458] + src20[459] + src20[460] + src20[461] + src20[462] + src20[463] + src20[464] + src20[465] + src20[466] + src20[467] + src20[468] + src20[469] + src20[470] + src20[471] + src20[472] + src20[473] + src20[474] + src20[475] + src20[476] + src20[477] + src20[478] + src20[479] + src20[480] + src20[481] + src20[482] + src20[483] + src20[484] + src20[485])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255] + src21[256] + src21[257] + src21[258] + src21[259] + src21[260] + src21[261] + src21[262] + src21[263] + src21[264] + src21[265] + src21[266] + src21[267] + src21[268] + src21[269] + src21[270] + src21[271] + src21[272] + src21[273] + src21[274] + src21[275] + src21[276] + src21[277] + src21[278] + src21[279] + src21[280] + src21[281] + src21[282] + src21[283] + src21[284] + src21[285] + src21[286] + src21[287] + src21[288] + src21[289] + src21[290] + src21[291] + src21[292] + src21[293] + src21[294] + src21[295] + src21[296] + src21[297] + src21[298] + src21[299] + src21[300] + src21[301] + src21[302] + src21[303] + src21[304] + src21[305] + src21[306] + src21[307] + src21[308] + src21[309] + src21[310] + src21[311] + src21[312] + src21[313] + src21[314] + src21[315] + src21[316] + src21[317] + src21[318] + src21[319] + src21[320] + src21[321] + src21[322] + src21[323] + src21[324] + src21[325] + src21[326] + src21[327] + src21[328] + src21[329] + src21[330] + src21[331] + src21[332] + src21[333] + src21[334] + src21[335] + src21[336] + src21[337] + src21[338] + src21[339] + src21[340] + src21[341] + src21[342] + src21[343] + src21[344] + src21[345] + src21[346] + src21[347] + src21[348] + src21[349] + src21[350] + src21[351] + src21[352] + src21[353] + src21[354] + src21[355] + src21[356] + src21[357] + src21[358] + src21[359] + src21[360] + src21[361] + src21[362] + src21[363] + src21[364] + src21[365] + src21[366] + src21[367] + src21[368] + src21[369] + src21[370] + src21[371] + src21[372] + src21[373] + src21[374] + src21[375] + src21[376] + src21[377] + src21[378] + src21[379] + src21[380] + src21[381] + src21[382] + src21[383] + src21[384] + src21[385] + src21[386] + src21[387] + src21[388] + src21[389] + src21[390] + src21[391] + src21[392] + src21[393] + src21[394] + src21[395] + src21[396] + src21[397] + src21[398] + src21[399] + src21[400] + src21[401] + src21[402] + src21[403] + src21[404] + src21[405] + src21[406] + src21[407] + src21[408] + src21[409] + src21[410] + src21[411] + src21[412] + src21[413] + src21[414] + src21[415] + src21[416] + src21[417] + src21[418] + src21[419] + src21[420] + src21[421] + src21[422] + src21[423] + src21[424] + src21[425] + src21[426] + src21[427] + src21[428] + src21[429] + src21[430] + src21[431] + src21[432] + src21[433] + src21[434] + src21[435] + src21[436] + src21[437] + src21[438] + src21[439] + src21[440] + src21[441] + src21[442] + src21[443] + src21[444] + src21[445] + src21[446] + src21[447] + src21[448] + src21[449] + src21[450] + src21[451] + src21[452] + src21[453] + src21[454] + src21[455] + src21[456] + src21[457] + src21[458] + src21[459] + src21[460] + src21[461] + src21[462] + src21[463] + src21[464] + src21[465] + src21[466] + src21[467] + src21[468] + src21[469] + src21[470] + src21[471] + src21[472] + src21[473] + src21[474] + src21[475] + src21[476] + src21[477] + src21[478] + src21[479] + src21[480] + src21[481] + src21[482] + src21[483] + src21[484] + src21[485])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255] + src22[256] + src22[257] + src22[258] + src22[259] + src22[260] + src22[261] + src22[262] + src22[263] + src22[264] + src22[265] + src22[266] + src22[267] + src22[268] + src22[269] + src22[270] + src22[271] + src22[272] + src22[273] + src22[274] + src22[275] + src22[276] + src22[277] + src22[278] + src22[279] + src22[280] + src22[281] + src22[282] + src22[283] + src22[284] + src22[285] + src22[286] + src22[287] + src22[288] + src22[289] + src22[290] + src22[291] + src22[292] + src22[293] + src22[294] + src22[295] + src22[296] + src22[297] + src22[298] + src22[299] + src22[300] + src22[301] + src22[302] + src22[303] + src22[304] + src22[305] + src22[306] + src22[307] + src22[308] + src22[309] + src22[310] + src22[311] + src22[312] + src22[313] + src22[314] + src22[315] + src22[316] + src22[317] + src22[318] + src22[319] + src22[320] + src22[321] + src22[322] + src22[323] + src22[324] + src22[325] + src22[326] + src22[327] + src22[328] + src22[329] + src22[330] + src22[331] + src22[332] + src22[333] + src22[334] + src22[335] + src22[336] + src22[337] + src22[338] + src22[339] + src22[340] + src22[341] + src22[342] + src22[343] + src22[344] + src22[345] + src22[346] + src22[347] + src22[348] + src22[349] + src22[350] + src22[351] + src22[352] + src22[353] + src22[354] + src22[355] + src22[356] + src22[357] + src22[358] + src22[359] + src22[360] + src22[361] + src22[362] + src22[363] + src22[364] + src22[365] + src22[366] + src22[367] + src22[368] + src22[369] + src22[370] + src22[371] + src22[372] + src22[373] + src22[374] + src22[375] + src22[376] + src22[377] + src22[378] + src22[379] + src22[380] + src22[381] + src22[382] + src22[383] + src22[384] + src22[385] + src22[386] + src22[387] + src22[388] + src22[389] + src22[390] + src22[391] + src22[392] + src22[393] + src22[394] + src22[395] + src22[396] + src22[397] + src22[398] + src22[399] + src22[400] + src22[401] + src22[402] + src22[403] + src22[404] + src22[405] + src22[406] + src22[407] + src22[408] + src22[409] + src22[410] + src22[411] + src22[412] + src22[413] + src22[414] + src22[415] + src22[416] + src22[417] + src22[418] + src22[419] + src22[420] + src22[421] + src22[422] + src22[423] + src22[424] + src22[425] + src22[426] + src22[427] + src22[428] + src22[429] + src22[430] + src22[431] + src22[432] + src22[433] + src22[434] + src22[435] + src22[436] + src22[437] + src22[438] + src22[439] + src22[440] + src22[441] + src22[442] + src22[443] + src22[444] + src22[445] + src22[446] + src22[447] + src22[448] + src22[449] + src22[450] + src22[451] + src22[452] + src22[453] + src22[454] + src22[455] + src22[456] + src22[457] + src22[458] + src22[459] + src22[460] + src22[461] + src22[462] + src22[463] + src22[464] + src22[465] + src22[466] + src22[467] + src22[468] + src22[469] + src22[470] + src22[471] + src22[472] + src22[473] + src22[474] + src22[475] + src22[476] + src22[477] + src22[478] + src22[479] + src22[480] + src22[481] + src22[482] + src22[483] + src22[484] + src22[485])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255] + src23[256] + src23[257] + src23[258] + src23[259] + src23[260] + src23[261] + src23[262] + src23[263] + src23[264] + src23[265] + src23[266] + src23[267] + src23[268] + src23[269] + src23[270] + src23[271] + src23[272] + src23[273] + src23[274] + src23[275] + src23[276] + src23[277] + src23[278] + src23[279] + src23[280] + src23[281] + src23[282] + src23[283] + src23[284] + src23[285] + src23[286] + src23[287] + src23[288] + src23[289] + src23[290] + src23[291] + src23[292] + src23[293] + src23[294] + src23[295] + src23[296] + src23[297] + src23[298] + src23[299] + src23[300] + src23[301] + src23[302] + src23[303] + src23[304] + src23[305] + src23[306] + src23[307] + src23[308] + src23[309] + src23[310] + src23[311] + src23[312] + src23[313] + src23[314] + src23[315] + src23[316] + src23[317] + src23[318] + src23[319] + src23[320] + src23[321] + src23[322] + src23[323] + src23[324] + src23[325] + src23[326] + src23[327] + src23[328] + src23[329] + src23[330] + src23[331] + src23[332] + src23[333] + src23[334] + src23[335] + src23[336] + src23[337] + src23[338] + src23[339] + src23[340] + src23[341] + src23[342] + src23[343] + src23[344] + src23[345] + src23[346] + src23[347] + src23[348] + src23[349] + src23[350] + src23[351] + src23[352] + src23[353] + src23[354] + src23[355] + src23[356] + src23[357] + src23[358] + src23[359] + src23[360] + src23[361] + src23[362] + src23[363] + src23[364] + src23[365] + src23[366] + src23[367] + src23[368] + src23[369] + src23[370] + src23[371] + src23[372] + src23[373] + src23[374] + src23[375] + src23[376] + src23[377] + src23[378] + src23[379] + src23[380] + src23[381] + src23[382] + src23[383] + src23[384] + src23[385] + src23[386] + src23[387] + src23[388] + src23[389] + src23[390] + src23[391] + src23[392] + src23[393] + src23[394] + src23[395] + src23[396] + src23[397] + src23[398] + src23[399] + src23[400] + src23[401] + src23[402] + src23[403] + src23[404] + src23[405] + src23[406] + src23[407] + src23[408] + src23[409] + src23[410] + src23[411] + src23[412] + src23[413] + src23[414] + src23[415] + src23[416] + src23[417] + src23[418] + src23[419] + src23[420] + src23[421] + src23[422] + src23[423] + src23[424] + src23[425] + src23[426] + src23[427] + src23[428] + src23[429] + src23[430] + src23[431] + src23[432] + src23[433] + src23[434] + src23[435] + src23[436] + src23[437] + src23[438] + src23[439] + src23[440] + src23[441] + src23[442] + src23[443] + src23[444] + src23[445] + src23[446] + src23[447] + src23[448] + src23[449] + src23[450] + src23[451] + src23[452] + src23[453] + src23[454] + src23[455] + src23[456] + src23[457] + src23[458] + src23[459] + src23[460] + src23[461] + src23[462] + src23[463] + src23[464] + src23[465] + src23[466] + src23[467] + src23[468] + src23[469] + src23[470] + src23[471] + src23[472] + src23[473] + src23[474] + src23[475] + src23[476] + src23[477] + src23[478] + src23[479] + src23[480] + src23[481] + src23[482] + src23[483] + src23[484] + src23[485])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255] + src24[256] + src24[257] + src24[258] + src24[259] + src24[260] + src24[261] + src24[262] + src24[263] + src24[264] + src24[265] + src24[266] + src24[267] + src24[268] + src24[269] + src24[270] + src24[271] + src24[272] + src24[273] + src24[274] + src24[275] + src24[276] + src24[277] + src24[278] + src24[279] + src24[280] + src24[281] + src24[282] + src24[283] + src24[284] + src24[285] + src24[286] + src24[287] + src24[288] + src24[289] + src24[290] + src24[291] + src24[292] + src24[293] + src24[294] + src24[295] + src24[296] + src24[297] + src24[298] + src24[299] + src24[300] + src24[301] + src24[302] + src24[303] + src24[304] + src24[305] + src24[306] + src24[307] + src24[308] + src24[309] + src24[310] + src24[311] + src24[312] + src24[313] + src24[314] + src24[315] + src24[316] + src24[317] + src24[318] + src24[319] + src24[320] + src24[321] + src24[322] + src24[323] + src24[324] + src24[325] + src24[326] + src24[327] + src24[328] + src24[329] + src24[330] + src24[331] + src24[332] + src24[333] + src24[334] + src24[335] + src24[336] + src24[337] + src24[338] + src24[339] + src24[340] + src24[341] + src24[342] + src24[343] + src24[344] + src24[345] + src24[346] + src24[347] + src24[348] + src24[349] + src24[350] + src24[351] + src24[352] + src24[353] + src24[354] + src24[355] + src24[356] + src24[357] + src24[358] + src24[359] + src24[360] + src24[361] + src24[362] + src24[363] + src24[364] + src24[365] + src24[366] + src24[367] + src24[368] + src24[369] + src24[370] + src24[371] + src24[372] + src24[373] + src24[374] + src24[375] + src24[376] + src24[377] + src24[378] + src24[379] + src24[380] + src24[381] + src24[382] + src24[383] + src24[384] + src24[385] + src24[386] + src24[387] + src24[388] + src24[389] + src24[390] + src24[391] + src24[392] + src24[393] + src24[394] + src24[395] + src24[396] + src24[397] + src24[398] + src24[399] + src24[400] + src24[401] + src24[402] + src24[403] + src24[404] + src24[405] + src24[406] + src24[407] + src24[408] + src24[409] + src24[410] + src24[411] + src24[412] + src24[413] + src24[414] + src24[415] + src24[416] + src24[417] + src24[418] + src24[419] + src24[420] + src24[421] + src24[422] + src24[423] + src24[424] + src24[425] + src24[426] + src24[427] + src24[428] + src24[429] + src24[430] + src24[431] + src24[432] + src24[433] + src24[434] + src24[435] + src24[436] + src24[437] + src24[438] + src24[439] + src24[440] + src24[441] + src24[442] + src24[443] + src24[444] + src24[445] + src24[446] + src24[447] + src24[448] + src24[449] + src24[450] + src24[451] + src24[452] + src24[453] + src24[454] + src24[455] + src24[456] + src24[457] + src24[458] + src24[459] + src24[460] + src24[461] + src24[462] + src24[463] + src24[464] + src24[465] + src24[466] + src24[467] + src24[468] + src24[469] + src24[470] + src24[471] + src24[472] + src24[473] + src24[474] + src24[475] + src24[476] + src24[477] + src24[478] + src24[479] + src24[480] + src24[481] + src24[482] + src24[483] + src24[484] + src24[485])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255] + src25[256] + src25[257] + src25[258] + src25[259] + src25[260] + src25[261] + src25[262] + src25[263] + src25[264] + src25[265] + src25[266] + src25[267] + src25[268] + src25[269] + src25[270] + src25[271] + src25[272] + src25[273] + src25[274] + src25[275] + src25[276] + src25[277] + src25[278] + src25[279] + src25[280] + src25[281] + src25[282] + src25[283] + src25[284] + src25[285] + src25[286] + src25[287] + src25[288] + src25[289] + src25[290] + src25[291] + src25[292] + src25[293] + src25[294] + src25[295] + src25[296] + src25[297] + src25[298] + src25[299] + src25[300] + src25[301] + src25[302] + src25[303] + src25[304] + src25[305] + src25[306] + src25[307] + src25[308] + src25[309] + src25[310] + src25[311] + src25[312] + src25[313] + src25[314] + src25[315] + src25[316] + src25[317] + src25[318] + src25[319] + src25[320] + src25[321] + src25[322] + src25[323] + src25[324] + src25[325] + src25[326] + src25[327] + src25[328] + src25[329] + src25[330] + src25[331] + src25[332] + src25[333] + src25[334] + src25[335] + src25[336] + src25[337] + src25[338] + src25[339] + src25[340] + src25[341] + src25[342] + src25[343] + src25[344] + src25[345] + src25[346] + src25[347] + src25[348] + src25[349] + src25[350] + src25[351] + src25[352] + src25[353] + src25[354] + src25[355] + src25[356] + src25[357] + src25[358] + src25[359] + src25[360] + src25[361] + src25[362] + src25[363] + src25[364] + src25[365] + src25[366] + src25[367] + src25[368] + src25[369] + src25[370] + src25[371] + src25[372] + src25[373] + src25[374] + src25[375] + src25[376] + src25[377] + src25[378] + src25[379] + src25[380] + src25[381] + src25[382] + src25[383] + src25[384] + src25[385] + src25[386] + src25[387] + src25[388] + src25[389] + src25[390] + src25[391] + src25[392] + src25[393] + src25[394] + src25[395] + src25[396] + src25[397] + src25[398] + src25[399] + src25[400] + src25[401] + src25[402] + src25[403] + src25[404] + src25[405] + src25[406] + src25[407] + src25[408] + src25[409] + src25[410] + src25[411] + src25[412] + src25[413] + src25[414] + src25[415] + src25[416] + src25[417] + src25[418] + src25[419] + src25[420] + src25[421] + src25[422] + src25[423] + src25[424] + src25[425] + src25[426] + src25[427] + src25[428] + src25[429] + src25[430] + src25[431] + src25[432] + src25[433] + src25[434] + src25[435] + src25[436] + src25[437] + src25[438] + src25[439] + src25[440] + src25[441] + src25[442] + src25[443] + src25[444] + src25[445] + src25[446] + src25[447] + src25[448] + src25[449] + src25[450] + src25[451] + src25[452] + src25[453] + src25[454] + src25[455] + src25[456] + src25[457] + src25[458] + src25[459] + src25[460] + src25[461] + src25[462] + src25[463] + src25[464] + src25[465] + src25[466] + src25[467] + src25[468] + src25[469] + src25[470] + src25[471] + src25[472] + src25[473] + src25[474] + src25[475] + src25[476] + src25[477] + src25[478] + src25[479] + src25[480] + src25[481] + src25[482] + src25[483] + src25[484] + src25[485])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255] + src26[256] + src26[257] + src26[258] + src26[259] + src26[260] + src26[261] + src26[262] + src26[263] + src26[264] + src26[265] + src26[266] + src26[267] + src26[268] + src26[269] + src26[270] + src26[271] + src26[272] + src26[273] + src26[274] + src26[275] + src26[276] + src26[277] + src26[278] + src26[279] + src26[280] + src26[281] + src26[282] + src26[283] + src26[284] + src26[285] + src26[286] + src26[287] + src26[288] + src26[289] + src26[290] + src26[291] + src26[292] + src26[293] + src26[294] + src26[295] + src26[296] + src26[297] + src26[298] + src26[299] + src26[300] + src26[301] + src26[302] + src26[303] + src26[304] + src26[305] + src26[306] + src26[307] + src26[308] + src26[309] + src26[310] + src26[311] + src26[312] + src26[313] + src26[314] + src26[315] + src26[316] + src26[317] + src26[318] + src26[319] + src26[320] + src26[321] + src26[322] + src26[323] + src26[324] + src26[325] + src26[326] + src26[327] + src26[328] + src26[329] + src26[330] + src26[331] + src26[332] + src26[333] + src26[334] + src26[335] + src26[336] + src26[337] + src26[338] + src26[339] + src26[340] + src26[341] + src26[342] + src26[343] + src26[344] + src26[345] + src26[346] + src26[347] + src26[348] + src26[349] + src26[350] + src26[351] + src26[352] + src26[353] + src26[354] + src26[355] + src26[356] + src26[357] + src26[358] + src26[359] + src26[360] + src26[361] + src26[362] + src26[363] + src26[364] + src26[365] + src26[366] + src26[367] + src26[368] + src26[369] + src26[370] + src26[371] + src26[372] + src26[373] + src26[374] + src26[375] + src26[376] + src26[377] + src26[378] + src26[379] + src26[380] + src26[381] + src26[382] + src26[383] + src26[384] + src26[385] + src26[386] + src26[387] + src26[388] + src26[389] + src26[390] + src26[391] + src26[392] + src26[393] + src26[394] + src26[395] + src26[396] + src26[397] + src26[398] + src26[399] + src26[400] + src26[401] + src26[402] + src26[403] + src26[404] + src26[405] + src26[406] + src26[407] + src26[408] + src26[409] + src26[410] + src26[411] + src26[412] + src26[413] + src26[414] + src26[415] + src26[416] + src26[417] + src26[418] + src26[419] + src26[420] + src26[421] + src26[422] + src26[423] + src26[424] + src26[425] + src26[426] + src26[427] + src26[428] + src26[429] + src26[430] + src26[431] + src26[432] + src26[433] + src26[434] + src26[435] + src26[436] + src26[437] + src26[438] + src26[439] + src26[440] + src26[441] + src26[442] + src26[443] + src26[444] + src26[445] + src26[446] + src26[447] + src26[448] + src26[449] + src26[450] + src26[451] + src26[452] + src26[453] + src26[454] + src26[455] + src26[456] + src26[457] + src26[458] + src26[459] + src26[460] + src26[461] + src26[462] + src26[463] + src26[464] + src26[465] + src26[466] + src26[467] + src26[468] + src26[469] + src26[470] + src26[471] + src26[472] + src26[473] + src26[474] + src26[475] + src26[476] + src26[477] + src26[478] + src26[479] + src26[480] + src26[481] + src26[482] + src26[483] + src26[484] + src26[485])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255] + src27[256] + src27[257] + src27[258] + src27[259] + src27[260] + src27[261] + src27[262] + src27[263] + src27[264] + src27[265] + src27[266] + src27[267] + src27[268] + src27[269] + src27[270] + src27[271] + src27[272] + src27[273] + src27[274] + src27[275] + src27[276] + src27[277] + src27[278] + src27[279] + src27[280] + src27[281] + src27[282] + src27[283] + src27[284] + src27[285] + src27[286] + src27[287] + src27[288] + src27[289] + src27[290] + src27[291] + src27[292] + src27[293] + src27[294] + src27[295] + src27[296] + src27[297] + src27[298] + src27[299] + src27[300] + src27[301] + src27[302] + src27[303] + src27[304] + src27[305] + src27[306] + src27[307] + src27[308] + src27[309] + src27[310] + src27[311] + src27[312] + src27[313] + src27[314] + src27[315] + src27[316] + src27[317] + src27[318] + src27[319] + src27[320] + src27[321] + src27[322] + src27[323] + src27[324] + src27[325] + src27[326] + src27[327] + src27[328] + src27[329] + src27[330] + src27[331] + src27[332] + src27[333] + src27[334] + src27[335] + src27[336] + src27[337] + src27[338] + src27[339] + src27[340] + src27[341] + src27[342] + src27[343] + src27[344] + src27[345] + src27[346] + src27[347] + src27[348] + src27[349] + src27[350] + src27[351] + src27[352] + src27[353] + src27[354] + src27[355] + src27[356] + src27[357] + src27[358] + src27[359] + src27[360] + src27[361] + src27[362] + src27[363] + src27[364] + src27[365] + src27[366] + src27[367] + src27[368] + src27[369] + src27[370] + src27[371] + src27[372] + src27[373] + src27[374] + src27[375] + src27[376] + src27[377] + src27[378] + src27[379] + src27[380] + src27[381] + src27[382] + src27[383] + src27[384] + src27[385] + src27[386] + src27[387] + src27[388] + src27[389] + src27[390] + src27[391] + src27[392] + src27[393] + src27[394] + src27[395] + src27[396] + src27[397] + src27[398] + src27[399] + src27[400] + src27[401] + src27[402] + src27[403] + src27[404] + src27[405] + src27[406] + src27[407] + src27[408] + src27[409] + src27[410] + src27[411] + src27[412] + src27[413] + src27[414] + src27[415] + src27[416] + src27[417] + src27[418] + src27[419] + src27[420] + src27[421] + src27[422] + src27[423] + src27[424] + src27[425] + src27[426] + src27[427] + src27[428] + src27[429] + src27[430] + src27[431] + src27[432] + src27[433] + src27[434] + src27[435] + src27[436] + src27[437] + src27[438] + src27[439] + src27[440] + src27[441] + src27[442] + src27[443] + src27[444] + src27[445] + src27[446] + src27[447] + src27[448] + src27[449] + src27[450] + src27[451] + src27[452] + src27[453] + src27[454] + src27[455] + src27[456] + src27[457] + src27[458] + src27[459] + src27[460] + src27[461] + src27[462] + src27[463] + src27[464] + src27[465] + src27[466] + src27[467] + src27[468] + src27[469] + src27[470] + src27[471] + src27[472] + src27[473] + src27[474] + src27[475] + src27[476] + src27[477] + src27[478] + src27[479] + src27[480] + src27[481] + src27[482] + src27[483] + src27[484] + src27[485])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255] + src28[256] + src28[257] + src28[258] + src28[259] + src28[260] + src28[261] + src28[262] + src28[263] + src28[264] + src28[265] + src28[266] + src28[267] + src28[268] + src28[269] + src28[270] + src28[271] + src28[272] + src28[273] + src28[274] + src28[275] + src28[276] + src28[277] + src28[278] + src28[279] + src28[280] + src28[281] + src28[282] + src28[283] + src28[284] + src28[285] + src28[286] + src28[287] + src28[288] + src28[289] + src28[290] + src28[291] + src28[292] + src28[293] + src28[294] + src28[295] + src28[296] + src28[297] + src28[298] + src28[299] + src28[300] + src28[301] + src28[302] + src28[303] + src28[304] + src28[305] + src28[306] + src28[307] + src28[308] + src28[309] + src28[310] + src28[311] + src28[312] + src28[313] + src28[314] + src28[315] + src28[316] + src28[317] + src28[318] + src28[319] + src28[320] + src28[321] + src28[322] + src28[323] + src28[324] + src28[325] + src28[326] + src28[327] + src28[328] + src28[329] + src28[330] + src28[331] + src28[332] + src28[333] + src28[334] + src28[335] + src28[336] + src28[337] + src28[338] + src28[339] + src28[340] + src28[341] + src28[342] + src28[343] + src28[344] + src28[345] + src28[346] + src28[347] + src28[348] + src28[349] + src28[350] + src28[351] + src28[352] + src28[353] + src28[354] + src28[355] + src28[356] + src28[357] + src28[358] + src28[359] + src28[360] + src28[361] + src28[362] + src28[363] + src28[364] + src28[365] + src28[366] + src28[367] + src28[368] + src28[369] + src28[370] + src28[371] + src28[372] + src28[373] + src28[374] + src28[375] + src28[376] + src28[377] + src28[378] + src28[379] + src28[380] + src28[381] + src28[382] + src28[383] + src28[384] + src28[385] + src28[386] + src28[387] + src28[388] + src28[389] + src28[390] + src28[391] + src28[392] + src28[393] + src28[394] + src28[395] + src28[396] + src28[397] + src28[398] + src28[399] + src28[400] + src28[401] + src28[402] + src28[403] + src28[404] + src28[405] + src28[406] + src28[407] + src28[408] + src28[409] + src28[410] + src28[411] + src28[412] + src28[413] + src28[414] + src28[415] + src28[416] + src28[417] + src28[418] + src28[419] + src28[420] + src28[421] + src28[422] + src28[423] + src28[424] + src28[425] + src28[426] + src28[427] + src28[428] + src28[429] + src28[430] + src28[431] + src28[432] + src28[433] + src28[434] + src28[435] + src28[436] + src28[437] + src28[438] + src28[439] + src28[440] + src28[441] + src28[442] + src28[443] + src28[444] + src28[445] + src28[446] + src28[447] + src28[448] + src28[449] + src28[450] + src28[451] + src28[452] + src28[453] + src28[454] + src28[455] + src28[456] + src28[457] + src28[458] + src28[459] + src28[460] + src28[461] + src28[462] + src28[463] + src28[464] + src28[465] + src28[466] + src28[467] + src28[468] + src28[469] + src28[470] + src28[471] + src28[472] + src28[473] + src28[474] + src28[475] + src28[476] + src28[477] + src28[478] + src28[479] + src28[480] + src28[481] + src28[482] + src28[483] + src28[484] + src28[485])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255] + src29[256] + src29[257] + src29[258] + src29[259] + src29[260] + src29[261] + src29[262] + src29[263] + src29[264] + src29[265] + src29[266] + src29[267] + src29[268] + src29[269] + src29[270] + src29[271] + src29[272] + src29[273] + src29[274] + src29[275] + src29[276] + src29[277] + src29[278] + src29[279] + src29[280] + src29[281] + src29[282] + src29[283] + src29[284] + src29[285] + src29[286] + src29[287] + src29[288] + src29[289] + src29[290] + src29[291] + src29[292] + src29[293] + src29[294] + src29[295] + src29[296] + src29[297] + src29[298] + src29[299] + src29[300] + src29[301] + src29[302] + src29[303] + src29[304] + src29[305] + src29[306] + src29[307] + src29[308] + src29[309] + src29[310] + src29[311] + src29[312] + src29[313] + src29[314] + src29[315] + src29[316] + src29[317] + src29[318] + src29[319] + src29[320] + src29[321] + src29[322] + src29[323] + src29[324] + src29[325] + src29[326] + src29[327] + src29[328] + src29[329] + src29[330] + src29[331] + src29[332] + src29[333] + src29[334] + src29[335] + src29[336] + src29[337] + src29[338] + src29[339] + src29[340] + src29[341] + src29[342] + src29[343] + src29[344] + src29[345] + src29[346] + src29[347] + src29[348] + src29[349] + src29[350] + src29[351] + src29[352] + src29[353] + src29[354] + src29[355] + src29[356] + src29[357] + src29[358] + src29[359] + src29[360] + src29[361] + src29[362] + src29[363] + src29[364] + src29[365] + src29[366] + src29[367] + src29[368] + src29[369] + src29[370] + src29[371] + src29[372] + src29[373] + src29[374] + src29[375] + src29[376] + src29[377] + src29[378] + src29[379] + src29[380] + src29[381] + src29[382] + src29[383] + src29[384] + src29[385] + src29[386] + src29[387] + src29[388] + src29[389] + src29[390] + src29[391] + src29[392] + src29[393] + src29[394] + src29[395] + src29[396] + src29[397] + src29[398] + src29[399] + src29[400] + src29[401] + src29[402] + src29[403] + src29[404] + src29[405] + src29[406] + src29[407] + src29[408] + src29[409] + src29[410] + src29[411] + src29[412] + src29[413] + src29[414] + src29[415] + src29[416] + src29[417] + src29[418] + src29[419] + src29[420] + src29[421] + src29[422] + src29[423] + src29[424] + src29[425] + src29[426] + src29[427] + src29[428] + src29[429] + src29[430] + src29[431] + src29[432] + src29[433] + src29[434] + src29[435] + src29[436] + src29[437] + src29[438] + src29[439] + src29[440] + src29[441] + src29[442] + src29[443] + src29[444] + src29[445] + src29[446] + src29[447] + src29[448] + src29[449] + src29[450] + src29[451] + src29[452] + src29[453] + src29[454] + src29[455] + src29[456] + src29[457] + src29[458] + src29[459] + src29[460] + src29[461] + src29[462] + src29[463] + src29[464] + src29[465] + src29[466] + src29[467] + src29[468] + src29[469] + src29[470] + src29[471] + src29[472] + src29[473] + src29[474] + src29[475] + src29[476] + src29[477] + src29[478] + src29[479] + src29[480] + src29[481] + src29[482] + src29[483] + src29[484] + src29[485])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255] + src30[256] + src30[257] + src30[258] + src30[259] + src30[260] + src30[261] + src30[262] + src30[263] + src30[264] + src30[265] + src30[266] + src30[267] + src30[268] + src30[269] + src30[270] + src30[271] + src30[272] + src30[273] + src30[274] + src30[275] + src30[276] + src30[277] + src30[278] + src30[279] + src30[280] + src30[281] + src30[282] + src30[283] + src30[284] + src30[285] + src30[286] + src30[287] + src30[288] + src30[289] + src30[290] + src30[291] + src30[292] + src30[293] + src30[294] + src30[295] + src30[296] + src30[297] + src30[298] + src30[299] + src30[300] + src30[301] + src30[302] + src30[303] + src30[304] + src30[305] + src30[306] + src30[307] + src30[308] + src30[309] + src30[310] + src30[311] + src30[312] + src30[313] + src30[314] + src30[315] + src30[316] + src30[317] + src30[318] + src30[319] + src30[320] + src30[321] + src30[322] + src30[323] + src30[324] + src30[325] + src30[326] + src30[327] + src30[328] + src30[329] + src30[330] + src30[331] + src30[332] + src30[333] + src30[334] + src30[335] + src30[336] + src30[337] + src30[338] + src30[339] + src30[340] + src30[341] + src30[342] + src30[343] + src30[344] + src30[345] + src30[346] + src30[347] + src30[348] + src30[349] + src30[350] + src30[351] + src30[352] + src30[353] + src30[354] + src30[355] + src30[356] + src30[357] + src30[358] + src30[359] + src30[360] + src30[361] + src30[362] + src30[363] + src30[364] + src30[365] + src30[366] + src30[367] + src30[368] + src30[369] + src30[370] + src30[371] + src30[372] + src30[373] + src30[374] + src30[375] + src30[376] + src30[377] + src30[378] + src30[379] + src30[380] + src30[381] + src30[382] + src30[383] + src30[384] + src30[385] + src30[386] + src30[387] + src30[388] + src30[389] + src30[390] + src30[391] + src30[392] + src30[393] + src30[394] + src30[395] + src30[396] + src30[397] + src30[398] + src30[399] + src30[400] + src30[401] + src30[402] + src30[403] + src30[404] + src30[405] + src30[406] + src30[407] + src30[408] + src30[409] + src30[410] + src30[411] + src30[412] + src30[413] + src30[414] + src30[415] + src30[416] + src30[417] + src30[418] + src30[419] + src30[420] + src30[421] + src30[422] + src30[423] + src30[424] + src30[425] + src30[426] + src30[427] + src30[428] + src30[429] + src30[430] + src30[431] + src30[432] + src30[433] + src30[434] + src30[435] + src30[436] + src30[437] + src30[438] + src30[439] + src30[440] + src30[441] + src30[442] + src30[443] + src30[444] + src30[445] + src30[446] + src30[447] + src30[448] + src30[449] + src30[450] + src30[451] + src30[452] + src30[453] + src30[454] + src30[455] + src30[456] + src30[457] + src30[458] + src30[459] + src30[460] + src30[461] + src30[462] + src30[463] + src30[464] + src30[465] + src30[466] + src30[467] + src30[468] + src30[469] + src30[470] + src30[471] + src30[472] + src30[473] + src30[474] + src30[475] + src30[476] + src30[477] + src30[478] + src30[479] + src30[480] + src30[481] + src30[482] + src30[483] + src30[484] + src30[485])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255] + src31[256] + src31[257] + src31[258] + src31[259] + src31[260] + src31[261] + src31[262] + src31[263] + src31[264] + src31[265] + src31[266] + src31[267] + src31[268] + src31[269] + src31[270] + src31[271] + src31[272] + src31[273] + src31[274] + src31[275] + src31[276] + src31[277] + src31[278] + src31[279] + src31[280] + src31[281] + src31[282] + src31[283] + src31[284] + src31[285] + src31[286] + src31[287] + src31[288] + src31[289] + src31[290] + src31[291] + src31[292] + src31[293] + src31[294] + src31[295] + src31[296] + src31[297] + src31[298] + src31[299] + src31[300] + src31[301] + src31[302] + src31[303] + src31[304] + src31[305] + src31[306] + src31[307] + src31[308] + src31[309] + src31[310] + src31[311] + src31[312] + src31[313] + src31[314] + src31[315] + src31[316] + src31[317] + src31[318] + src31[319] + src31[320] + src31[321] + src31[322] + src31[323] + src31[324] + src31[325] + src31[326] + src31[327] + src31[328] + src31[329] + src31[330] + src31[331] + src31[332] + src31[333] + src31[334] + src31[335] + src31[336] + src31[337] + src31[338] + src31[339] + src31[340] + src31[341] + src31[342] + src31[343] + src31[344] + src31[345] + src31[346] + src31[347] + src31[348] + src31[349] + src31[350] + src31[351] + src31[352] + src31[353] + src31[354] + src31[355] + src31[356] + src31[357] + src31[358] + src31[359] + src31[360] + src31[361] + src31[362] + src31[363] + src31[364] + src31[365] + src31[366] + src31[367] + src31[368] + src31[369] + src31[370] + src31[371] + src31[372] + src31[373] + src31[374] + src31[375] + src31[376] + src31[377] + src31[378] + src31[379] + src31[380] + src31[381] + src31[382] + src31[383] + src31[384] + src31[385] + src31[386] + src31[387] + src31[388] + src31[389] + src31[390] + src31[391] + src31[392] + src31[393] + src31[394] + src31[395] + src31[396] + src31[397] + src31[398] + src31[399] + src31[400] + src31[401] + src31[402] + src31[403] + src31[404] + src31[405] + src31[406] + src31[407] + src31[408] + src31[409] + src31[410] + src31[411] + src31[412] + src31[413] + src31[414] + src31[415] + src31[416] + src31[417] + src31[418] + src31[419] + src31[420] + src31[421] + src31[422] + src31[423] + src31[424] + src31[425] + src31[426] + src31[427] + src31[428] + src31[429] + src31[430] + src31[431] + src31[432] + src31[433] + src31[434] + src31[435] + src31[436] + src31[437] + src31[438] + src31[439] + src31[440] + src31[441] + src31[442] + src31[443] + src31[444] + src31[445] + src31[446] + src31[447] + src31[448] + src31[449] + src31[450] + src31[451] + src31[452] + src31[453] + src31[454] + src31[455] + src31[456] + src31[457] + src31[458] + src31[459] + src31[460] + src31[461] + src31[462] + src31[463] + src31[464] + src31[465] + src31[466] + src31[467] + src31[468] + src31[469] + src31[470] + src31[471] + src31[472] + src31[473] + src31[474] + src31[475] + src31[476] + src31[477] + src31[478] + src31[479] + src31[480] + src31[481] + src31[482] + src31[483] + src31[484] + src31[485])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbe1dffa3697a237b89c43b0bbf8cc438c0cf3cf23ab9591a6fbed7e2e84eca2a8ca5a0ee72fc70083f41b86c5697bac7fa41b3842f5f97cb150dab6e59c0fdcd21bc449d5313670f52114cbc39afdc8a1becad9b1423dddc959c6fa61602eaf26a8b84a23ef257ccad9e8b0853a923e784dc70381f59727ba59d2ee213ff732149864e4c9d9a3e0e63977c678a8cdf9e1646a9087b83706046b9d55a8c8b570633f6b50afe577c28ff7840e0ec905b2176f6f5fb51e80956cb0945cfe19b02abb32d14d65011958f8365fb78c2de21e61f8fe948365227101aedcb5ebc5a6204453be493e8194ec97439b1e349a2bcd201ecf4764e253d6c3c32ad4e24d1639e184289411b27a99647e8fe62c2a940eba05da14e830f0e87cf4232b808ab3f0522cde4471a1e8e69b37eb95ff70689042f34e719114e94db4a54c82504d09ee7ad939ecf32413029ca9f9308e7510230fff53900ab20b07fcae16d4cc2657891071fda45d16a73edb591460591e39c6d60e81c1421b3a5329c7ce2669d0914f2a7e56dd6d2dde52ffec54e1757c5f3d4b392a0231f2457b77e13313998a2be3ed18b8920c4cc89183647590bf72ead42b4e164e8d099523258dcf15c186555f5f47c71deee4ea0697e8eb7bf643a0f1a30d47e769f4efab2a10cf8ba0ebde69cf0f2110b9c132f73817fb6ec7e7d66c870a724fc540f6231fdc91a5ca6a752c751bf461468cc7dd68c220a0026288990c0f318dfa6b7cf25481328c5200bce70a076b8fbe33d6f923f89fda586c3ca27c0f5740bf200d1099bd413567f409a80fa9ee6da63dcf95d1f6b1d20b723fa7c09b9a5147eb51a895fbd5d5228a1bb3cded962eac5837da010a8baeb5d465e84e3d03c07d09b58a60739b8257185b96c86012b5453aa6a32d9af32479b611fa6e5e92bdd4c8dc6e844259c3d224f98d03bf661a0af2864f54f3ed03dbd7903d9a302bcc925c223479be3fffcc949401b768b76dcb195c386bbd94bf6a4fd8d30a0096c404b64c7093b53ba3ab041c633397d45828d83bc0c57ffcbd881c3c1217d2b8d088d14c352d3de1289c52ecdb0f3f6b8684d2ccc2e6122f7ebd5fec0cd9c7b198295e926434a5a4e30154bc0999ccb0895deaca9459c4a8df586da5eedb8bc353ea209db0741359d3b061f166d10fad39af0d2c91c3e732eda37ef2007173828c117779b6abb7b4ca868b2da98fea3c9f43ee70c2714ebc0a1457069f7fe03c51304eace60ff0f8d0ea86bdeb7bf22ae55f85674ff0024f1a84e585427febf55e0a14677a245ec060c193f74a324cf8321203229e2b839c1ae7c67e4f63908e64526e94ed8d69d2b61a16ac808b131ab3e609146a8c13df5a49525bf33becb05c0ae533055d367686e5288c4eccc5347a3491cc8e9925d9071a0ad8280f28df313dbae3a3d8b8baacfb16e27d61aa18fa457a30fc2eba5fe68f66fd76cda75a8bcb7af9a92a0eeee550398899af37061975ef999cb2ed24ddb07a9deb4dbf6db3cc9d017785f0608b998a506ff379257f3f39c8ccf6e4b7cb2c13eac237551d9db618682e6d5eda43320100eade9107c7f5c4c8bba580cc6ececa9aa2626efbeeddd9f9d80ae18f860c5d108aadbbadc2e1b50d55fa18e635fb3d6f6b6309c98ab5fb96f7f5dcabfa771674dfc89749db07c8c41bb13e75ec07491669a660c18dc182ddb7d546570c7221f88e535861b02282280a0d9e4a8a6d755b5d0b7f053089df15327579670981ae9441cb22fb14528b56d0e4b63baab8074a3f7cead9556c14fe2211384307d7593fb39b52597a9465e94ddcea4c6e63f489547752f1fd9bc84a5696aae9a107797102778fb102f0ac9d8cce56d2a8972628c669352cf4f7ce00fd14b568048653f3687d7cd10cd7b266a41e64e331f3f3bafdae3ac4962090935920eaa7d955772038fec55cc84691dfdf66199761da58682c40d96c159f06cf7a0604f7dbfc58bcd1569e26935e0aa4bf26b6d8000ef3aa887c7f64aded112584edbdfa30a7522302ef9912ef8627d5a571cccdbdbc4b729122100fbc3af02ee42f4c94c6e1dcaf6a4034f4539e6c356bb49b6918258cfbf3c468b9da7c4b832bbfee582f773016b318134454c2ce49675f5e3685444173466ee34fb6ac649493e8c529d90c4f2ad0479fec12a627ba402cb65f64d27d798c3a77583ec587fb6451d7eef960e71f6a82b323528349c705fabeb5bbbda3766f693f2a4d13bedad9c15fb8ab6ef12b1eacc668dad35f5039b7239e3c57e60131b2cd7dd5b6f1055eb66a5ff4c1f1307473eb07c17332e2326b5a55c7b8dcbbc20b0ff149b7a15f95eede770d738be5c55f264e20fe5b169eabd46685201a7bf8a8b61b9139fd397100c58833919e956f13c20ed78fd4538c3a5c0765242fd6b8e6b59c8d82945eaf4025371af2a8de9fc6c560e1d0a993a4f93ac596b8d063a8fcc739a1438a7d54ee63cec687f8b482d45e8c573f8335f74dc6aafd8ec449b6d1f9ad41856130b73e24386750935864c90c105fe8b3f0a40a1ff01b19bdb1096e4e1f8a707847b8b1807dd0fbdfa9ae6b4383e57fc82d35241db1e0ccb95f4d5aab8a07e60389d54c13307c4345b148d581dbe3cbc450de4f566df7d56899bd3fc61660dca54bd70f0ac459fa6deb3f4ffce9b0a3c9fe3bb2708e6474fe4ba5e046d131b7e021c2e6a8413ad695de8ff5836889d99b041c2616c9ef72fb41b04498ea7909984f3b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6e7164006fef69371cde2f9cf3d732c4d6d1e4c8e21456bc17babf0332b82e791610194a1a8c3dae39931fe181d08b948dcd9e123f96c42459c32dda32150d4e6f6e36f6096cd45e45237869214da3d015d8e7e7dc8d1ca48062a59e526f7215362f48fd89b4286bf1a74ef4ec2ece89b7cd0e50468556e6ad38fe3e482dd712b69b9cdcd58c9aab0d337c6493b3aad120ce2e454b41a8238918a9ebf35992002a17269c0c8f527f0481db42582f4a47e3d103d49b015033b493bff9ea44aa891b4e88d3a495ede995ce42c99bd0431650830ba1e6b3cd7723f1d785fc3ff8e6bba1c9942fdc799cbb8144d8f77acba0a0c199136dd59a817dec1411d3866497c8dfa64b0242fffde3f987ddebd94995cc2c17549cf5aa6c957d7fb060794e26c0118a615046e413bdf63ccb0ee1f63cc7e5ac3f249e30e27a53e01eb1c1f559171297c2d17ef17796756f1d99974b46d5a8b4a8383a3015b56af0c8373c83da0dc8758cc24b0e695f80aee996d573c0531562ad1263df93460cc5db9c90192f135a061d1701a89adf1f0108880cea04dd52efc71524425ff21019011b59bdcc53a32b64a643111b28a69b61ad2cbb7320378aaeb17111bf08b6d7f159f7ef58388be785992adc1d95978b24c8463b85da1aadc81db87c048996a596b482aae54c27122d04454c07dbf072e25d99ee1f30a2027126e6f5d128f8c8f0369486edcbce3c33ac4f36756de8b2c6165ff57c135e5ac300877f05934d82b66689c53ff085ab75972c39d3f96b1e2fc3c6b94c038154835fbdb8ed14d0b373202e3fc80ad9b862cddfdda094ce59e6978a728a4f1bd8e18de4bb618f8d9c96e4560e0c45c1cf81f034371ad85639f360b6d07389592ea992f3acf79fed41c6bd9bf5104e6a5d1123f348b123b6ce8c1ba7aeb14a90b62f6b3df5e32d877577e15696ba7a5f91555ddb4f225c6318dd32a2f92ab78a2b3e420e546079b42af50d3d8cec86601563678056a0e0c02858e5e5d485d317e91c687aa9826e1365e6c49659ef1dc26397e7a3db20825297f3640d850205e9614e207ec0093707a2f7a2629711ceee891583a9972c2637fa2f16e541a5df4fb51ef9f6bcbe19931f7a183fa872b752cf39d65492c243eed0996dcc6f012f1e5b889c34291dc81da2daa199b5dbc4ce7b57202cfba750cd2c6e4d7d136149cf51716c6e34bd5b8dd533131612580b1075c27cdc717f3600c42afc500e313d74b8421817ebdac57c5dc6fe2fd6b125cc769b1e2c8e94579c8ad3b19452fce3eff85245b112f26b13c59fc43d1c779f92841d29c3a98a6198cbd80ed4aca1e8b6c9563cd543f059255b144aa9e397109c7704f32957d2163a9f1b654a98e70f4b088f50c66b96092bc624788d19920662f52af9a20dadf0c5d37fbce1d4515708e6e33b302681b6034089880955ac2d02d27ee99f7b0adb6aa5ece8a75746ff25442b0175c9e16caa0f8b8ccf2a0ad883ae0a83505eb28d72e5c7960ea36f1e1b3dc533f452a065cb693cc8caf6464dd7bc0c3b945b1c11071ca8b0c371a1bad25ef3d025f2eec438bedb1ea689c9f4735adb0401130b8f400c115eb6c2770be1c856a77fab7795fae233ff6575d33775dd451c63107d3028bf8b19079fd5a2a9b1b7bad34083aa83a59013aa1284d3a45f2e175da738e47c1600a4a9632c6a5a5842883d31120433535018b56a5328073887869c4dbaed6e6114846f043ce7aa32bcfd8016add74407b11e5a6e4200ad9804ee3b6ee6766eca8d43d8d744e8ab6265d5cd8ed8554c834a0b1a570f271773dc31b1d9a6c28f2bce239e97d819d8f1d2532c1ce5b34a236f0c4880d2aea2cf12ed3f56dcf5ad012a8065b7fe3ed4a1f9bf4f6c829927439bd7e31759900aef02c25066bd44a1be63ebbf1177f2152f844aec7d63a77d0b4dd989ec18f606b1adacce9cadc96c6476a08ea6117a083e9b853399641a20c9f716e68bd961eeac71db82494cc4a122229c7dddffd54862fa29030f018bc2500e16a5f0a85a8cc0b7f223d5aa269c9a0ba00eb65adc2da56b72b39ccb8d0637b642dccae004de7dc615cada266a8d0bcec1bd7d034cb42a555d945a398e31bfa8d9b21599c65060c45ef1f55c8d22f438677d21bc90710a30e27777783f645aa9c354815213ef2fa0060aff591b75ae66d045e3792a690869463317f7621391f436ef96001a8773ea6d9be236a6f1178bf826e04a2ae5ce25c644d8464f68ceccb8b13ca5401a0b99e4b9c7bfb8dbf3f0a4986b3b261d362b3aa530e4a763b1519b1b7d12d71a3dcafdffb6451a816e9814c632cb778787aa29a6a978c759d6c7d7cb069a35bb4541a381821c0dfcf1d03ccab91735b4b9b9c03dec3d08e890cdbf9c68d17dc4439cb0e0c38bf62aa481e7917dd080650264ca0547d761689d48acc1770eedee3c7830a6890dc57fa0f31a4d376d8b8393d8e2167289c2b644c4df0c83958d7b55b75f29e3afdc92b56f8eed9d87aa32ca49ae275763c6048a2b2f2784e21c1eaa9bf1ced3990ccb521639f9175607dbf384a2f257e08e039df06f12914ba076d6d30a64251e1c9bfcbd5789c7be5ba153b38ab495b910a105e53d0f124409d233a370a2c7c2c20ead9aa32d13776349d82cdbc1f5e12d4a098688e41b1ac90bd048e214ff5208544b0a6b2622e7089c3afd1fc1efd3ac1115e06b0b44624d5f6e800447fc35a4d5864c3ebdb2186df6547ad6c010b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hde102e80ca0a58959e5d37c2e085dffa9365be0a779cb94927119b690b2b8f6d9b496402595261f189579144a96734c55bcee2509c25b3ed4f38088f5b55ccb262e306bee3dc5e2df6b71454ba3ffb38ed34e04062f4e77b17027a151634b258538452c8982ac8a0e836ffbb656429a3d82db1039f65b95ed173b8b9c5cfb41e4946955ccc7c32e7fd08ba07d11bf8ee40487400965b531dfbb8959304c0abaff1a51c4d0a684a6b173255dad1cab7441d781bb185f4709daacb1b9695ab77703805964dd391f0013d441ba6f89f2e8eb1c9fb5f4b0e1c0e10a9888119e139a4c48884608c65a3660707780fb0f1ad145f048937dfb0a79171327c5439771d169d57f029bae315d7d74bd8c93e59500eb25dcd9b136a97ac4ab87ee153626874b4f65aa600f27d261366d8ed01a955e3c96c15f42818ec41e27618f4b493155b8bc41af477b2d5eacf267da5cdaf10560d76f7a5f25866bfae89374903ec860d8992b3a46c46edd22f44c4c7eed2a9b8355757b8f29c272cb67eb04c58676ec2993287a891e11e5dc52b01bbebc546fe29ad467f10e60f265bfb5d34b1221cfc814902acd1ed7724b98fc6ea4d59ec59c9fb4345e808205227a5fdb0ecc39e242efb44900a52f0ddf272560b5583a92f008b2ec81c7b4891712143057953ba6db45b1107d7b6dca6b6f4b0d46f33dc8cea2ad892504684154d810d3c50ef51e83e010cd8b2b63587d708e70e89343cecde2b35a02c627e9524c68e3ff84914fb898c4a4994ef9060860d5090d36fe60e9f1f47458722ffa346c73d6f65c7403d1ef9066740b8495360b96c784038533c86a6da100798ee7e559a8ba7ed38a40a74a80c6ff99a36f4b124fb3009d6f7a7176c34307c6a9b4ed6c2b7730e2630daee73a73a9c93527344de029176f1a1cc611c68a14737a93ebe865376126f3b6ce140422f6daaa1091b38a472661617b4ee91aeaf1a3c6541c041a09c28e9bbb94284408b98d8f92f0074525c834a442dbcafd709d5afe13b6b1a45f6aa5ed8f6266a91e5981a87ee4fc104e768b0c8698aa82ec10a65cd7b9be06da47f1443a52ce6b9bb346301f1224e9fb991f1ae2a7a5ce428dd698aee258728f6ffdd186534f709a0507f79ccf6454b58646d3c8091ecbb7342c302328fd6e50183c330d60365b4691e6d5e5659499372f744eeea510cdbc1680cdc9d70cfe741d7f8ff95a10e94048c8e97d334150cff788fbf1d9e8123e1c215f7dbe7ae4ed392edbe15b71f9e0a3e768e955f3b447d8f77a4737805ab53f07d813064e1f77d747ac075c8b7d4cb3f00f78e6edcdd3127a5761aeb6aafd415879d5a593a7b668da85b9acff9ef16ecc1828b11e2a1d3df15dafb7d9919f78af8a07d6f046a90e3f7784f8de8fd10d2f1d537ab99b8c1e643583c045a7edad8da7db9d18611fee42dec86ed5fce0fa1f8cb5932afc7716424fc2ca90692937e924c43dc1534a5fcafb81e7aac5291e1c9780a488be2e50f66f009ba25c491c0cda55868a0c7a967fa6af4da545bbbb2876f7d72024a7f1e8a61145b57c61d4c9c25a34aabec4387bf9e911fce68b5d952f5ada65209ccd6bb2172c37fcf8a834b1d048701d2af44b58ab4941c3192e3ab44b4b6dfd482aff041ff26bc14ab41d350973374a0b5c78c1c4125e94c4db0bb9d4fc93e18349a026d29407aa89b5280b4b30bcd0facb4c43ed60c434e4ddc2b57c2e9b50c1c74155f03cecedc9172645ea00b96500a6bb1d05be713158b51013aa7b99ac5c496c126cd0227d7051e3a1f4b85b95d27aea74c19dda61de47b11187a63e07fd6a377848524d49e6daa3dcb6812886a275185884112b7b89008669a3d53c464d24cd0b5d2aaf84d249f82522ae7ee1e27885e768b78987265fec1305e63a97266f30625360022bae3ef63f768d546d9a36bb0f09f45f07b9596a2ac21a8a1890f2abac2e9216fedafd53b7975acab231d75da3a1f1b6cca482d7417111f897fa42c3d198b364532083cf26f34243db891d0fc9bf44600ab2aed65c0b9a806aa9b60460e8ee711fa23edbb0b00fab806f304b7684ca4690dc2a743c2ed5ea9c49f2ea63d1abb770b2c0633327a3d3887586f8af9c510b702e1f0ceb01413d83e37bf16f2cc4f32e9ac9530ebb531ca506a240f9126d653fe52d8b2ea3e083223e8194d2b9f69eb72d3b52099e80d69cee0c89c56ab5fab969ee50af9bbb5fd6c7e502d03feb3e385d5ded35ca6ddf0c21eca1422ec2a40f9b1847465e868fc3f1fc1a98597105529b8e229918994e24e9ed03951cb90036545d388049e0663895d6c6f1a28d11dda83851dc2a61880f63abc4531a89c2f3037e4e238fa5728784a48ec2b2dd09d1f8edc8a0e680215cda9b015909caf42438cf0670eae241362cf75dfe923745773927067cdb5680cce54f5619ed9ac04af265514667849ee26a9c55a1fb9a2d74f373ff6888b1b7a4b351b83286758a8d1e9c1b8d163422985d1338e3f68cde4d15f3505c5be9e2c968c430557540093e0d335a27eaf1808d3254d64ce9e8202c8d0c0fb9612d4c6c9f35933722efd4aaec7fd87c69fe5ec69b2da6ef2459e52e570cb1cd0fe84ff743314a905d1bac5106d25967616d5dc013dbe5a5a9f15b175a729c79862c466ad9f6fa2836f85705d2de135eaed138b881a0b56e89badbd74002f654163d8ce316265952e59cc88121937b665839e947335a84bc0669e14b9434417bd4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h23ab36cad2cf8f1674e105ce3c75ed1bc796e0d60e45fd9b907f9f3c1c5823a24c33bbfe99e5034efa946534d3043817b7d95c3ef26d03db108f29ed18ceddddde5bb685a2e6a4a3e00ca25c5365132b04d1ae7e8f48be9c27fd593b53138f9e4a0205a38371037c75eb88bda9b385669566610ba6bacc0842f4e5dd59bd5b2c0e7dead7b85984b48f69d44cb1a4c72c1bb45838769377b02c0d010202c193441b5bd2ed1bbda2f545a2ec4eb506728dacf01c4bbc4ee8de8ec1d02939b93b59409e017f5133aca3b83a7371467eb9c0c01ddc08179e6357e851013f7c6a03adea40237abb8d89c809e4fb70e01550cd75c0243a4d2590e7eb2308d1367f9c397eec6d0a89aec1c5ec6b219ab82917f360eca13092e5329b44fdf983764f17fd35b506cbcdc4f5122983eee724a1a19d27def277abd2263ce026e34d636222607e5674cb54ef94e93d022e6cf36543bdcf6ce742fa23553081704274a38a6870193076c3cf0500c25ed1feb6739ef4579a0a6cd0f74d7fe85d4d1ad126fb0cd12320093e1f63dcd3aacb405525b038a34ec89be0410296f531d305dcb82625222c7700049df38cc17dc65f229dd54d4dc54aab19ce8c1e64a016004bc1212237cfc0dc1070765701651398371556d4e5199ab88e2dc3f8ff8d0f4570957476e8389c921c340ee30d3ed38a3a3785754c71cee5cd31bae4532cda88a1400c58bdd708d22a76220f6fee659fd556404a76d2ce5b5c292d7d4003d92b44ad361c87bc9c1669d910094734d56007e48f71890f4df08aba915c375ad8888f35ab621bd925f303ff9e41b31f8e42f43985632cc907433db5c183831d58c35b64bb1a140a2537f2a632e8ccccf61032a8ce2e48a4b99f40dd1c2207d18a2e42ca13bb2766d62f60757bffad6ded92cbc17c783d8a53578fe9a831b79d55e2e132fa31c616a1be0e04e78bed51162b67f985a65fdd0ee610a50c5a05ab8a88155b43e4a1b061f56248ca6d95f6f521e8193d243845647497092339b996c9c16454416ab79cb0c24450095b5f9bca39902dd2376a736df74ffcf107c05d2b31e9584e7ca9fb66379089fe7bb0968e040d0e9e76cd4104c5a9e395bae7452467c13dfd80c9d76a0f50fb93bc3f7c4865921cb8f2b0c5f37a1bd2eec07cf9a0966da0b95760bea03016696d3fc6aec1c7b79d5a881b9991b2c98d4134ec179d96dc593b88ad5e696d8f43b5a0f4e5d1205cef1b39cd84b58c2415c78d4e4fcad2005fc1d4c4efcb31b38afbc11de79477ec09faf39a61bcae128c9539643cf20c6c91769bddd5f3bdcfcf54ba811ef5e4d7e8aafee3fe0718f7e1168f6a6a1ce2aa595d7c34fdaef56317ec23e3079d9c49591b3c20e56517a4e10237af335c151765256211c9d3fa381a4b3160bdd3908e35f03b2b0f13afc835ae2c285ae9dba92eb0eec9be88e406e14400587a481655dbf7d6da4ebc0c9b5ddfbc4374784771424b7f6c85dfa2db4b8c80626c768d5e9e48cc51e8f330a801ee2d1830395a05ac6465af5718b791d2f7dcf9d0c52e1c010ff2b6651af73489b7cb67e88feec25e3ab52137463712ee5e36b6de9e9ba53ca307578ea6fec8183afbdf22b725e5a865b07dc31d47a1ee75c527e138bc4c65c95a14c7335e37d0dbb4a20539a297dd88f4cef2ccc1b216b9d3a0b22ab93f9c4980f2d334f272d18086a67db07d2dd0f790896cb9bfc7ec04312250ac8705f7eeef0253030ff872fb2785af737f5d446b1f183c097e52bade7fb710acace433b991ff9c225a13401c42fbbff7a0b40671255f9791d5592d42dd6d6ce4e362ab6436d8bc4bdf44d3e9e9e713caf51825b1736f4e7ba74a323ba8ffde8e1a3e89741afec6a350be603708b463f5baaf617e3635072950730933b0280072e80d7d4550ae8b66429507f285d93aa6cac546fdb016a93edb351a344f9085ab207ae51aa33bbe503f0f2e823773e4084d8852cfc449ab149fbe14529c55996e835f8ad7b5554880e7a0fd12c8b295388eadd58945aefb258479e4bdfa11f664394c41db0475cf3a30a02bf6383ec71d6ff243c1969bd44678b733846562e3c6f41594837f2a85e3d13f1c4f33ce18c4a993d3000a8fdda606b08b2ec1326227c9acc649de7a3703d66a4764399b5fb7d8d891103e2413058d5faf9b6ff5babbdb7d90065f905a789faa6fb2e0df5e9305d209f6a2dd9c0f789608aaad06f3c4dcf722fb003606ca6d58508dd3480094f8548e6cd8ca6d186d80a2dc3e37c6ac4542ba2b9a72a9238a51096abf1786d81e7e89f7ba2b1289e58a46201ded35a4f60bcc778d66b2132bd8ae575a449222468da6f5442e4f6dfb530aacedab09dfe01f96dbcb2a52ac84a32b8aba5dd4621e0f9858d1e152b89f4cb45e10096a0d8354d401d2459e6849eeb6f99f74c6e48b0297a98534d34a2edc446a91948ccebb25e36825dbb65019ebdeb9c0dcba5d52f5448dcf96aebc27448afc3293b450bdf29235b71d7e74698b48c4df3163d54aa101b0dc39702e40504a0fdddcf4a572a0a94f0cfb552d92e65db0a95551472573e8899ddd7b69c5fa47247286992bd702184c3a154bca8dafebd6e87a7d7a79349738bc8ac7bbaec4a6676cd5537b574e4241b8410ef69c25d39050282a9799faaa47207829c0e3efbde03d87caf6c0528ca9f4984b31bd5b6ec78b83ee34bfc3466f91ee64684563e8b5094009f0fd66ec64bb362c2ee4f8b1137f3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h9acf6dd6a941caef12d56db479637cd29ea64e0563a17061a735f6e8d7594bb8f50d4205bac9d41362e793a471d6808114a05794e1c7762c27ffbc8ebea91d5d7f0d357b6159603adfcf2549f095e05686cb85943a17c9b8f574ec84fbc6f0d335774ef681f8c9aa1d5bab7839c51378ef2cac7df0b9bfa892a8f734552ed9348e8acaaabcc0ef8f06a0766923bf44b74c0ee484ec3b5db4dd13aeb59e1c7be81c00a0bcf21fc363ce86821a56098d0cddc3a16a4a05cf2cc14ff78ad7eb1e5f2af4cd53b8dcab64c8c1d0fa052d4590c1478029402aca7a38c6ea275463b53504d03cc4de78159e0658dbb72f0d593359488d97b1c294d2557f65fb751cdb5720dbfa52e05b2ec9ffecb4b5fcdb533ba617fb5c20e3e480a29c5636e61d416315d74f57312afd49240908ab1c57af2d7001b7897dc60524448372a69570a5cea58c29d65b17c55ad3896e19b0906cb4f0e979cb4647dbe51657ed337cec6f0eb695ea6f77ede2df3dabdc595464e8ba6d604e98a716087ffe0ba9e38eb053988d2d65f7c2a4bc15879603f9125492cd3ecf309a7da913237df57ae6cb974729c39b4aed80a2174e2b27bdd2fd7beb0549bdadd0b9946f94cbdb5661160057df57b78863f7cff6960c5fe521c8dc6e57ba5aaec78c5985922672009b32108b1a3d862af6464976609a16f41a863d747371378539eecb699d6c15ee86a41f0c7d22ca1afbf4354bff2af7c690a0f7121b25c281629cc73375ac618b1c374cf1b5cccb1d6ebae88bdd0500b974e7782521a0b26a1b87fdeefdd0f77baecaea673d7721ba8f7d0fc79d1ac44a08227a6154c91d5d168cb12dbceaec098c9e2902f0c08495dfbca4c5387fff8a143f2853beed8576c4651cc24fc47430816557496ee4ee7c79d7f09ec5ff6cbdab127a7b757cdbcf40cdf61019bbe6c199bb68070cc5024e04618cd6a5494f5e02c2d95eb80772b4e70b7c46779568d050c56d2445a361dfe7d18e7abc4f77e2a34415d7a53fe3c3fe92c5cc9a7a7ee68c5dfa43fa552859b7c4a7af1604689818bc2922eca2914790a310b577d5ed3ae695f1f945395da765eb6d2b9252e628f740c6b43732f484ec3800bdefe12a59da9da5f01e29167d3f00fce0c6ac2dab75edc7ef7bc76d52f4f4b298f7fd81eb0a9c93573650ac9f2bf3783b3f377ab781ac6b4e2f615f9388b55451451fe2bf90cc5a5e2c1d57b51e0ed0b5a0ab2c8a09ca2a097c1f05491044541f0a37cf8ca29ec313a7b9cdc3e4f27b9b33a7fcae739f55f4de6e93845aa4e1ba20cec6ddee3b2cea8bf695e8a564f0700cfe0a8a1461efd518290e0f81e27221835c1f4c1542b6a7af3e698a7e6e7aeda92b30f526e6dc203b4af05a70c16d52a6fa26dc07d3fe526ebd99b2fbe0ac39ab179a929cfd2ea783930ef5e7b32cfd74512135f007c1480b82dd26d6ad0f7707b8dda0f4fc8962794ebbf632f87ecb866285402f23f2365b0bec0c625a13c3cef511a4532e4e1c1229818397d774ea45635df9ebcf18e6bb03a5c9b55a6616abc0b0ed9ad394d9bfecd76c883eeeba408f037c943a61fb6342f2befb4abb6d295d357bf4fa6ea2c6a77c76f80f7175e3de9a07632f5557ad416869790352be7df32285cab90b34aac656f2e766755ada2355aede51b2cf8fa6da7be4137f0f0c3c854cabfcf01741d326c70d449512065ade4d206dc073ef5c53eb9f51a607fb5cb095463b28437c086ef881d563ab373e523b881b89f5d7e7c4cf130f76f7028da62a8f207daffcb4d7be495f63c3af2610f5d5e714df32ef46a70ba4613f9852068e3c261a87a3db21abde90037a606999fe1a2401f8125f4cfc8417d0353959ec3b0f9069ee5c29c7ff529fba37a22aaa870b7e202a098961e8d7c4d0fc0aeb1b547c7bed76535e163b99caffa2bdc67143170bef80e58fc9305ed4f76b3a2df6525803c929b7d76ebb24ec51fc286027942648f11c9bba83e41526fd3d820d42391c44b4abb240f32fce073cb60358810927a893d735567dbae3dfa2c9608b8e01171da598975328548f42eed990e262c05d7f5ee310c0439e5eeb20876b383e031f6a60b07e0025634e05fece0e74f4cd0836e4741859ade71ae4aa19f01230f5c4565352592e4fe716cd03e42a5b0267ced07d47ce49ec2c39b3eca8cb540d98a74b359c064ddd52c992fca155fc4eeb08d1148aac89f8bcb06ba121a11a86d02d225ebde751dcf760c7787d981b2dc8b0f2ea9d54b4404daceafeb0fcf49aafb9cb71294b57eee6ed2ef56a2d3eff63d7093c94048471080022a09216e4353a6111fdbd9c55a3cd09cde337de451ee7a800de57e19654e6a1afc8241a9c6366e058f550658e5309ecbe91952d4816a292eb7847849ab7115ebd2b5e3abcd8f7f48bbeb10900cc20f8dd253236ae1205b1f8d8a976e5f2f7f5ba6b81c6ed720693b0cf830ec96d747491235a9fd25121df4184427a8d6c80ab5e116060b9f997b9943e647045d44ec8e2a55ea022d180b22bd28bac6287c58cf28665888bb94ad65a410a5f36500626ad746eb2af685210a4cfeefa0c654ce9794f725605bc1edad4c27a2a2fd7c38d2ffd345203e3b5572916c664906f676304b8b024ad65b2bca41ee04f0979d9d55115bf344b6d51ea71bbd1f732956af9e15a500268e3bcd0c3440c039d3a754ea81b1355e3040cc8c915eafbbf13ef22b0ad9928c8aa0381d0fa0d9cbb66b94272d936bf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h2a406bda7ff36027ddb07aecd45eec8c37a163554c2b0d77aa64efd886b6383150f53b657936dc3b5253f398b04f348e33666b13f4c7d8aed21e573682d48b5d76edcbee3c93ae866ee5c7e121a0484bf877e4103e7251dc6f670e536c95577c2d3a07d7c3ebf47b83decc91dad4073dd40b85e69b8a4a97830f010cd57f95cf4891439e21c901bfd710a5f9eb123ebf198a7bc248356cabebe81d9720d981da29532a6e943754ef6d46454ea39f13d719a5d3b29408afac6f86b8e341b076e90a295a3b29d21663f20fe33d58fe994119dfabbc8a12a821b487822f34a8171ac5f70523eb7608ae849dcf1967806e8f53fcc6faf8da6e8e7816f8bae431200833e04280deeeb22adceb000cd2ba46f912935e4267f08f5226191f279bdc4ca873b0ffdd97fc866db233112c204e9c178170f0792edd8a5d60e0961a70032ce781f56a0b1efb298d534062265c2850382ed4e8ea0a4dc2bb6eb831e24e272501d799b967aa32e4b3bdc381c8b2dbe6feb4fbab5cc400fcb1636275d7d7b7b0ba75d112e925e07bb8a3c102bbcbc9b4da6b1a9fb3815a667c2d91c399d29ec4854212327f1ee1b6440c4c5c9d0e79776079470183b34a580243b1ae1d7db675de9c6f06eec278aca24ee53f72b589e4f0ed6b9b87e2f554e9e2c5b45836744d1319826c3d85f65698fc207780e20ab27784ebdc4756b03f3b9aafee648bcd87cb64d0bb1c178c06ff550150af8f97a06ab6831f73eb4b2425bb4ef68caa3ebe48a521f08708cf6e483c01dc5a063f80ced8e375fdce041dc7866c37665feeff616a177c551a41af73e023055a6fb81f9bfcf0465ed927d9175f1ef60bf862c76f3c89ea4435aeb1f210705d5f8ab5932792713db484ad40a41ee8381bbb783fc7384b2ceb5dd2b157649cde99157a81be1c33265cdbfd547826ea97aff1def31a239a6c7ef5524ce7df33a3db71e5cd0408d5cee26eaa6adddb1c60fd13debe519725e478a02cffbbf7c2b841aaf73be7dfe6bef86368ce6c5bd09b812d1bd2ae9269e2613ad87d167e2d08c8d1a76e831195e602d008d6c04ffd5fc078a5b649239264f1b415e2f0ceefdf2f9ec7cdd5c7d8301f130596604ba619d78f169a76fe713a44e0d18f422ed8b746d69cd4fec43ef9694ad10e2e3ca37eda274c0bad2e8d452ee0f94d57ec56090c68a10a7de38c9d7ba024b3d0e73f8a322a2c245391ffa94867a96f94a6c688a06f46f462964bb676784dd6846895c56659bbca1cf3ea3ad42802b26ce344a9b6d8a2d54cd6fe6117ea80f3736f8dd1c7cdaa84452da7b215b4e10b7069adbdbd758b45100c7618840e0fce93690793f0a3ee8cd961a95ebdde3d2065ea8c5f769c650b7a7ce7efd345458a755db4b13d5611f552c359965bab605a9c9cf2efb88e028871eaba12bad9d35263211b5efb180496177067ed977c4e116c5723017a671cf3965b4c49fd41aec7770025b2f5e1c7738c5da3639ab6b3e58dcab5a107978e9386cf98a5e252973accb8020b2947a723b1e89fb915e6c01732fbe4533e941593c3c87eccd78551f2eb3f917fe90b1f80df16435865bf56425502e90d9fe33f948822d8c221be25ce10209df9822e277cad159b55e95eb870902b1150f215bf2c2a721320600090eaad1c364a96596494e82a6d9a1885a9c57e0d49d584c753022c78ff3354c5e6b17f9cfe6ce1dc10770ebc6994f87bbbd4f878f054c65da6b4fa7f29baba2b19c99888ca057b91ffa14181af17c508e39c9c199b8f25f7280240041980e60c2c8f755f1154c9b96d1a465dcb8206fd71c5f5dd11d0333dabaa777e8e15fb188ec66a6d43d640fef21de1be23d5a40bd7f648582dfd28f53fa4462139ef693d9e579ca6bbe5dffa8be15fbf5e227008fc39403362842a4a3b6dbc7f893657a8cc11c51684b0571755849adb3e7f8449feb7038dea9bc905fcd052f57520d32e0494a86200481830a4b3d3ae84eaf3e88e7f2b97df965c6000b924c17589648efecf1b838f3da5e19346c54f60d3aa5a4aa61a8e0075f06153a57ccaa787023b1edec6a6145fa0a6aa59b88f20defa42e529a78b15b92ba00afd78a870a8b5b9187c41b3a786bbb79ac79e55da6cf7e4f2d1d2e4d6727e8de04706f88dd5aebc9cbf2c088206de2239f9d69ed69659173ac9aa80e4d158db6dfcc23c8b7828e429eab8058279b76cb6e7d624785781bd7ad9405d41e9b213619ec5d2e2fd0bfa03f322cb16a8e369bb5a3d667f4b56232f94b6d8a8cd1ff18fbe234dd57e23cfe2cb3ae51e766541b7d89b023c01c259f6d160dfc480a2928b4dfdaad8f2567e3e9d9bc311047c23f5b4d83f048f7a6c0cb80252d900dfd6c48c864243030ad416922b198818a5badbbd0ed151bfd311eed49cce26d0ba2e9aeaf9a2c6b4d8d1b31341c8d79a715a2518a880d921647a7403a34cc9008a0e58adcdb6d6035660b9baaca4c909ccc3f4cfda49a6f26750df481d0937a206b3b69c89a8caeb12b2ec818c6ecc79c66f5bbe02755d2a6f678628e1745c5bad2bf3866cc951d57caba1023ca9277b525ff4877e508204ef8d27844fa2def03bd965498206a4e4b9afab1bfdfd7fde9743ba1e5d9cc12491d050f8ff04a6d19bc6c426d78303c68e50ac595a74621694715b1bbe5e343f9c8becfdacf78ce5d477e5b4d55b25fddc86ef46ed4c4dba0e7a31fbc7f8f5605f59d00e045f1b15adc6576bb5eb84d97ae676b220;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h179d028948acf593635bd55b46ae211527599a14891795f959750a088daeaa11a937df80bec1e04912738ebb196cab6cc368e7a79d12af70dc4eed42eb0a8f0aaa7964a0ee67300561a18c82a5473f235bddcb1e75aa32a22092a52cfbe7eb14aece5a0ed405ecdb337ddb8cf9de9cd53256f5e32a280c8ceabc000a5424ffd1cfb1d293dbfc05164f2e6291260855f10c9b326d94201a6efd683df786bc2f55be381dc66421f50fe3e151b3cb1cea5b6b04fc8ff7ae0ddf349f3bd0322da73b49fbebf3027bafceae60e3556e19200980c20baece88c10689d2bca33714233071598c3321b98fd95ca0ae8a6c74b62dc461060f086be025da2c1409115163a6f55dce77f749221fced83424aa7a33f767c842ff324671180686e6da86c54a5ce693ded7136290471de0b596a9f25f18d7d97d4128338940b3f92482fbdd8aa294971a14696fca6a579d2475b69a0e6fd5cbe8400d12484278fe54fb200be931cc54f023f18fff0963efc140ee65d80f75d5efc8ab1c1daaf5df1a846ec10524192a5824243d0212ea507c9abd1e087a3b4571051715dd18f64ad9efd130aef6165e45d9bdb382b47598b90f95450d8c070a2e6f6b97be8c2c56bb77b3acfb38c05ee8ae8f7f93877af721128c929be226f47da2e11ad961500d9c67b7fe9308b9b33dc88554a2905c4b78b21999db4f25746699a43ae7dc21fe9ad038b268556b5d8c0f4b77903c9d28b53a84f9cad68ff5bdc3afcbea2d23a970386edb4b085810457aee1352ed22e840e44a6040661d915c2f776d905b16fe60c3b15a107baec7d7e43a2456b3aff69c59ae96d076050c9d6c25b720b2a70ef793d5f6e49d2d18e2fc107f3574206e3e2946964507de4b904cd45142ff737463bf5f5e3c3981bcfcabc0927f5accf69653b0375e51b9aa0b7c550c850ea1eda91c1b74bfe034c597d0f80844243623f90a6559d021370ec3f0eb4dcb9cc2696195e4545a2b678d24cdeb2ff4118c4288559cd913b4a13bfb900e66cba00d6e8e2b9bec9a4e4b0cc76f425d634dec4462d7d06226b61197c9b452f94c35e095f1f82efaa6a5999d8bb04c78a3f7aa5ccca0b8cfa908cfa329d6beb2b8bdecc582ddb1422366afcb36cb2cb70f4e51b67e928b429ef8025d37fa99e6f2c6ee32c98c6fa4a071ec13d69ae02737ad380b31afeb8b132a0b88172ccedfcc059959ceaa68fbb8eb7959f44784d293df71b9e16f7142e48bf78ea0c95fbf75dbdaffea8e59c08465cc6d811aa391cbc4154ff5317555c52d0ea827f1bd98a6717dabd85b78ceb2bf2894b4c0320f4b9e4fc55a40e7ee531f23ffe3336be2b2b70324f3e2c96adec5c04db19720a8e71333643323eda95c99e3f7d3c5021b95b4dcd05f4cd14f9f1f69beeb9dfeb400151fb040754be4ebb4d2cada7ab768370a9b6726891b5c1f33ef853552475148dede9d32b1cc6ed4f0c4a379282e3cc6099a8e67f09c2fa84efcf4205a78e83e3d05d526450d41c22075cae528df7cd134e89f9a126545782803d1fc6e956516ca651c6427ab93c97a72f7c6d1372a3772b8288ae34920e9d5d46c21c7d0f90979c99315383342a28096b6e907ace414c2ea9f35da4c267aa242fcca1fad6edc65752ac28e088e1d9a608d98e80e3888d8aded2d9c92783ac9811f1af2f09d64c4c6da547587d23dd707fe6c97d8928fd3cf746367fc4ac8503de931d57d39f0230fbddff6a7ea7052ec8d402e3286b1d8ac5cc5fb859fd6618b8fa0f43f4c478d8724677261107efdd6420aa074e23c4e7e9047a55475787a58b25ae8530f1426128c3a1a4f318c381282b303c46f9734e32bc682e8a74955200d4b35f87a76fe30e1f3d039646edcb876f8f4781b3c419cab9f0a609375c8ee840d3ed89fa5fc600a38a22fd723e25ed565a92fef069a7019f114561903f0fc1292c8ba8dfc3b604984bedcf637eadc33508118fcbb10829899ef8a524870077502038b2f4ac9133bd72358aee0d25c94038502733ce1b089dbdd922c35055ce58e89376d5beaf09000e0c6ca7a3eb9e817b28a827892cd305531808a09dfc5e6f364ccb1adff2e22dff0599cd033b443b80eae3de71dcee72c8f42720959a178cb4a79c4b2e72bc90438bd1e1007312e0deea40ebe1ed857776ce66eb38f9d9a572483d910dbb1ad3ad0ac0879a6c9942f87bab2e6daab24c2788f2551dac90ad03a4a4e1204b3d1b415a2a37567ac80ebdbdd47a1041dca45579e04b64f1e4aae9f985a6ffbb197ab58cf931cc5c02e3e831bf7bc58d17caf4c8a31dcd3c10180fcb4a7c20df7faa891b5ff20cbecdd257009c71da686bce25574f2d09539bc11e42ba3ec5ca5ad06bafffa9cf69c53c730fc73a3bad2cb7912ba3a51fb5385728cc021e63344da00b13fd05bbb536352966a00cbc318024599e7e59b83de804cbeeac5fdc95491f67a3904f0286c46f8bddd9617b0d343e59d501cbc0fb104b8e3a85537dd107f9bf38182302b289352d3d26a077e5a730247eafaa4fcea78736a847b86511b7ccfa21dd2b40766302a3a0f82202c9af6831ffa79dd2b234ccb46e6a5ab0be67bce0ab0e823e4bf06e11a7c8e35dfa72f1c12628ed6debb69bd70e915690a088d65dbc19b165d8a3944962a1437cd4b3b9cbafa20afdbc9e1e8fb06291d892d60d9887ef1d11287155326794533d42b1750d56e9eac31e15b18b00542f94539d772d4682d33a10fd6b243db3e185c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h41295ab0d00ddf6f7d73ee01970f5733ac90b8187877c5672aafd973699376d49db5bef600d54b10cda227fc46f0bc1c50274e75c16ef441afdac6591dc5c00e328748c5068b912220bed66250c6d63fcff1b0e5619e0f9d59c633d3d268f2dc977b18d555ac4826b50d33a56c3eec8a502e1b9205c5ac9e68434a681f57c30398db753251418e59d4fc23650a638b7504039649399ff44dbdf42c303f74c14967e76d0d22cb09d6f6bcd7ef3430c1ea0ddc2d897e6075e7ff7cc68819bbbc5290cd79f7ad99c39f74bd44b21fec7bf2716e435cf5f0d65cb3a36cd469e146958333678e8b62ea430b3bb7557fb67c7a8ac5973f767841564a2d76a6bfc9c3069961e0f2f252d5bd3db00c5b39904ca68836847c85aa0fb15a483a01ae99b4e8d3d2ee357032d8400176eaaf62960cec548de2dc3d77189bd215332ba7c36ddbccbe713295e42cfa4c0142621c55ec91e43c8e7d80043b366c0a5cd0ed01056af00fcecf295382b35e9610458b9f5128295d3d10e1f6dfe2e618b5b09af738fa251b5ae94c8255634d65cc7272200c8ddc7125a486b16b5a457fa5e4a611a7c5d47495a614e94e995fa6aeaf5ded45df9e4402494592324b400315b1a249f92087fd5f041609e8de1502657f1459906a01e75a9f8b82ba00102b826ea5a57506b4546ea3e598230e706adebb2c0bb11977b519125b103e3ae2b017d7b18be0f1c366b2265b33a98e2ccf7f7359392f1bd5bf779311c276e1cdca0fe7590e1ecfbc56146888927d9b5ae4903e74c34da1b303d98f9c7b98053c4cff2c2dc157a3648a94ef1f0659f6fe16c4ff509b5d09d680871d60a071821b6cacaba46c26ae03731374a7d45d5894e2365f10bc87ca1e486ebc8fec5d9cf9ed1ad7a661194734c22a9b0f6a504278453e1e7341b231ba35c58af7e7150d405cb4d2692f3ae9f0e37ba6ff6a9844a56ea1462e47e20dcc2ef48392fd7356d232f2ba3f16bcaff36bbb7d069c1408da5d86df72ffca84db38f60c2f75341a7a59520324bcc51a7c959d33d5c9b78817ec8c690f47c5d7bf46ea86ba3d2b756b68e72dd86b96522a82cdb457eb50a59cec2cfc1ecce7bce3a43e425dd54cb67829e7c46c981ddfe6deda12aeedc122126d93ef69f9a01f64205caa27ff6d17157c61761f24f41aa410386f5bb9448660ac134c2e8bcb54574ee629a653156394ce5d12a42ff28443c43092d651f3582e25185c2328c62e42ca46a34db93a868677e938fb2effc067bb8668e26f776b9f484775967c1b5ad18e13fb6058d8e4e9525c5bdc12795ddf449f22f9da575911328ae334ee8a83300eb2f2b7c00bb68bfa733e55d228df5ecdc7cf9c7464d3cabee5200e4d5faaf86c4eee97da396b48fa07a8c1091534445130924426539ae2a347d09bae448273adeed09b08e65a20b05387e436619f59e517b985c4c87ad34514908ab3a498088179f3bfba363c693fdf908d6affca2858795bbd81e56a1f94602705fd77d5da92e42d3fb11407f2244aaecc1b54de866ad6f08365c3369c4ace34edddb02c7edb3a22066bd02d76244157ada4138f4cfe549ad66911413cfdb4d60125116910c959d49570ce1c1525c983d14cd40b7702bb8927c31d6216a7a3468485d01e554e93c2aa0bd443e09b2cf07b095a45a513b54973e1496b2055ae974b1c5b49b29a06381d4fee7e25e9f9d716af5c7a184157c6f621261169ac4f2307ab47f6e8daa7498df7ecdff022bf21c68e558d3046ab3c3b445e1211d456158b09294e82ab11dd6956284dfe03bc7395cae1915a45d04550fec298d39c88afdbcdf627db976321dab9011d6bebd3c480926333d924cc11061271235e73ea52574314a9be9b7fd99ffd288dc94d8fcec609adc6e4739c2a6e7d3612f9456b45e87995d5166d9b1b39ee09c8a81f67d4049fc9ece19f4ca6b88be92778afe2ff2967173f606aee77fe613a328073647b3ae17b0eea45152c6cacb570152f7f3a7fd83e33bd1ea1c629b674fccd3a63ea29ac203ad0bbf84348af06ad0fa0c7981b67322051d3438b24ef3c4574500c8303c30189db50b893f550875f5bd1a7e00081b283bcbe4b327d5a2282de9c3da05a19eaee95b40ffa01b450e39312822d0a988117e701ae3b07f40c789bc233c07046a59a1b08bdc71ced6c6dce95ecd89675476587c11390534f83b41fe55a80585893a516fef939b58a8d7a8d6dfd91a07cf916b5dd041fb59e6f36f18f4462476b0a946c006e152b8857ebc4203861c9ce845654653119d9b3a9b98b43cbf74b9f81bddf5e9062d6137551965af399d96fa32f65e702b1f91b7181d7c8410e4ec7c5f704f3fe1134d0caaedaa5725fc9d9197908e38e5e8e017afa21d80c321990a6b2999e080e0741f947fa7af7914df9ee543c6e78af444f6b7e1e52d977bdc00395720d53d26a9919cfb86d4b736a822c2d7e6455f4ac041279b5822d74d0ee35472bc1d41931b058a9c83a30ba2a0bde8e3383abe4cc21906b0be3ab20432fb1c3e08067fffb6e504178d663309148ce45b8d5e69db43b62cbf92d910157df8bc2885016366058a52e546fc7b5bf12c379b85349dbd997cef6051df0d5255dede0a490cdabde46a44adf4857db18db37891056e1596fb7aece8ad7e465d1520d339df7c0678c5dea7d26916cd8de4c3eb41ad3f5716a19e263f1148b37af1daf8de139542447abe710c47f210deadc564b9b991f2f03a7f498;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h4818df8540785c0c16211a36c2e1ef6592ecc7929314ac4a33c0904f375b1d64ab6a98eb94934f35a43008042f44bd6f10252e9f003498bf55f7590ef136079ecd59ea581fca470970b2422fbe683f4deb6a84a23bcafb382f1084b0a5f9b9dc967f89905f42940604341ccebc88ea71b10d9cf8343d5fd79c523f6464eb1be82420b6338a5be28144e9a598b0d0b59b67955c491db1b346455e23059c6b86875265cf125379488288d138824e4926a1498b0035f4b485e88c1f00aa567c56bcf6f72dc34e99c0e7e5d597d26b2e755f685c72e0641ea224c512098466c6be691b4e5af4ed92661b6780184047888546b8e56514de3ceb4876df8d8a062b752a7b0b6f4b121d89a80fea8fa9b567707394f1794c254fe409deaebb9158314f9945b54b81b8d0a1c3155e4b7cde7d481873660a114e05f4952fb84faba18578cafbd5224178418c17d51573f35da7f3cb732ce09c1202cdd3e9ecf116a34053650bb630207ca511c2d190cece145d1845095e224825a0e39071a5d55065cb601bdac2571609f61fd881d7d30d20e51687ce2e159e6193b9a4187ae3ebcef45f9ec4a847d738c60aa11088d116726734692e770b9c35fae62d0a3f09072893b8988702f6e6c3e0170643416003027866f1e9e3e12cc7a6e951237bd52d59323bfb01d3cfa226922b7bd0914f441dc4e69f7b9a87679bb9bd53a8af9940c81f081d026dbc9d5b735991285bae9c655b01faafbf819e62290f0f8288afc741f550b30da62f5acb96ab82929f0dbd42317c7dd5e38a6f9285e47e0f8274235526fe6ddecefa65b5d5c2ce90991678f65e589888415b02921ed633e80decc331942161edfccceb014c3f969e80bfe1fc6c42a159d750b2cf4a1561e7c29ee53078ac038b310d5a1b102a9c743a00c360a0778469f1119235fd577499d55853435553748b0a56c7fad2d498bf6815dafacb2ba5aa01d8989360eb2f6660b39f62aff6c5b5ad5d58f1dc6f96d4dfbb6bc9befe9ed19b329e6a1cd4b7467dddb39da11664826359d0d9a7bcb7d56141d5cc51e450748e8459cff47ae5bf6a6cce0ce2c20cc22263d59ab7ed6a537facf5e2127cd3264b8fe7d6eb5a373e7cf741e131fd125f7ca16514e14ed5fb9138d99c3c622ff211f85bcb1b6ac7eb64624c9d5940b457aaa0d2edd6ad1200f17ed225326fffca35237074f9271a1a42c40d53b3acba2d91f4ac6bd67ebe84423e3f8765c67910c93f2eab5f1756e783db1352d7a433f8f6f7e9db9b29770876838d3a20d87082e259c93c692c03c6473a5c9d9b66ae76d1757357f794b3ce3389a3ce776f5e405217bec21d96c5e7a81a2c1470ae6ee3912502acf0b4cdf0a26e5ccd47771f4b05f7ca1ab59f90ab1a713f9c1dc805c9663c3b636be2ca29de94b4671550035ed688ac030d817916a5f3f3a6945d2c298b9b8e47592f111b6c9d809d6efc92ac58cffadd10039d9365b500c79adc91c0a1ebd1db192d266adb68792cd3a519410fbd66f141f03dd776bd34dd323f9aa9abb0920d27904e11e9f2f3648881e1551699d6b6aa9309a7fffacc2c3dd549bbce66988b2329b07666ec9b248cbda48e1f080526d6ca24177c8d00c3c44281d7327b11f3a53aa0d02833693d956353f490a0cca7af9a8020f616817a08337450355e11f54d142ff4503611594d1f7ed498699e958aec7aaf0c5f69c5563044026c9c36c894a7f774b1d961d0f5679a1a5e72f53668018ad45076914d3e9b993c6d490af3e066bdbd4fc4216bddcc072c442ee8053cb646e58fc61be797b1ae83a4858fa7a70ca36dba94c164047338e2ed24fe8d0feddeeed718c8efc4bafd72fe03d78d2f88bbaec126c35869279c1df1c59508eb777df990a7cc57b952dca15a73e562bbe793440e5004221ecb9cdd90c805d6c2ea393e772a201bb394ffa65f217dc823ea3676e07c9f5dfdd6ab37ec7fe05b39aba0428910e2818a3fe5998ebb4a2c868abe32d546b6503be666592295c86b809ce5ac304efc4228aabbb0f87c7a6ec5ad7892178e12a80921f65c525990effc43d21244ea2ca8eca98b05f3c48128d0030f7fb7abfb4bd4a29cf922afb907d0a8eeaf73c7d451c24ec06abc321fd5038dda11cd7f21a717bc8670958f7707ac72d5d7e9492c421d32506fc91bd4e5b5745ecf206beec81ca9f16a2142d1e31659130e74384c72d01bafaccab8c7eef7c06ab435f0bf8fd54140a0c2ce44730c8c8bdec10246cadf63c47986701d750ffe989b4db1cbdc0d6a5f3503402d2283016cf2417c0b20e94deb01910a073aa4111917894b6fe01ce7e48abdd5dab25baec6c2ec715ffb5d8d1c9c785f988f43b1368dd9f260b11ab9492537dbb465298380c1ccfbe0e7bf74f0cd672f4784656120eab119415b48c548d5bf46eb89110844bbd75980e9a19e239350d9df8d040ddfedfb82570050d727eae2946dadfe2338e2bdad24f373ca45f0f6e346f5c840d3626d5573edce2d5759d28ce365d951d1b24f058279e2c1f0c4f268ab0d3de0021e55e198f799c35d688ded12b6300f9a62a439061a51c88cbeb96bd18bee2d1b1a45489e929b76cab3af65693b95b8f24e7a164dc40ed6dcfa46f2e3367be2640ee19f1801bcc1a56e3c8c905035b537b945739b874db70467a278f0f4335be2a28f47f3829462e5c17648f3ef85cac9d6feebb589a27ae926e7ef30f097f124e9683bd6bb319787314e32574ddda2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h572ed673c44314ae69a2a507fa9b48b501de17e1aab68a3308fb17fcdbcf048b255d1d92cb334dbe8c432cde538047def1f67dbe2fae99d1c7631c9631cc9715325c65ac9ed1c116a7bf2464111bcd2a6ec23fd8e495a4894757b3a0b7bfc092f58b10b82c55817c8595015f8f8dc1670c31172e462a261d50afb649189a8639d28afd68a9f1927496466d21e27d8ba5fd8352d6b0a34f184bed9794719b93ed7b282ff05279d76d6f48837c1386d2a7bd8073a3e674ad219e6fbf3650bde08fdbfa0e55b0c40e8fd06376629c301c85ecb09b8a437a697f2d0314ee4403dc145e872f383074dd22f9fe672192d60db59882a80917f96de6b2994532c90be522066a5865949dce84c0b86bdd08968dcf85c60683a8eaf64d6354163a896ec13593dfe1c277ecf2e341ad127e4f7653ac561bb40456e499e6b7a2b20afcd031fa80d75f6e9d5ce191e45c6ae0af0f6a138283a4dcd57c155ab302048595f06ae97cbcdea93c0ec058cfa5d4cc6288720e289ac333137bb28f4287517988d52cdbc4e0164e952577a74681b359aac8d460c139a923897c2f476e5f7605cf4be09c9cc0e67e6be220a3eee8ad90111755ce7d82aecbd3a1531f8fadcf54e21094674b2a633cd3dc3beaa46068e1cf97aa5f9736a4da53dbdf1362d16e6b9c9156617ddb199b03752bcf5b278a89e597089e67d3374033967593c4fcae3ac438c10c1854442c154d7dfb5b153d6222e4aad80743b281d03158e0f9fa91a32f4cc78811f2332542df69d4d4b5c07668ca6de33aaac26559faad017e8e86261e25d0dd8c9aa0eb9371130de2b1c1cb88931f373915f8c247cae3fa981e92f8764e9f8a619ebfd83ad3d9c74a637ed6137d03ae2d67e29631975847293420a3ce48db613d104962693e9992ff5797f8c79f1ffed20ca56fa1baeffb46bded0efb63be79b68d2ba2fa9abd2ab054d68e312d90195cc92f2dc5ec0fa26bb40bb38e8668303936919c5b0fb030034e9627e1b77ec07704917345e9376e2100995dd90edd464c9056513c8288d0dda4b9bd71edd06ec3353af3c385b0508e18e63d1f46d6309f1c228eca6273d9eca4062eace19817640f2fd9c31cfc411623eb3621057e7e494fcc1a16dfbb7939c690786ead1e8c1ed24e4081f82cf9919e0c193fb0050ea4eda0bf8e59cee41ed90a99150a6867d5cc8c8d606c5572a424f6485d6a3f448ab389138c61a08d8d6d7e44457c410f7ab76ce1cfca8a0b9828252a3a4d8015df9ee71169694a82a1ec5c4362314e36e9997b881d5ee6a809855010e26147e6bb33b64694ee09a29f30a6131d5f44a2854b20451056fd27076c0f31a3a92727369c8eca64956acebd1f3151b0f36cf1c43efa610c2e8b8dbd3916eaa06b964e58aae41e63ce52b92e373a0e8c2135704e7feadc4644f1fd754834577a38c180b6e59c67abe4af0c4ade9e9b2233429708dfb3b560b0803b4c2dd91af68552e17fd203b1bba642792bcf8cf896c47360db763c9bd048d2e5ffdeab84c326a004736ffe3aceee543fb4ade30779c44f1eb1fb298b528e1913d7dd08675f7e5c36c5eb8ac828022be1e5284bc840e88502c681d2ad88eda132e0184e2cd4221b1158d779b89e1883f4a65308b8f97123aec997062a78a16875ac9e052dc5203b8e046355f6796376162908e512a23db9159fb4c409b0bf85371556ade8bd7dcd54937e62e89002e307bc5745cdac9005610d0931d311440dca3f29e1e440b6dd8b4262288eb5884b6ffb088ece6651e50bbe351dfb2042c4949e7940502e34d38a96129f67815177a7cb772fbb1c9c4c89c2755307decf7dc6c160e2ea41c8bbcf2a81ba8cdef9626fcdd1edbf61ee46208b434fad49d107298efcbbc58b5aea8730b2f6bbf92b2c4f424d0518f3f2e3683aefc7f33a1aa417ae1e6e1409845cf0fe44ecbdb8f010c31873da393a63906d9e6f4126943689bc0605650602393ece0962d3a210dccda5d9d407bd8766468528448f2ae0a43c692af84b46829e90d4688f1a0ec1ce85f24ca79a61de18210a6e213c0ba539ed58903d84424bb10008594ed666e8f27b384d74468e362f1ede90b4e5b805a3fe410d27d47ab87a0a9c0c7af6fc347b4762961dcf20d0ddf0e6bec88ab90ddcea3528d7ea2222d85ed562af3ca38cdd2e2073af69d7f5fc43e3d35a8d20cff6cf32f3f9679d5417092c829f601d1891cae1dfee37909a36c0274f66e3106ee1bfef1d0d1394504393d26496ed51a30bde6893886e40080589e955b4e50d5144a1aeda43f74c15f86c2bcd4ef79569c990e16721dd9670bb46cdbdbce767c466869338189fde7e752a3030872906ace970f627c30fe6d4cc7bf1a2e3b7bfe0d88175827523bc115b5f167ab2ab341c681fae03ab52bfd1fb9c8ee12e34b3ab89f094a05d646a7aefb81a5fadd437cce3124e161bb98416c10c92473c0b20bebfda015f42cdf10071e7313811af40e053db3d5f94eaa7916c783e743a37c716020f88ccaa63082fe2d0a75fafc234d8df29115fa5190338ffc252c170587cb64e44bb0c7d2178e1d6b8675ab6e47484317c3adcc4f653beffe35a8bfba0c4254ca5a1afd9cdd61fc17a62a018b55a944e51741a75ee2e94e2a037e82a5e09093d0159c90bb3c0d4fde41b8d9fe51aee8962aa9d8816b4d0b0e02251b0576edd9a203abb8eb85ee16b66e667ad59be8fcb82bc77aa1c606d26f837b589e3210d34a97;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hd8d1a6bfaba5198e3e57b178ad270626adf353929c17175b0068485706d507341622d4befbd73cf9509c55703fc84ac6ab5f29a0b8ca85f8833ee9b2cfec47b3c98b6e9f12625355866f79f7af873e335677bc5878c9949a9baf4736e51cf30a6ba1f66297d55ed06eade274fb90dfc9c57eb23cb04645244e8615b3c36f0863303275f973ff8117628d3447d1ded48c3bcab72dc359f033af94545a119e2ebb5472eb132b905f5cc00748eef7d4bef26f4f190639d1543e05a2e2975f8d8844bbe62ebafcf11a103193adcdb99b0550164821f100f7f85e02bfa046066bcf8be81b668d9aba20c84780452d41aa54a0306c4f1fd407c482108547a14eeead3e9e1ba7bb74daadb28066447a5a2928428f04d781e080688839f0254ed81ac4670b70daa1487fecf08b8ee1180e1f62fc4f0ef1111dd9d95be430656d475665b533679a24beeda7723171488fb69e790a7eca664b22aa0141b492745e4c819810bad97ec3147c3dd8581c23bc88cccd40c59dc5715f59392de1bf0f94f6fb07de57504cc8a863df3b60540b46b20d681bffda9da52d3aecdb5d300216a79c8df2fa740318643a9b2b01fe792f85e5fb1b2ddff1ebf910e6a241a61060d5b4f1a6b4fff822b2846b578ee389a2b14b986b3ccd7fd1da40ae5fb42d31009a64d4e9f5c17f9c3b735510e64f8216cb8d37db0ddd7a5ee1c3a9009ae353a0b6ffce06c466a839b7014702d749aa5ed9b982b3482d3a428345f927b76fac232cfb0c3c2249eb60ca2145a18c6d7993d5acebd5cbba58151a3b494d8cfa757fbffeb6830a3f7ba0124deff2a7b00cf0d1656cda853ab6867e938cc86444df5cae92177177ba2e874d294f3d534388b9278dfb1351bf899f18152f3e894b345ed747512693a20dfc8c6f50b0cb18097663163982f491882dece9d58b403e3df3060cd2d4df5cadd3ffb597ab11ced8564ed5d2435342cfdd7b89346e029f5449432576238e7e02e12b9fe8ee6ede7a6f19766e968bca2d303b8476a3886d6911cac7cfd5183522fa43a1b2bec72446c04ee3a667526fc5166f8dc2de03ae5480da94fb0f179a10481287d9e93d8a10440e4daf43c1e2a3c0c3f2aadf0e6d2927a36d385245d63a1455ac6fec858fc8aa40c67a747753869f618c8d8dbe45d65cb38c1621de9fece0719714d1c6f66e536fc1b67208fac3fe48aec275e06fd990bcae903fe00ce1990c912b3f69c9ae0f15ba6fef803ef833ed804ac81a6224a4a4416b31af862ad755b42430963d66280d54ba6dd66947ff0beabbb47f5610449928ea8bf4804a2c8d05ac89daa16fd36a6908b244dbf1c4c6768081663d525a2d87f1a2a94b4f419400a953f0e3d169ff7c6b96bbeb8a4ca88f562dc3fbfcd775b9b2e5c48888e2e605de8b85b87eed0696a0d7e7a64adbe23f58911d2bc21e0a93bcc83a604698e173b72bf07c0422c529ffc6ab076b351937d13d04c6c06862bb6fb8e1700f464946ac2413d416354f93d11cd3233d87737e6947269cf35cf08d0a5387d3d987222142f6724bc26d2c4265f1d9d5edef6bcd866c2e1991d9153448f635342aa2622e9fc6cfc694ef98415af892f9fc9bb8493d37b19ee0fd53f08c47de1d0260dcde710244acf0df39cf40f59e6507eba58a13f1a537ae651300aa46848054a5372dc47a98166fb326db858749d7fd78a6241e9b4ce307aafd6226cc4d8855edcdb430f67ea2ff81774bc7fbb01282911419b034731cc3a84e1b53a441930b805f22c16263c406fc86d139cf4311d48cf7f11f26ff0f24c58829c0dae64b00ef6525a8a88e0d4fd8a5a655f809569a526330aed19f1767cb49511d069759ee03065f96730d8b0540fd2a301ddf4947e8cf0cf62304e3425cc0a6c627576c4e30839b97a27d36cb345e5d349207990142dc99a7f9486e1e187cae204ab2298ac6d69b56e525be9aaead66f432e27ea9f5c85355707da14b09cda7fdccc5f3bbc5e28de8e28efb17346ca161eaf96475bf7eb22359fd0ec068ffc85ba0a1214c008265fb4bceee9c76a4b6610193e028eda1083a3b66aa7b5633ca97e63266e4be6d5af6bb245d94fd2843bb6b1440eafe61aee1aa3794750ffd957afcb2fd1082e2b1b499be0cd72f87c742ad623d755217a2d941d4a30af7267fb584284345d9b62ff8f734d75a941e4a79a1a71f6c2e6455749fbd3c578ddcbb22b89c6df7eb1c7b442e8f5d079054b0989088a4451e73177cf6e1805be4ae1ad35f1aaadb6397be12f067c6f5f61a58b5214919b77f3b2e7493b0f3521a416f1c8304219c678aa462d4808bcecfeffcf75fd6f46e945b90a286f2d684fe7c678e81892886e4ebead98dd6d6a582408e568c84cd5b95a7dddf27614e547890ddb924723eb40ff8c1a38fabab322847f3eb095150bd0af63c23a34668742a300bdc036754572fb984ca8978f85648f9338f126eb1d12fd7525712a56606a5aae9b28f5160b8eabfd03812b7242e2f8a0d411fdc03f917351257b73604737af532ff999381a52361571aef92a32b8316ba7419598e1a929ef57950461be743939657bc407341329af300661729d955662828478e5be31f3a47900400e8ce81914d8fa4553a0262770dc326cf71c97230cff30f4cf581b4711332c0a4d1a21bebae163c8679589330b75544765bf867392dd4ab6075053fce56b63646ab056c8371c5e1e97c49ee3a6b6895dc5b5b1b3383536c5f843df08fe5bd0e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf7e04e62f6537ad0f00d8658fa0cf030800f004de86d1824d7570a9da52d95a2a5ed0d7f870ff04e86d6f0a1718fc77f172b0e2b67af5bc0aca77bc4edee4c0cdc2635375dbc090fde9000556c3d42ad2e19b93e4b3d3f9745fcd61f7cb7e5e59d6a97bdafc0d801f5b984c3090758ff97747afd56a3cd7ac1f70fca6d685db10d0b83529a772dee41a6f8850206a69c77be546a95540210f2bbe1481892925f924e7b3692f59a134882a8a5587fc57eb8deae0ef43370e4786e98e3fca76a994bf07216dad93e7d98c7bdc0aa4291365219d157b7c4ab748e5962f92d39011d83017604455dd7aad4ae123c18f8135c3c72b4ed286f4da018f7810029a8edd419e76642b6cfbca36ebf24f5a5e28a6f582083d65f9986b3cf35c1b395034ea59b461d41749b7abb30dfda522db9af3eb3f58b094a94c24fba3863fbd1b1b56adb79a0b30a1670c0f6c01b12ac889c3626a0e2e342b72172da83aa49bd14e9a913cdf2e250bd3f72629440e61998a815eb4766cc7a0564fcc78f24055ac8c89d09828fc5cfa9317ebe60856b4ae7491a00617a12271977d70e3c55bf921236c015a393de14e3b3e10c051c0de2b4982cc69879e4edadbbf8a7c03834ed1f5e9b069c8c57f86dddf299a0cbb192e502f9120cbae9641575a282760c1b55de1d7dafc94a0468d4143ac67f3ff4ab791f1b3ebd67fb87599cdcc6b1aa8974d97936e725da588c045a6a2bce985799a6e015895e3c0e27e0e215427fafc97fb8ffd5c783fe021e3957ac8a467c61ae31adfe8e1848696ac2a4163b473bfd6b0a5654b47ab7411a132912a1f3ff56fa142d095028f806716eccf1e925718a9440d5db43a0f78a2a33a28f015e38f25922180775ef20fd079449ccd5a5c041f3cdbc718a996a797922c16071da830d5c9f5fc693d439a7f31fa8585b778aeef7e6a279a206a5ab810454dbd9e907420280f910a7b0df54a88b005ca08e5c44f1e7fe3c592bf4413b3c4231e1aa8730c682b2694e861dcb86f3c1d0de87db44a1eebc166c0135934f80ac70846ce9c4c39444f670b6455893f80e9d148f0a8032865a7b6a02096b159a9fa39f8e89679de4003943899098323cdc4e773998d4f4bb30dfa6564efbc43c1c8bf15d725ba9b37eb421199258680f2ade98bc7274d60759d13bc254967ae807a5c46beef1b18ccef2ab657762e71270c7206814d81069d2d70ff8f98e4d714d396737001002aeacfd44cad2651e7c7f76058de5dc00437e6428caccf7bc3b51e1fe1705475480ebc310dc45ee5d86f537d59db90b19b3dad6b0152c52dda21340437dbd885b31e79fd09cbd137e03991a0f47744cd2b1d1e0b547ffccd2ac3620559fbc737ef4a93e666f9400951431890460488b3a500ed42e61de9d2a4792bef876be27c1a3044ced90ecc92d0bc33763caf666fc9b0f8bbbc10d3a565741dcab9ca52e3286c0b35f590c4f357d77a858292d6c022b9080b6a3beab03829bb8c1fffab8d923f19b670da3604b49ecbbc53ec68bac560904c53c854f1b02653dbd7fdd5d1287ebf0fd6cf33b3fca1a8e5269f55a3528b454f12d3b10abd1ac2767311dca45a2f1b2493bbf5ed7378180a55f0b14bb17b0e8a6fbde9dee69d1b046a9ab593301d442eefd4365357d43e87f956dd9e7ecc409eb914d8fe30c671b5cbf512b48e2b5cb18e7c8fed0d0616fc99cf53f0900b554303ea14a8a480aabdfd679308839bc2e0600c308d719f41a93787383c9976d79e3c08cb2f4a86894ed3c74f3a1cb937824ed9ac148f3a26c2414b7eac272ecf38f1b549c5e8a41cc67d164b20cd3f4173039b97e6d7661d356441a6fb0c89ac10218b650af8a5831b89c048b2dc24b8fd595f155ad4563fc91029ea591b893f7dea6ddf4f80034d9931e035755c2b460f3176c29849976b7b04a066b1e03ccf38dd7fa5d74568639eaab21df33eb490c5b0d77fed9c1dc0c8beed1783c046fe6b07e26ad6a7e95567b5184df944e4cc6c08ffe7ba91481814974dc144c14f83be0fb8d1f6af8111c86fa46bd391bd414a9e117acefb497a2afaa82a8692b2da1dc634231263cc44c7a71ed5ed889e64abf22e7f1466205f498816691e4e8c52ddf5307acb02c25057bfeaea99fcf03a2c7d197ad3a92eeb26db946ab51067037342089e1e19e46db671eef86a2e01be53e3dad765d3ec16f22db7f46a40b77dfc941f9c63df23d86527f379cc7b39e41d5ba04f9038fbcc68110c9e99ea956510eebbfdd226b6a8ac6325b58445107ed2ffad19cb9c46a24e52bdf37363ef1c17e775a1cbb5cdb781f698396552c0f6f081a3d26962c6fb9676e8289d879d7e195caa4168bd58cd1ad68aea91cb1a46d7924367e998303754aa647825beef755c62d2ef3e54e91b24e1164f232921effa5588e706bfdd7c6bd848b7bc873d419dd06da3354c6b2e2ceca3812e1ffa03f99f22b4b6b3cdc84744a3dbf1e259f4edf3d41373c2f54f04ab6ff3bed8f080f1f8854aeadba887677943c52388c444ec81d9c9d04e0f2d28564accda9424eb1bfd01d3bbee313dcefdf3d4b34acbaf1fe813dc39bfa73a5b3f1f8cc9d52af991f940c7b449edf4cb8ec7b151260569254d16a47d1e747114e4f1053cfb1876622cbe1634592ed26611d9f2348d9a94aa0c88fa324415fe5480e3dc746fa331f09ed2dea6d32adafbddfddc356a738b01cd4cc4c7d3efd3adea43d06acfbdc8c44617d803b6322f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h4a0dad9518e1e0c85c098bb54581a7d8e724332982d8510e0ffbd4d465f24b5f9af6478628a06b296418b809cc48c3d59691ab6eb3c4d1f0fb14892216c697653d29ed897c7276563b583a5b3984c7ecb667fa7692caa58210a81f61f50536092b8a73e2af91bcc35d83d4f296ff88582dd515aa217d48c2716f8cc1bc09e6d98b869ee8d5a1d07d5640a4534e4751cdf66f9500820b6f80364a995606b3eeecfb54c4c56f1b518c3c44179283b0fb6bd3ea9ff45968160ded80a56e48e337cca81dcaeb17e8bed5e102ab5f51d0f12c0f1773eb80f3a6c710ceed216cabdd9ee4a1e67cc07e3048a2578fa59fd89fae369992f2f7fd1c0abe7e3d70abcefc8e48070330817418d5498de08332eaf9fec6e25821b1f617a60ee93d3b09f1106224f575d5204b55a35b7399ebd04337c2d17d0dc96fb08da1de94b591dc408dcc6a23eeb6ec016077510305e0254759596187abda33451ef9886f5a7493dd3121e5dc6b36436ee80f265ee5b9b47916afc0a87e894ecba05013241760b7bb5b5f0642d3aa400b0a62a23c9048cd64e37de1ebbb727ddbae1cececb5541fcba7caa7bd54c1408b8a9f43c08846e7d5fbea6f0bbd215b269dd38950f1c45333fa32f5e2fbe54dee66003e0fa7a35df276963b9469abb651d31007e72e1679c9ca536f35ab1df0e71749439d67c216d368d105ad7b58eb9af37a556db86a36323f98217bfac7d0b4f8c28125165104f84aada45857768a8d1fdb710c3ddbc0e5e99297d691cabdb72549c30bb32d6e91782d42dda871927041c6fe3d8acabd04d9e30cf2c1662146bf5ce6debc732b8f22f858d3a17058c797ef4ffca2df22300ec33704afeb9ebc375fc4de2c418e23843734c7d1a35e86b6d347fbb7983f3afa2f35e4766a7aa78aaf37e871c5889c4a9d174bbe838001f3a16075b4a22449888dc181b6dab09cb3754e6d59a494f53ace928d063dcde016ef2b3272109d1920ffa969d3d56fda02075e7dbae331f050520a56dfa85bf6f92364416162afca252321a9a247f6e7506d697d49f6002bf5fc9735952d94dca87d78adf3c5ca34fa31ceb962ae3457fdfedde98d1d8463c2ac52613656e5a96f997b91263d27f3937797ce6abd88e7786964b2d947ef973c65e49487ddd3bcf9fbe0f48d968b9fecef1d6d0136c18b5f83bdfe360f3b4b32223af710992c0ce0f490217e315b630dbef803a9769f7695575ef6579cd60b19c70b453929ecfed4f9cd81e64792d0954413528537be93b2dd7ffb8857c60e11e481ad660a791b44c05efd7ebe7ac4ad2f40fdc21dd44ee4e65598448e64abd5b71a5e95ddaf86fcb27de452315e213b0d1db3bab81d6b90d5f52112702a81c352649984ad31542dca9dc6d81bdef4ca5846029ce48642884f4fb3f865d8262bef192563b3a3070d678a95e63b587152ea0a378d9f70bdbb25dbff05adc3f057a9e7d01765fd278f5fa4017b84542c3f856e1609714b5b50a877e122daf2bec233fde26ecd94e0e3df9d79ed7d85fc408d633f24e77acfbac6c6a5672bbbe488d5093682aa7a63fc2897c10b284dc332a4a2c256f394f4d677039b0cf6ec40b57169af9357f70becb0dabd181ed83975e767f34029a08ebcc114aadca683628e97dd59781c3638596891009a21ae965ffa975c93222664fcbc0af367c3f0cf7468d5f7d4ca439c28e5819956bcf3b9e76569f3c870fd4d56cf77fa884de8e1af3e792d060765a8042d9e60e1726f0fbc13ef490dcec0fcb7cf106bb3f6d5bfc0456117936f0fa74226e1fcb1360e65ecdf73f5cbb4ce562a43bda49b056b8aa87a215208208962ecbdee07b285d51d6a9c2f9988082d65aef1c3a23376131c40aefbbda5d7bb3ff2ba29784689f9f21a92b1024975b8169d9c288c21b444fb5c6177a1580d2c4f3ae7b5a2df90284d4fcbff731822d11a9caa182d433c93ad755e5544a445d3c6813923f1d259cc2f80b46153717364ada56076c7e720e245b600034c00d9bf01ed7b02bdfc15f703437857943aa04c8ded10495afeb53c60e127518372faaadb85919174c43cb451ebe20e87e40c21093de7f368063e22a7e8d7c47584f0110f0204300db5bcab77da588f729c2d8a8332617a08fe9b8e9912dd61faf51bcc533a9254e17e462e408aa6124f0f7a262c1bf3c6151354cffb5ed1640fd6e9ca26ecb476b6af6787e36c0a412d9d87bc8fb4300cec9c2e3f2dae939531570b39357250e95c37fdea128c1771fe794f898b0450b6d215ca74767b7a8e7ca8780bcce551ddf7f6567474755d51b4e2d2d99fddeb3c87834e95f8607e86737efff9ce82f92aaa6c0d6f0d2d9b471b5502006f42c3a88b706ea37fc27d45668c9b1c9c811631e0073aa997e6b36030e3e9d80c9fa1902ba10d2b3205ec50568a202a16686fc545f710af29d10d73c43e6dd0d87da8fd70682dba3c8c768e0348f76134f1c71853e59fd7eb2349c0db33ff1691b3d5821812539c554cf345c3b45e0fbb7b43e89b77c98c233e95486fd93f9e8e70a9b33a70681d973456900a0163d246f079ffe2337f4efd6b7d8fba1e8f905d9c7e7db16fc7074c0125139536789ae8fe3353d7285c1561de4e6fa10ac43590ec3499ad846c9b01ca611ca100e9a1ac9fb1f4fa52a4144d7ff4f2e868ae7cbecaae67a2cbb6871af6967b22a54953036160fc434e18943f8dc9da28703c2f5408b33e5424046347c2c1a9b8a8998d10e157;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he3b762e1998ded9ae946f1d7efddcf3f0e048d09985b5487ba49086c1c73530dbebbb0398071715d37129b89c02afe6056fb85dc9de5cd5ae22309c60eb5e86d8dbe563b19f6cc7cc2b4be36dc8dc048f6cbbeb2c0978eadd55436e0943694cd299fab116bfad7c52395f3a0e2bc134adfe3ef7008e34b9bb375f35e6e6ba30dd16d945e24fc25e3879a01ce975ed14507e8894df8d21d4719efe1343bf517f474eff8ecafc80642c81fc3e9b0a822e76e7b19ee10b52b5ec1fef901b0ef77039c52fe5f9a0ed0db0bc1f4eb38bb52022813799cd0d0b3d553448ffac2f40bc795a3ce38ed189c929b6c3a5706850bc820bad6c5fce967a72658283f3427261c94b9000b4768a3e82bfbbeebc52e65614743091ae6c653a7823a3cd68e1cd2f6df062fcbb272240ed4b23b9b55a61e97dfc638b4ec76698cb0959f1f6adb5ca198d98cc3cae9e5cd0cead01aebbd24ec41f2df5671b813f8d3528f30a5cce34aeedd106bc35ce2c6153f09b1840c7d0ab112838dafb85e8969950b24d8e1a80d7a8cc1fdf4cd50ffe769e8eba1997ad5567d84bcc08b520d4aea7b6d7f7d469f0aba90038366d0df5057bd555f7186963087f00c9cd364a75f6e8c23efd1e2dd974c6a5c7749200a626324bbeacd71ad6beab425a48c6f1098a9abfe0d36b551ffaa9574bd73b2a34db9635a48c30e310e23767c5ef1a37f1f0d00c72386915fe35c2ef2fcce38209a982473afefda0f8cdf058bac43ae64d4db64072c99b4f7d7e9de6614e7cbf1c4cc4430edb66aff9659b2a554f5acffb10396c7dd70c5770f8017a3dd781a4a426bdc599053eb6942f6b97a638e3b6505fef17541a746ed98276c12fca2f0a9502de0a6b9130433540c4b4be535a9f44178f3c41d5dd3c761fd09d3e4d3ba9de296ac463731ddc4d2dd71e489fdb64936e7e32ed58afd4683e1a840fe7b51d2eeba9da6dcedf90fd70316d3be547c9560e5b72e80dc06c9ee2230c5a3e44210e487f5adad33ad74334f33bf35dd60639489e653a41eb97ccc55af069e1313d87881e338d11e4a22bca7dc387db9e40f1db7e8b01098b86f00e272c17228b5ee23fbc9414b54982c31719cb2818bbec75a0424f9498d5303c235957b3693132e043140e6b6f1e0a6b3993ad18902380f9b32a8bfbf519f6e2467e5ba04c958e4e14238ce988ae1fb1a2a4d2f486c052cf01d2b2af529bade808478edb888ea9473b3ae0a4bc111cf6487e3c084970d5b46ba0780980bbda14b8f01383c1316951322bd8af6a1107b3f429d7235025ef131ad0927d5ae83490ca8c2dfdaf96eeb7526cfc0cda10c1b6e63701f6fecbe54983b58a932a4c3209b537998806ad48d686b16745c5c3bd6350b26721c1cdaa7a25941e206f19d3c8a38903f58df0a782d33983ca1bc0519114002e80eb13e7fed94085d1d67a37068fbf20dce00379c639df036da6eac0a2c4be9ae597c6be1774a3a79ec4cd2224ad8b38788d1cc15c25de60298007ed0b5835068100e7e53ac03025ab260f87fb41ed552b08845e52eac43bb40bd3532694dfaa8f7d8ff3062f416a3480654a065d488b10a5916cae2e94a9e42ef136b9974b475dc741a2b383998bd4cfb6d320249efb6352971862114eed5b0857f23cf8538fb38d5379cf9ca5cd1a61f5231c1b8acbba09ff323a2feeb83c9a99016499a200d36cb53bd77226107963eacd8e6b0964fae8319c6faa9ac8e4e352f438b828c522019d376c72b88ab59f1ede30b9bde5a3b6ce3250eb0ed6d732bfa6e36ab6d4777dd47d4d84d96a0d65bd46692d6dd11567e0557cdde910da71dc2415de89a455c124388a9c44e859d257a06d4339d03d902293377d106ffb1f4153a968d8aeb3c56a880e77730ee0816a564d083f7f57477a1d074b0e3b721718d28d2af085c97bf79017e2523e4398bbb8974617531a539b61c396327bfe2c8c46c2b4d0429e91552118f3e792476e57b452d87622931bb5661d6e398c1f575ca4ba82144edd82ae3ce9d3f8cf53e0499ee42fd3a31619251cd5d03e4e8976b8d1b3e3d2e3d5e613c13d4f2ebf1cd03fdc0314068ca064acd30dd24208867b4d7064fe5c28178bf85adc7d654b1ef11ced460f78f82c8198c5d0483ae105269a72b0da26b513ef3f6d752c68d68d4fa9c53cedf65b48cc2a7dae044362755c197af1ac896c9c2226b1478078bad3b6c23dadae66b470bd0b6c7b69b9dce0e36b67ac7655b12cb1c479f246b9964d8095d7ea5d305177095e8c7fc586b49f8147e0f2c8e5e320b2b6cb0f9140a681ab1619cdaffaa8c25da2baa0357368ddf8f3014af58b3a8227ab6b041d0c6140e1c38e5e293bdf73480b2362ff799d094e83afdce8a20120f48736ba4456cd55316d0fec4bb7cf157cf1420f28d5634dca6184c961c26811287c009c2dcfb8b2678e41bfe90c011bcf0317a575b73807e231d5438df3a97648603adf4691f59333a8fa8c71f0c14f0fecf00abfb3975657949880ba428ba504e5ffd78e5de0e0dfe2c521a4bc7714aaad6592d2403b6c456442cc63bfbc62255df661a69a4dfe6f0e99aa70b11693e3f42b393c34c29217a733db05ca7d0f1361fff480fc0cf96c718c95625d78cc7ed0b0a0619e2447f6c432fdb835a5732d481de04d31cc15ac2e73be159d5fc2c768a569b23621aaebd44aa87cd28809d15311d541d326f4a8d8b6e3c05708c3a80813459efbd623776520832b1a1f9a94b3d00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h4f7d978fcd16167b5c13d98862f288704253de3f9a760fbdb3c1a4b62478c34838fddace62ef227e771a51a4348d7f85a24956dac667b2d98dfe2f13635a9b8d89515f1b6e2e4d7bc70fffb5e69b70eb25c7e2bf999e7fdbcd72dc6466d3ac7c90bec0bfa42aa42721ba4196832ce5fe6c1377632c47394d08ac333f7273009da29fd229cff997a8dc613a55e159e979a6bafd49eb1f4af50c75d5a9eb61eaf2a5c669a1f01ead66c86d0fe4137a93c254543440f3dd5310a39402fe3912eb87c528a713b934ebd1db45552d8642570c69a1ef72414c0b226743a0b9bfd29bd24e4fff0963ac385e6197a74cf2935f9506ba52c3b7fd092f5aaf2144346c3e146abc68886cbbb2ed225af264f379e891849ecb95fad7849383a093f6f347b66fc6fa4c6419e3f67edcb1ec0e0cf11a8a70190e08eceba91e8b1aecfd1084c0b3041f5a1ad02556969257e30db94276fff7211f1a23dbcc869084c19a1a30869a9d149942980a437d1b73e17749ace7bef0fe61cacb9d1e386fdf0912e71b162378f1ca5e65124430a16fb9dc3cf7c82c99831a565623ffb905b37ff63082e43ef12f246bfa44b5f9d3b24b373cc5aaebf22908915dd4f9641d156f4028ab9179bd52bceaae7074525b708858ca99a17147d8d55b138cb99f72e54c1cf9d49cd924f8a2d8bd324935323a696c154c56fd31f7d2a1068efa5c20476866f2aefa6bdbf1140899f8b47c9460b2db7ca349792c9097873b9a822ddd44196a6d723aa9f333ac07176a14bd6822c4eca28b09fb636e1d707abd3b7960bee2e4f02d71a64ee2ccc82325cfb1c4778fee1220587b6b18ea20baae02e433a7f8e40e1d0abacb84ffd504423d6ade30add432a781eb3048e10fe5e243f1bc2ce9d4554752e29f46e3716fc4d85b88a8ee13dfeeaad5fcfe523b3fd1c1cbc5aa0815d19f85e1fb94042e2e6c1f2749d055bdfc76f719683effda2f65263416f993d6a87f232f06fe265ea5b64d01959c542399254e4c5f545ec2d207b73d47334be5c769e46e9c2d80067f022da2545c8f296e21b645300834876e51782d49cd98e095b56eb211f287c6331353ed9ec84e3f57512d14144a447882fc9a230e555f0b9e567b503dcfdf486c23b5f99f55a4741369ace581442750f433e8fc61bc679d9cc5d4292f19cc109fbe23a855d3f399084772335731f4ab18cac5ca90c5baf61f78759f6cdada02983ab24d849790d44b8129a20bcb64f40f6797e6ac980f42959903ba41e10d2597f5929e75d8bec405378003496aad2089b3c59dd3221fafa6d5bb2a4716f875d44f63a606bf776d6057e06cf293dcf31abaf10115450327900f1458aec90df2bc7164a7078030dad473ab59bdbf4786681d893087151958324e764d0140452571b09a04f939677fdee8dc386362d75e73c698b55b4b008a1cda1b65ffdfbceb6168ff5713faeb9c769e9d9b95942a8e636cb90fad41c29f34cf6218f2ee2c89fd20aab27b8b94663b6f8acf6d18579ed72074fb302ebc37b90524917846ea4bbae55d1cdea0e6ecb054af0b8d0d50feaf291cc6fda1b40e9d89dd38b2e3848dd64072eabd3583f4eaee1fbb94b90b998ba6c13480b58107775a5cc76255714efe5051b34e1b9d739edf0cdf3547f9fc25a8e85bd86ad86f108e6236493d4735305bb38bc751c222a49e443ca1fcfc73fe589218ae136722d3547384401f792622eee7763950a895d388658762c0f92c42e15c8a0c9d05b53a0fc52e4cee926d2b5ac91c61fe3523729bbc8cc7daca43598ef9a3383a08591675b0ed03c5326ecb92d95681b81e74799c050699b740ec634996babf964a06f81b3ec37e8b3c4ff000740e35b1a25e64f71b65cdc1b9aed058abd0e4e4433ebc7aae7996a925176fd8879173d7498115529705f42468ba8afe7a7deb5e3e9988b871d4218d5b466b22e332c4a04ec989cca2b250bd755389016c71c333ae44e5ce07f4a2702cc264264b730e688f3d28f596b5473523c965f3405ecf0c0dc2ecd5ef9f8a659e40e10e963d83cb002850750fafeba771dbd1950ee85174130d1f81e29819481ee026c9fed2a13befa7fe1949413dc6a1e10e8bcff09208588c5be03739a2960d2990a11e7cf9fe5b1b26edf3533354ec305e8c0073bc95483ed9fb7f5abf2de7994edd9deb8bdaf8de84399bcfa4ef8706f91da390891cae6b5f9d3c3316065b1a923379934a5609e2d4d38cae72043a811be66f9d6c2b33edb21bfff63e88607b4a958e6d9f7aec2a69bde31de9b79bcfe2c4354227655353a7424ce07e51b1bd0d68d91c5eced4031cf1967566dbd8e343410e5cf3a999c21e2902885fa607a12ff8f95220c0538c322137a88a349260f7212e90dffb8e650beee0ad9a5447a7bfff3323033c4eec301c0149e5a5853283ee724238baa75e77602c03f8b869660dc706569874f2d4f01ae5768bcbf8ab548f58e4a1c8ed325bb3f5e1cb6e04f56742a84d57fbbe9fb30571fed34229489e499cee4ebd26453644297c201f015566efcfa1b6b5e9b1ac4ed634d0784c6c64532ba24f12bc68f2c83e7689b1770a3119879d6a0dd39f83a5ecec1169dcc02fc51a43da59d5c24d966e36b6704c6f80b9f3b400c060c531e3d06a6129c4cb920589e61b400a899adf771e5d2238238ff285ecf01e7a81bb5beef3e9dc4f86d7e4281195eb159ecfa26955fb6b932997ddbfc9143629e2055e6b922b152ef2e4dda389;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h7d2fd55b4ec380550ab2a2dbd39d203e9331c025b23f8bebd6a45536c5d920d0c45316bd1a99407b3f5b5d411dbbaf08976bea70820b6d4408d1318a1f00c9c59d3346b1185d370816ef25e5877867ad871e08deb7cc1a841cafc94496a19a1fff47aae74226b22a0e4cd15b45a44f1c9a72297f30eaef85f21e0e5113ff4e4425cca0644bdd7f74ee33a5907adcb324820467be3d8482ee9ecfdad8a4f7d9a6927ac65b28ea2a7fb1f5a6a88c4e1d75a8571de75210821cc4e7d60bebeea1af660f7d59b723bea64b965a855c4384fd28fa150e9eba0e01e0032b58bbaa291e82401e48886fc9e2b4b08f529203df519965b94a6970565734f857ceb427af21f8450a16293ba7fa57b20bbdc6e49bfa498bc37a12fa3ce217c602dc7aa25faefe90df6bacd3764a3b8907290884a29c6aed4ea2eeb32362e538dac32eb4a62926a23e1d7569f16101b5cfc483dedddc717e231232b31922bc9c4b43562dc938a3d4570e5057c0e967058476eb4b069cad1d611c4adee93e18c38e37406612256a1535a58fd345938652b9a6b537dda9d0d4a31050cca4b7cc014dc4fa0f491803605299783a3ca0170ab85f5f4e4581916b1f02fe7089c9220c7b65abf1596b8917e5da7be77ab9fc6733685b3400b3b82bfa4376ed8f8a07641be94b9b8d7ae95b97213b233079a646270d3c1d9b2d8ca63f372f7f0c37174e54c148e4ffa9afff6973e87c1ab7a89f9e1a0ead62adf9df3a561c3c5ff7d411cf689d0b25718d50e1ecafb75cda7692610338fa7c3ee95447a3e40fe31aa92670b3030dbd2c7c2e309f0811018f511f7a77ee0d675ce015bcce876faa2a279704d0138ff9b085eb4fd3d749b9a2d9d3b37ac2c89155b816d9eba9c0b32e577a870e3934820d59c91de18c1b82881f5a1f25618d82226a220bec07e10a354aa3b8cb4075cd6afcb4ca5a5b54f1a0f605528c01497326fc373a6a6d5b6dc1aae36e225aa31010a71ebcbed6abd241d399b5417446322ef1dda32ec3928c41e9073729e7845ec53ebd8d5f5eb553741f0ab90844a1383109704b5a74bc929bba617827914a436aaf96924ad5dfd2d2fccd19e53f973fecd0d463852bfaa32eead9f01589800a9b3b99c88dd23d6819662a1daec9cbac86319a6b990aec71729f6c09857e495ceff6185668261a8dccf2c3568aaa9df87080ef83e6a1c9fc724764c6a3f533148ea3c992b15712bae8afaee07fe3587b9a525f495e9d1997b0c5ad6d833201e1eed82dcc8fa4f7f0ea39ee5033988af9f8d75df7956ba383032dfc36cf95acf2274062c7944dfba69dfd4a2d8c40c4a313c5e7dec8cc3531d727b84baa28a2bc3e6c00761dd6d14320fe59d583eae91768bf13ace639a9b809551923a6963068f2ab4fd19f9bab187d8ec2a7ba984d34a87c07a7322a771c2dd639edc7a23319180daf4830cca53318e7035d4667aa20cb3f5e48440a56800b09035aaf81497c60a4b5650a4c48faa8400d3cadefe320a18bd8147ea76e93bae7d4cd638424eae112d1d01ee4f975388f350e32c210ae1009359af98457b55f3b0336ad9a5f2914e580c1550e81b533535c3920bb8f4a0a49b84e311a25dbfe374717bb225b5334aa699832945117806271783a7c3fba21b1bd1d040e54199ea320ea64706fe040b60880e8131ae8c9c9a6fc1dcb8716f6202f6b5f1d1fd870b8a891ff97370bea0e3f329a767f3d91c05c6f69a5600ded7a53125fa2a43c518a2b5b9aaec6d47b8181e7fddf69f08a2fc13c601a0726cd92ea8fb0163fae76815442be392c38c576945b33f048a96c58232f6628a20d6a2124cd8e800b3a361787f004e9dcc22435810f3449a5a5f18659509e264b13a508ddbeebe3fd5783cdce274c233f9432f8ae7c9464b9054b42e4f2675b9429df31d9009d5e4b7e650b4aed0e8908361aaa556fd9657b2e5b546eb1e1b486630a6f0966edb401cfc3fdcc8d5a4d92736801e82489e6b28429be4d7ad1219f3272c4ddba042aba00391fdad04267ab467ec6c0a9440dc38d16bafbb5caf41176ac8998e229ad881731f14157a8179cc95a15406db28e8db36fbb95cb51d4f8fb100e675f28a3b99be1f7141badc174c01dc9bf76b759c1f959b65b1363757584ff486d3c4a5f14d4a6e2f10bd832a9cb47bcb2fabab0663c17d1ec8fdab2a0f715a5451671f3dd328c7a09179ddd6807ffbcd1ca7a9c012cbe29251a45965656170a74b332a29fcdba92caf62ed46e7919e3e22c2b1829e1eb26ea1a96076fdcfaf0fefd65bf051ca18df1e00b869469556f697d9a4db6990adff09554c5deaed0c51e8c5b98dd5129348314a12f0bf83ddc41290db8fb3da5c473def8dddbf94022be91054ff58b98747a20600da5f33eff3533dfe61eb0e78021dd69e85c736ada49f14d94dcfe051f59347b366cc105d31d00ae3b6442d798e46614405120f08781ebd8d2b5726fc88ec6796e5cb5e96e17cfd1ed9c61902171b14beb29ae38a1f55ec8ad9392604b8577d068616bda68cfefe57c25e3240023468c30828b3ef14c09d245cffcd75e160aa0e4734fc51edb6a01a2d37e0f939e35aac3a04537b02c99ac1aa474dc6e2adb3d4af80dfd39d70cc40dc4047354223c66c5f2e8ba48a597ca318d883a1aaf143bab7f0ffe98715c9a1c7ea7d755df62b2f49f10dd4c6925f74eb8ea62c838d62cab3d7bdda9573082e0cbb2f5018cc479210f5cfaee667267783bb778;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h736c53471ba336866850c4f01364b6c749b2ba66d62a8329e8ec31c9564b104d207fe22f7fde6f93ab713f0c22dfc809d35d1473522b3ced004dd3db3dcf665e9b1f88e4bf798a05c79921931a4c4cca1a7f8eba288800214342339d96e3b5c50db7536749c7c4db4d92c49d992ed9810da776a0e6968519c37b975ded94502bd3c44428b2a8a153880e59fabb6af8f4d0f278b2cf700c1fef4619f228b6462ae0d1eb35901773de2afa5b0ae2e55755571196645e122963a4754d8ae10d9cfdc96ab390e43a6e809479448519980ddc037188925c12555d39489fa44c4e9d91b314af78a3579017d7fc97d2b8cea2a6e8acd86c38789f7439d80aa97f00b308db0672b26dc9f4f8c8cbf3696c45954c38bd6933253d25571a5bd035aa5b876157fd0998a7fba17ed0f49b6f0d2be031dbd2c255a263bcb0e5656004eaedb9f2c68d98b55c1f0e314cda4b0eb096c0c93423da4832b4882a512dad810613b77899465de67ba02939ef34535983fe4fe99a0186c86965cf0a0b1951a7ff45874c76fdd16181a076b0086172a4c5e3ceacc63af2f843d9e8d096a3acfabe6b1690e96b29d059e5c2e593b5fbc0bb615bbcb5668207ee4cb8a3281c839c23de6dd4fef3973e01458c1d1f4109f3741cc67b7d8e76018377c6edaee9eb07dbe22c6464c23c2777e0c435c217582e557a39790ad224875dffb2703a336b6df0e9a1fc33323495388cd65a829e745c39109e47c2b58fd8a058e79c716c1459f04f5bd939f31c0122511a868fd016348c6bc803236367e165b841f8393b533cac3740bd8594111658c3749a9113d10519681a680a94e2adf0f13c319be4b603e8d556e51783b7821aa114fde32a34235d55c14b12cc1ff7c37ccf0f4076d77eb961d74340733b0a01f2bd077cfbc528d7b56005b9baec8f3884a9e8c0a0a8a14b766e6ffb0edf90cd944bdaae590c6df5b5836f893ba638189e78bc9a0b56d2a9dc71bdee4a167a591940213c73b3b3f7fbd8ba1afb162ba8659ff44d7b035a9d7f87ebceab823f87ee49398f556374cf4dd63beb74af7ba7bf0c87f3e898f0b535eb4582e7b82afb829dab4dfb1d2996600a0431cf18a85f212ad8fb2dde89494ed0a72a4782694538ac90ab05c396e3f5b59343c67e3e85bb76851041517eb38caf5fc531348b4881322a40059e5e1c944672ecc4e992f9f3c9955b4edb5a0c068b673909cb3ed3073a608cd6d6fa5d8d70d60119bf8e6d5c3e7808cc98056915191754fc38129298b7bae90fd20e05b1dc426d91f90351781cfcfc9ce89cc6cabe714a4255f1b3d25d012c7cb22fb8bce6f6709430dbbd0b623c3e256654c56fde913a8cd49e4a66aa28e4807d88e8c6591ebbe6d0b0944be918b7887a50b0ba4d006419f6f9cd7724d205acd19762615ec49f9c44d8585c1e73a3ffc5a7cfb04dab5bc40b3735cace39dac3077e0751f5203dde48ece62f0c85b46c477012434a608c80c387bff86d29e202fdd28ed513c31601e01e30f7172037628c43108877675eccd4891f1d29375dd744cf87f2c30a14f65f1fe81f5226e6eba801a7c503e28bd5c0a74bab190fbfac7d992faf150581a718f303764529abb09b72dda9dd2f21a22f8ff9d300acd356677a9a1ddcdaf7118608a38e4b0ad8d493cde2ba8bf4cb92ac8667c8110da148c4f69e47a75317ea1a5442d73df162db1618997505bc18e733a2fb3d72ccfbb0f0de35d0a9943d7d4918a4f7b6a78c4e737ad8b03ed8aa111397e14b2cac5cfa4c1de82f6a7e85fc26a17634ddd487f5920e00e46c4f2d239b690ab95e5e0b1df0ada2932602a4168ee29c7a94b65976907c2ef24326641598ab11613a41e34985aaa2904ff4d30575b501efd9643388a9f4efba7bcce83b97823f2b9948c7765ca1d7d8ce1c2abcc4942e3356d6816b00a00c30b7c557c29942bc5766ca51b9e1cae38fe28ae12195d59a68a4ccba515be8f153651664d84a7c0ffde8dc25744d62a5cd804b69397beb57f044c933522ee705582404c2ebde137bce0b03a8d8a52edccb3bb716995fe48f53d692ac13477b055b12e4a54b008cdf2c48b1c6488d5abce1e156395df566a8a1c0a77e667edde76cb4c3004bb468957ad7eadf5519d6ad13b762b48dab5661888933e986b37b4e1985bcd4a4645477f5f2f059bbcf910a2b9e75f4400bf504cfbe6614b68dcdf7f9a05fbf802e7590fd89ab1e3305a861b720b387c14fd92a1d8af11ec65bda8b6272d36cc5373a30a5cca8329d3e0c11fac7551bfd70871326c58600fe64a3601edceb1b53524721737b8326e9d2ef75f545a25b3f844dc22295dda034c8894366dd1e7eb48a67464be1aee37324e86e4ff905cf8f1279044df36275a6ea3aba17726ffd1c7f5b37e2652608829b982fc1b4a69acddbf36b2eb44948d009e9e87fb1a0d4b2387b0b2aabe7554007ff981aff3840f86de4a541395dbeb270e189b57ad700dc6bf294ce59ab068e5c8562cf245c526bf0119aeedd0c881892dc3a91fb1546efcea526b87a8c9c855c5da7f3d77fc95f409c7ddcd015c9d286f1f4cc99d41ce2ca66e001e0ffbdcba01b36ccf10be9ed72611ec0bbfc288a23dc5571e379df46df908eb2f759d7d86c63d1647f98d4c555edefbec157c0e11d7af5481218288b22176049ed65526bb94afb372b4527bc9696124c980b2c52171e3936f3658a959197d6961098d38d21c76b5d6414de8eb0daa0ff482e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h85be625351056674b59e8d8d5205ee456b9faef720d567650151a0d8aa13c192d253ec7dbcda9474ccb1f23e4abce3052a5851e83fa2b6b0848a5514eb4253ac96e5f2cbeb27378aefce61485d6ac22e70469127e9d5d447326e655060bb13ac3d307c2c174f81a9936901a818e315d18b26c3b6cca2c2c618f21f878995141d2d14c334809b8fff454c41b2fe4bb3e14f82c80c695e275ab9f7d515efa5a6d514927933b1163f9ebac35913e93ccd99aefbd2f10d2076acb8e8e4552c13a0feacb638efb72513b9193dd461927090aeb2a3ea7ea1ef8a7e22979609cee62d1a6f0af47df4defe8af9b7c948baeb42aa287a01dad7c47853d317adde6f94eb60535a071535c79910ea4bb972ceaf806c181b6c4a779270f315eaa25fb72aeaf32c1797d943c29121cd1a5ff1fb5d3d10a75e4a9f2039ed5b1367d7d4e16d2ab0cab0388a381c86149fd233dd62e62a84d55ce86dd2e19aac7ae16a4f5cd4d90d9de3f2e7bb938058d3df9ff74ef25a57a57e8bd83ed2f5e442898f00126f265712560d469d85844cd8571c8b15429cb88880d63914b547cb4808ead235147c2b4a51ef26151de2d04906c7c36a4bf88ad264336e62ebadd179da9ef58211c935a90ae9b74477b808753d1312f7e14386039f9b5b404c4c42ee1da33eddba2a49fbfc25d784dee78be2d8d23973f747662c456c3775ac8e99b292c74ccf2545a40992c6cab4772b02f3b68cba0676d0fe5023445808becaf9cc7637cfa0d179152a3d11c388493c60048f0363311b7f54be8bfa8e83e45b8e72a5a21c17c83dff372a2b19ab8d0daf1096a974744c0edfbc3b592463260abb19529a3ba91950fd188456dcab96bc2b6b7e6aec0face9edbc799b95f1c9699a489275c3bb7e623d12e5200c8fa13939ba33f1fa758421f466d6ed63e4d820518d4fca34d8a7f8368e54f6e848f7bc86d15b0ad5d2c5d704c9301774b5d2239f13b03fcb3f06d5ccdd182f1e4e84508fc92d341ff435edbb44a6b4c79b25cb30c454c10a711a81eed93243df611b628d80c4c3c47b93a5b2378f32192361bc897f0019a4ccdfba764854c8c13e4404a9acb051eb728e2359ebc54626e95f857ab7fc1c6ad53f4287849aa75ed3ffd20e613e157580475b9cd76f41789a44c6097c9a91ff039cf470992bde6e7bc4f01ae8c1eb9d1f00a1521a19948d576d9969d1402112930a93865d3e3adafe5a3bd6fea368ca580d07b08e819dbb1b0d50e03358ebb0edbadbe5ada0cced86af845469c625319f6a1418580921d42f8db842554ae81fda06de53e57576e9940552c7bedb4738051170e1e3cfd48843de632d5625447367b69fcff56cd519501c31489f8e75a0ab7bfc7588baa90169bbbc7d4f9d30943391155066267083467ac536369d852390da31fea6f0d7b036675b1e8152c25d16c7168952eae0f97be521ecb5eb3fcea4f2ade7c8723e94dab2f76a3e26db2a371ef0fe3c0a1a4d4160b86a195fd76ed853f6137bcf6bdf9b5ca2ddfc5c62c61c6a91a857b8aeac7cbafd9643f3f488172dedfc836dd152a4ee5a3598f9699e8176929e28a11a20ef8081a99d42ae210812c1f41dcbcb3c05f7e9a0260fe93ad2242984c213521cde51cf337b4391910ca8f215002f8ce5e9fefe1b6697acc92be5c6a76cd232e196c06ce7b80af95bd4b9310d0b403edc8452e22e78b2c1c3930a523df7474a7957af2da3cfd71bf71122ad73cf28f120207ff0e8d2829d7a30cb9e2ea036a3e0ac7554c0a712e2b244fc3d9e32cad1c3e0135f03a2ac583182ca3bb6ea25f7057bc8a4bb8fcfca287349d4beb6bffb6b02a1fc52328fa2015a4d2dbc6e806d707935c2775e755e3fe8736ba3709bfe5fba8ba38b2d519e1abfc86ea800ccacf5c40d6b3d7a6d30f7ecf9497875c010bca946244257ff072a9abef59bef9c1e678243faf3ab379fa4acbffafe7f988a6f21ca28cfe995c282c54eb8342b3ef6b07e65b5239b8acd53f73bfb563e9c46a2454dd084189af21ab58430a259e442cfb46f76a16e08661517f2cee481b1fa872c4feb09b659cf54449777f2cc4cce7828f2eb9bf7433417a309bd5468cfcdb51e9a13501795a7bbddfd251392d5cec1dc7e29aaf0f73a96c0bb87e9b027edb5ab9b43908559f01d82084113f35f5c71ef7fb3c6c4388e0272d2aa6e86e4b65d41dbdc1dca15d4916e464d0d6a95c210727d710ff8ea90459ed7c33a883ad91954e1125cbf0519bc9360bd3ac2c958e7792487d395b5aa2e378c9ea803ceb93248b859275ea9f4ad5222752cb5ca8764dae3073cc217ebcafd10436ea233f98cdc50d5fc05d1e4c13f2dc23feaa1365ec21379e2e2a7a5f01139872b53a8c51b33b83575c88932b2565a748cfd136521fbc766f6ac43b380563ed7b50a899cb454279b724895d5cb08bc0e290c8c326e34af2863cec80d9502d6a90d5560a8db991f9a28623fda2d2752402c5e8844b871657d2fba20c7603b06b6933a1e4692eea1a45dfaad3b492eeea8e9068d1c4a05290aea02b5e5f50db06b7d41d5c936792ccc5e7a493d18a936b58c9a888b4586114f4bdbb3664042d9e60fbf979de159019979dfba77bf706ac0ffd96cc3d011cf29def3141469a4562906e534b78b95b433c0110bea8f9dd997d0eb125fdb9d10db2bb874396b5943e2ddcbb728202f4385c36145d07d5867fb6ab7b87759da16e9743d0d33b08a3cca4ed2dd72cf97dc2aa8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6f0206b1b9129f7afd92726df3d31856cb98e7353812b95740ec9a8daa82c1b2c551c2673d47c21003fc3edb193554d8e7501c56e433825dd5bffb367ca4486bd23ccc35d0d2153c1d580a4593443f30ba1c3fdc29854cdbbc1987cc0a21c615c53fb3ef0987c2fb79a12094d8ab84b7469f62675a0c8491c7d7dc0d3b0d44da2d5c698cd7f1b516deacd5e43c76b513c5ec741be560c6de0992312a6fd9405d3d2fc514e22d84d5c717596964d38dbe598e956cbf495bd2162518dc107dca9af362c871bbac29f59de79abd09156f4f02c2ad4399edfede7c11c37ec8c180be383be51412d40af121def8a3d13f034105101842ddaf21f903512173c17a0a49bd9f2bbe515cf9950ab8c9dece40d0c908113b65806413168dd55ab971c47b08d47665efbbd82355018c8090dfc8fe494e47557ee19c93b54627d3776ed6d78ca34698087a04cb60066c8b29beee16b4014a9fcd9401b6b3950b95eda8fc62bae9f10615ae8f020ba3933dfa44ae7e2a8a8bbf79c62c71a5deb9d34daa35a7605171d91f54ccc1d8c2684fa9cd34801e259fd2262161c035ad3798f88760f03a4a1195d5f6166194b5a96205c569585e1b46d892d53bf68004df9ba5e47888bb5c9c8acf7aea1fa70f895833099e81bc49e70172c73d66ed66ea001bc9e601abc8d207843b7c9eb6a9fd87bf6bdddc52fc9faf7650a045ac9c76f489142d65fd0a95a7b37f5fe63eebe8a273e458a04f97803a74dc656fda8dd954e0b5f8af03627edcee33f3f7fde9840eee2c907d057ed1d891e6fd6714bfb7d1d03f02f4b56b825b09d6fb09a20c8af937e724f0c183c7f07f0b705e17e7206c1e4c71f86809bb44ce0b4a74a8631e504f60ec949787c80b066811990a2507b561df9cd8c689181e34d935a56e380a8ecaf17e4a7e1512360e812adfadf2bf49fc4bd7a217b529b522ef31e3efc5f6226783a116e31869a2f051882646726cb7418d527bb74389903fa631047254ba32e56a6e13fd3c3b5e372f21a0f45bd18d096e10815533d3f6efa49958f350abcb531d98a12eb98583eab488623e5c8c6c622f9402b53986075460315823c8b61f280a6fea67b9b99a22c282ea1ef15b85c0921db6d8bb9c1a562fc0ed93f9386acf1a0a5f5f06ea54c3f455696b8c966001d2a9bd217218afce7cda572477ed6f6a04f713ca4005b30705cf88da2cc553db83288d22bb4ec0bd3e8412565bde7a945fb4d2dec78d792e3c522b39d3296392f901fa6134dee1de31fabd4749ffaa8dad883ffc20702a9b305dd03e1182ddcba36c5e9ea5300b2d5d2e9aae03e203e50e28f7108a882d452d01178c8b2208bbe29daeb09a648871bf7a43399ec91424104bc996255787f3612301827476a736d7f72b6aae41bfde7ea9dd5371e3135dfff7f70e6dee9780e1d061fa04d17dea643925256dac29431b0cb301c0b1b8fac05b4533fe4464e6bbe35336969ef67a4c7808e2b563cd6b29194d5be3f92f13e7323ef6b736f984ea84c42763139cdc779b60d72d5a00a3bc626f825a6afecbf30fb663f14443a3960f61b42fac3b83ecfb75b09c6911d78d90e52cee83e8873e89699bf8f079e44e621aa65d864312e08d8a8eac245e048d158a2135da29ccf07667f855a0c2dba77e7dfbb1d033ab46c14f09134263935589eacbbf5f37257dc76fd8d568574c3a62fab43483661b7cac654872eb88f86e58560007fac765cfe905e0213e1ac781e559faa78cd4f50e7467cf7050d93f96496a4711f13c7cd7383b259f1d8150a1f272c22feb0d9a6a65bc606ee2ca06ae2815c6c1f0fd78ed73e98cc330fb0dbd7110e1278d4b226909deb772629998d6d68734375397a736d5ee4506deeb881931858bfd9b60be3be8fcee1385e5af7adabc14ca8762dee8c20694ca5f71de46d4af266c4be22dd4ac5826716834b2abe3621d0a9621a2654766000006bfebf7bd34758cf7667c628b7bfe6baf8f4502bdb1aab20c5ea907de0acf0281a1d007eb1daf88907abe3a6937d17934d1420dc90e4cbf19ca62165f198e7cb56c39365f036b3969a1a07de0b59066ccea56bc76cbb906ee66267cd2d6d9230159b8450206e4b13e2df647d136dd5a14ab60babb8764c670b52ed98130c57d319ca51d922d45654255ea5e04c2826bc0378532e5332f05111dca9cde5aef438d07e2e5347320e1e531c0ceb11fe0986021abdca2a10507af97b6322247347ff39eb2bad7a92e63c616a70c2a2b5c1160d7c769f391cb38054fa592866d83853ce61f005bcaaf8032377a366f9b135976ba6b3a745ce49afef0ece3ca452ff7d0f40c629a67f2280f517d55ccb7d3b396a104d911b2d4c37e1891f475ee0931427babeb710ec1f33ce465e8cf964a7b756ab7660dee7b9e3214b7433e96d4620e8b36150ddff412b82099eaaecd7d48bfb0d196532fd36a43b781807934dfce8e7b093c510a38b93c80100ec9aa30e01879f822c360a027e34c2abf36825c327f3dfcc31ab0741b3ad1f8aac027bf1d3e430042d930f0a73666840f49e8e064b4bc006b130c7480cf1521926d26e05419e8ebdcee2f7106d2d15adee3c6e5cd1152fbd5a8e354136e8a434f2e966fc02ece75868dcf7fe8fde957d731731e15e26b855acd7bf9c4d77692e35eeee63da62ad15fba35a03ecf65ac4e0f1e1ea23fdf73814be4b8034aa7cc838d9eea77404fe2beeea56f47b72388a46e2f60a0839a6394ac124b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf222a165e131cb2777d9e0fe6c85d03fd9111b4e91b82b3c87f219a9b6e2bf2ca19aaa9968dc3ce5b621987e5c2ff1432e2818374a5fa796e906820265068af620330cada7f3e8a679ba6528cf09c8d11b36774f154135b30f0272995adf24021e8961f1f3e1ec179a43a6259a85837c429fdf340447fbad993e8712e526362a5adf53e1c941c1d73840a8d4f176dec8c883d0fd2c07fe7d35cff4d831af9253ee250e3c3f6c771565235d9db190ff7877fe78725e799e14f24537af6281faf470b2252ed447e0afbb60e1bab12a9bfbe6c44920da68bcc0e08141ff70de5866f34ba7626642c9b43c4720759fce9f1f17d0e1fc416face988b772b101f7e0686544394de87b367ee901ff1c3b44a0223064798cebc5988983c76eb45e180689e7280a88e98aaf1fdcfa8adf0d21b6692c29d0dc7f7623b6fb55dc6b49c777350428a254836c263629ad5a0d4ce00aa84cc8c7662c066064b42d80012035e5c0719b86095957429ef7d3a77a26725f48e9a057fa17d499202c41fde9dee2bf0a36da9a8807834305872259124c062a2bbdc7095c5219bc5bf4aba044f93715504104607f2f9b28bbc2b9f581a1d0233ddc245d62ce329ca53ced571502692aaa9cc891636133fdf70d8d17ea00fc639b15a8daa105c3f8e9cec1f7bcc2705388f4f07093d9a4ed8580b0386f44f049369b5a9c73bc1e581c57f96c8fbb7c0745ed046c5048d4393833cae00bc32702bff6336de00d18f13938fb38120595a81628f445831f0acf98171a7244932cba18401756bd9b401498d8253d6441b3732df67d09d0a239d0179cc7a739bfb9a209654d396d2085cfb926fd1c9d5d4dd8f6800795be6d3ed9396c85648bba31cd3db6c9bc8682c5c875a41fbe28ab959b81195d7a3aac597c7fca277c651af0fb1a31b61f622d840ccd320bf9df752847a638ede3d12c55ff3f741945427fd7d2fe5b59112f5b416615e1ba7d132543b3b0c260d1a06c98394b1a46147f3d54d2f29cd0a13eea80472643c6c1f880f0ac6089decb8221e53f4948cade7cf450398319b91626595c191c720f8367a3abe8fcf30ec580c4c02baffcb5281e34cdbd8e6da2a8f40b08ee8911abfee8427d40f5cbf28b332290d48cabe9f838da3f6c57eb8f09cef1b1ea52d5533d6b6b716400ddb8750b2206405214f1906065039db42fdf0adb532da9c67af578057d2e8ce4563979256f8b67bc7545307eff7b296f12cef1855b825feec6f30cce2b3a760a3c552afc1622eb021a97425bc0c928acbf21cfdf78d141e0134d3f045bf4711c1d391d44f7ed4d5da1a976c98a9186f3893d7b77a8ed8f5c07d1c9f70853dfe32b956f141ca2555386010412a3293357dd2682a0255d0d0578988edb754c147ac60ad59ffa530c24627349b55e81c74a90c1137d8b80e7e3f04f79c6a15b826d5ef2a6f38e9da0992259a217246d3f191a9c720d4ec669886a260b4ee50cc99cc2b653723c04c31502d678cbb4c5c1457583a46e720c3ebaafbe6a06be76273a26a0baccb272e576606acc5b1ae9ad312ab8c9bb8209de7a84030d09756761d759b348f2406c8ce2227845132a66a163d5dc1da2fba5a76d91a56b5e81118529dec8cf0db868dae33ec68ad01919e987ee8e2acebfdb030a852b5d4ed7ba72218d01266d4f4c6e25968dc00d5ba9b489eccc55b56a410ebbb74d790040b101d983c2f18e7db6cbb4824f1de4098021b51f0fc7bb996de1f5a8b5fd7539f1a64d26fb1800178e0c02cdcd7b5652b4c84b550de240e17de1f67a8abc2d89826a88eff44d903e362435ab901e68dd8f63b6fa15ff2b0a8c8b4f135a860fc44c0b130b86d14c5358a8b78d1f61f4c6e7009945ab8a7800cfec1a9e4b17332aa14721d0d4f3186616a93f1a9f5769cd8cbb720a4df7cf3144363ada3e1b176d9f6a770a9c4a4db60db20f5fa22fdf99ffaebc492769eb701f4fff0d4a2b6f83db531c57f74fdb98401830cf8f725946d655ae67d3a814025f8e384cb118ff82054329e8ffef2e902803e9cbc546633a785a6c8dbf1563370f8bd051f77891cbe08f072a523a205db9b171f15e620e0cc9a7e59a06a805d455cfa29091f7a5ea06b7d5b7b3a09e14da5009663eadb7c9e05d9076ab364f2b6caa87705606aaa1aaba3e7fb661b5d1b6672556ae8810f05d1ed8716f586d5b13638f78a1d96f472c94488bcdf45f993133b9b6d96d1bae547aea2a329ca2a1218ddbe4a72180133c6813d638eec536ad05b025b3c847c2e6116f03d3003725193be78229e86f688d8ae2352baeefb6af31210994578088bf772fd33f2b24babd9b804107136a29d8c214cd8e598f9c8ffb3d232ae3f496769e558c6d6c3d0c2176e3f73e4bde6891a5de57263888867299c3fc56b0ce8bc4e44ae36bcc0897cde88d799f410966c457e2110610f5dca5e6ec770fe5b30aef86b935057ada839bb270039463ad7c0f5b46bcd72334f92f0d8b19aa0483f97e8c907a9b78b1ec28d76c127ab7d48ab58d67a38a6f3342e19cb2102377f663654e00289f4b9f3e7c78756a4187a03561b85ca370224d32aeb0540b0b3d998a6f71490207e0876414969f2390dc6cd3a6b7e0986a7de17958ad1d93a765a25afc37b8905544c72b4ba1a724a19e475d8133cedd8a1343bfb6176e0df7d07a89ee083c4086e5af844ad2600235bf2e016ba1d2d30ceaaef4eadf099f68e828a92ee35171de24c40a00535b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hacdfaa72e76c8076f84a66793944392afa157675a7e363100bf2090c66254299fc4bdba5e991c5b380f6b82616c62bf22df571d8774a8d007e10534fa724a00f542d115cafe6b532373db92c29441b626604ee98bf0418361442e8bb0ef7d1d21cc1f39cda9bd6e61cb961bd56db5c21e2101c06e7451930098eb34fa3cde3646e11bf418217d823126d09920a29fdd3182bc48f8b616edc7a773bb5b1f8790e02ff1e955fce2ddbe1a2bf5d6e48a10c10f6ac99961ff1eb87b132ec9eaabf7526b159215db8136200ddd0d4c3aca573d34b2b545539ca9635fab5a99bd75f71c18cf61adae3b67737100d0eec3b71eded40d4779e78c808ac01b0dbd922e1c4893d9adf424b2870a46cb8422372140a1704046bc68fc7f22da53b21bb69bd2755e551b2f9b911369f292c61807a2f5cb370a5344335b98f4c97395a6f6e09c639911a023420096ef2d179ee38ac4f745f27e54f3838b9793bc5801761d47ffee15a099f7ceccadbf02de5ec26cdd8c9bea2d90d3e96e506d8a9d445cfb136e48f6d466b99216604441e4cf278f476ce47a77e42e1a897b19e04bd14b7bdd5bd3cc181c4976452c676e4d677c068f702dc1cee0cc196474a2599a9fb6f6cc8bb65430fb947a8c9e2cf9b05aff6fd2a3dd8bc759d7552487ea3923cbb0e844c0fe34b093ca4b12fc56b0de725b22b1854fe7b3cf86ca4b3d05927204dd622b4d3d75b41d5202afc166e71526b24ad8249556f9bdfe7dfe7e5b2c2bb0cb60635d5e4b39b473fc5e1fff86db2f8dfa0b61902cd3f94815dead8285ce85c3e445823397a124fb87915f0cf1e01b8206960e47459a65ca9679dce1ba26ac67d3023d741ad4158794755934d6bc2d1b193e14d88918611776cb367338eb4e569ccc032c2202797353d86a69812ffa14af2e3fa59ada86c8ababee557feb695567670d4e264e1f7dd4bbbeec3f6d51c649825efe2338f1eebf2464887dc1a119d9811b394c06e90168ff7e76be747df26feeb02683712a0a831dd4a813fb6db4c7df98f1d441d0c52773706d8614573c60c86ef7ae8825e009a03752bc334844bd846441fa12cbb674984dfcb881ecd32aa859edd24c19c90033a9a0760c3047fbf30e72cd7a98f562ed363b1f6aeea2bade54a8b727a09036ac3036bcab2a900478843256fdd7233fb1e8c4692366aaca126e4c5b996c035203252bdf6c35e77f69cc10913e157d45e4e8035f4262c0514fa5f98db57b16d38314fe77c54b48855831d2558a0d45323b74b576a0c89735502864a800ee9e5b8ef0d94039c9b202d1aeec3d4a670c8f3c53a0ceb4c8313244b99880cf091a4aaa47c4ec677883b813c933f93cdb3e0b163bffd911830aae3b9f0868cc3d3a81d49b198408abbb7d28a3e50fa33e21a239c3d3a1c5d5ae9f39cef63b72b593609f5671c778c906285812d79218136ddb1dce7577aca3f39baf197a2daf7cc4bed77996ab7b6f8e434f17d0e6733f60bb8ad71dc5c525e746ceae45604d2966478aedc44b18ca1716922320834892284f23af884f5eacc50c96d0548d914ebae4b8cd6057646079697a2073c5272e0366603bc1af79ab288e1e82038e48679148137fac4c77b85589310848d9e8a1429164c5fccd381440e0fb634b9a6a5d669d852ce45cb94c876c53984e9222a86a944668fa069e4c05da79e9918d3cc8c12e345f490f9014fea81af97879037602dc1be5323301ac6a46856a0eba5406909bf6d2b392a1d44c122209c1bbd01d6af72670335e26591e3c716c5bb3facea0f1490943e41a26c41c0e6578146c551b360069c6feca00a3b2c33b7fdbeeef02927256401565a0488b8785084af2583e611b299484b597b4c377341f86689b2b507c58f1d4cdd8cc20feb3cb0e318f7c4d0c497de4f5d6ea574bdb3343d605fdf2ac157ee6229a6a3c581a5be65adbbd89f009b3a486da87fcb077bc59abb90b12b04ac87c25be603cac408bade425b93dd4bd062f1f44810f51411d68077ffaccd437b7ef87fe6bfdae93cee520d93c9addd632bd61f32d3ca962ba2a10f9ac4f0e7bf389e1ad39d2bc9ee845728e666cf4dbc6583045cd14ca28d51417d8268194fffaa1bbe4cda908cc4a2ae32fe633fbebae4167b21369e2d0b4ef8eb09adb8c015e09287e4afd02b7e90a9f4a15617c7c86de8b31c5d263ec91c6b1ac1c18aa7d91dc9ca8ccb374f40aaca142cedb3f3e6880b92f1b2e715a1eb04c8510c91d0f792755cfef300776ed305c2226fba9fa466c102746640b76fdf7d4c62339d09dac3e785b7054e47f6af9d783567b3dfffc216c661aeb7338634da5771e807a765637e10999f34e73778cf2096d1758a4c71f455cffafb357be74817e64af3930a96cea95ee280923567510c53f87ab99bb44a31d7629cb0cbc56e5627aec7a5080d5d8cbe92fe068df0050f64bb63f44fc91c469dad43e38c9de69bcde2942eb06a9cc3ca49c8608d5f1c28681b5b06e241f35035e2337f0c45747ddace4801d7e4bbc4f9cba2e39f29d4eee300dd693cd9e89bef768b3ae8ab57c2672fec8c61720d142984d6a77ac15cd4b4d1ccd7d7a79a383c5840b5cf51c5c0f1c155b1c9ab9a7754959c91b714d778f8649ed49edebac33e373b80e90b111e08022271c0c2a6395cb6e5d6321719f617e78c95d7eda2c0880420d8b1cc60d0095e12930ded23c835264a40f456dff27ee6d1f51332539719aece769beb0406f0e3b89b50;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbdb1a451555a62fdf806fbe0a53a77bea90d62a1e49777f06d79a2f7b97bd89f7be5c5c4431b6f0bf3fb3673d8f0aa3d18bf06e6d5173fca630d30f1cb88720485a4de1eda7f73eadd13f6b9d4c157bc5974f4dafb77bb279cf03ac1e65862d4e0eddc5c23b4425bcf6e039b9c086bfed9057ae13b428fe8e2e6992249b354c28424767f4cabdb3309b7d2daa8f49e7530caac9d08a3896d1ba9c8239c23ac954d19b9bd6a5a05a98bde1d3a7312b48be200f80a11b7c0e15547e395860821631f1ce78861d9e9e54e976c1177e28c2a9340f158636d98403815d2e9b9551895075325ef738d69de10752b0188911cf930fc5d399e52f432b0f418f79dd83d99cc52c7622f8df0ded0df8fb2849beb29ccb72223a131d2ae91f2d445356e0c79791c5d135ae84bc766e42498f2f5d9ec5ee28d6ec619b2f8abcf3b991ec1d99647fbdb990d435720e4ed02123f960d4f2675767191fd9098c714711c1a566deb865b5a55ad38b985dadda87266621a26d39cda5d5b495b48216b4486ba31232898159fd3cc0b5c5d2a3ed062b0d928f904a5ee94850dacf77214a0c16dcdfe2405612bc839566c0fe6360484516564dad141ad78d8926bac6a0d8584404b16970907f9b957b334ed410630140d55c4b362f64b67df027da7a8b8a8f19fca33f4e85942c5d5a39de306c0600d78570cb8a23d0e7041c720c5df55256eb966d2fbc3fe7ae30d8f3ad0bacc6f3c5c73c93327ce7494572b32365cf75cad46888d17686388b85b46d7d4b40298f94ebc55d33ed64855cfcb5130d3598edca10d2d54b168ba7096a013ce55b85e524139685387d86b1f57032a525be2c0f347afffe84c57a3160088fd6e1145f5d439c4a18193d17f1e0a1282b21a3db9b460bcff0a1a126ac1ddefe44d91c6517c1c648708ec8b0e2241953f23a892be7c446b460e3e5a3075daf03ece670d8027dc4e9e51a58decec30405b877cda824a02da800e7250a07debc133ada52678060cd1258cd15015c3b7e98b5797187904018630b86182833d8f295ffd7b48c57dd0cd36763dcd6fdf5290a9603d4afc4e60af1c74bbd5cdf2233dabbe6531fcdee2a889278d7b977ebe85f21e6725b1b59cbc9f2d9847d1e5256bee6a9acbb97c6c2d9b35eb707bac040534fa69d074fca1ed12d296e0cf375a80f486eb68230a19cdbb850853b1353c1bca30c14972ee31bcf742e471c589ab18fdd290e83d98ab6a3d48629151a2fa2c1d727282fed65307372401df5d8ac18adf2d8ba435df9c18b5ffc28f194e3d48df593575b2c70e59f583ce52eb83e917c8f5fe651bbedd6cc982827b569f3e2fd0575155c6df13e64c31bab1d3d70fd83b71c15bfe44db90049850e185f70dd19c569a28fa89ddfc488d6363a8fe5bd8dda115ac3a2e163ca48c7ea86e185fb198738e8e9d3bff529f0b0ac17ee33628cab838583161e9cb7c858404414a8aaf559f3c05596760ff7b65e691b3e8f44e6146ad710770160f2182f8bcef90582c511896ed73b2bba476901e885cf6308c1dae95218701e03d96c66a86077b7c6154d25516400cd61f9d36c1a6c65bd9c06cc587be2c4b45b1a21141ae8ecd01e1729b2eb2833e3b009952a12cc286ce9f6347b89a255ba649284b21d9750e47e6e312287158644b48b0d6874c408088cc1d6be830bcc14c3889ed4e6c18cdbc391ec80fe3e60f73b9bd20f0997681716993989cff679109c515ac1701cdc6d8c38afe3edbe94eefbb26854ddbdb683cdcf30a0d8eda72d1930c74ec2ddb7cb82f7c028c6bf2afb5441eb2351ec5c95053d11a5ec2ecc5c987c7d5dc558e17477b99e7e7d6d78a33f3f1f56f0b034c807793213bd5e7da44a2d6db697a6306c6b6a373df1bf6cc540555890fdfff641630fd0fa28566d59e0f8a6ecc89f97619f972a1ac9c4182fed1897cc5aaa08e51c6e422cbf677fd0b24bc8f16389a7487023c465b25d9376dd9682b054e12a5f87a29c5a939f73300bc3a9a4368c146d018852d8da46918873b7efd12ea44afc4eba4d0a708ccb2d92949a1cbc57314a8020e01fc348b38b1d8856128198adc53c2fb13e1d725a8d044f27ed4d0f229657733b53608e7b99ab9e3d58d56de8a18e705a02d29362315d94d58375c16c74cb561667964b514c75afc6ce99bcf0d7f4fb1bf699626c47d34c517e2ad381aea4811d973894198fdb37a306569eb004a228a389b5a0c76f4626b86635b7b7b92db70a9307c22bf5c7f75de3cda025f243cc3730da294cc09b67eab240b5a353f19fe6726fa7a16d7fd29dc0d1d16abdb4ecc97cb424a427be7380bdd57e1c092f67bad0dd93ac65306f90503c5baa32e428445d375beb965848c606a7d8965926db9a439dc082d17cf8545aca77d21fe3355159a64f6783fa02f7559de068f5a4edf5a445a12cc9b545bbb1d05890b7e5bb7619047198ed43325763926791de8486fbb689797d5b8030de065022ac405a586a305e2679e5600e950fdf5ebba9c42482f560ec57a3ca143c62e209acf2e0169a02667f4133e4033852029d1f169dc2890c7c5cc6eb7b2c652d0b51459d9a46e106d230bd966eaa45aecbf1ffd1df41ff9662d052f636efe5b9e0791cbadf953b02418fe96e86da5c69875112f18ae88c8f1a26b63096240e2e0a2cdad3e58425795d5a9906de1c001fc53c0876281c8cf894eccaacdd833131721df5ae8ab43e3c7b9834d880bfdc453432b7e87ba5ac9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h560b1a80e2282ef154052f6b227a096e966ccfc67805143904ed931b1958d508a8dc126ed1833930f65dae33178edced6f54210b39cbe2cb04e5bbf72f87fb0ae1c84aa7cb25a72c97b5974cfd43215b0fa4e878b47f70c9f9eda935dff61384325062d5104ef1d25bd983d13b0a1182d21c8afb1cbd2d631091befcca8704276a316f0f7b04a09a1267490f4e58384f96bdac31a7af71f651ebe46667573bbb0661be8e52d2fa3c644a5a61147ae11b2799663df2f515943ae576f535b2e4f22bf1dd0d5ed6405a786514f3bb217ac61f06fbf956a3116408567c82ed7c9836b9b61ae571b235c703297f6abd0ec461b2b08ad2db44a7233c50f61e30f88114b2e8f9e0a6e12063c13fa7dc361565c063366243b9db4a08a61ca974a5b9a9bc6ad571129726990b37cc08b0152df64cdfad12cdf85ffc0da62b077426aae14bc32981496791f9cbac31e491da4d5252dd55093a9b8c52fd47c944c2b051734638ad255653a053c09802c0dc9dc8e65d11f43a008667b560a4fd84e19bc04078aff95e2a14fe82f8fdb8878bc85245efe3193ac931c44c34a3db437f3dabf4ff456108a93a7a5219d1b90062fdaf98785a0eb26173a83aafbe719483cb216aa0eb4fa49aba109ac8b1301260ed2d8e56a8c490f9cba3d38b275cff9178731fb24d29b9f754fe62fbc2c2411ac1cfd7793e9a38e16e9b245c98613f3dee2839f51227ab9eaf8836bffee3b55703d8b82afb21ea683380e3bfb1de2ae6f03d49dd1c16b952626f63cf0fcc8e697095df3de3204f2779b88397172519517d17cdb40392dd894838adb2d6ee64d8cb830e95ba123ef1c86b9c5d6cf306bc116b3df5ee7ff518c3a3b8ecd08a7551b67e7cc7ffaee5f203607db2279d59d841a4c34659e0ba6c5bd8a02628149da28fe39dbe3239ded8b2443319d33ecca8a1a3bd8eb1f42938a6851cfaafcf1e80a10a70adb722b664b9c379a24e6941c645307148b8c5afbe3b3916a689f5757c9f4f5756359c2253e6dd490f19d2941a65d6743d40ef02490f62b91e150278543b3ffb789f736e7744758becb51b2ab3219c4caaf1be2c5559f3e4c302f3ae88c32c11e4d018f5fa344a28d983eee0b3b967619756a662c697b40c99344c2001b577da160fe6fd7305d4d0de411ef32cff4ef9e9d02514fa9df25df31c6163788f08ba2f25ab2c72fb1be566a49cb824262b7539c6363b56f6b7ab2ebcdb1dffd4636bc252bfcafd59ab2cdea164cef4ec10bcb8fee6899ef5c3e1b565bd3e03e6aad7f86a220d31798822b49b31190272afad0609008999f52b72efd214d5d9999f88e21e9a0845d4011b73ad1d6b07f4823acaafbc3c1faefcdab4d6ba128458139c1045cd7e799e91f9cebb28ce7004b9ea8335931d29998d02702c16e0e72ed26297a5dbade5f9b3f08d6204638988d946caa2ab118c0d7ce7abf4b0306996fe170d8b3a842c5bfaee9ad2951b5de62a1313716dff049729c66865a6575b3b43f7f2e3b2f2c3b28fe3fe9b267d901bcbe96bde9711d3380b68afa5ddccc53387e3fec005f435779a331b0c5ee77b9dc9421cc8f8191087d1b6a4ab69eb158d3587867d8f4e79256a35fab553dff0503ab5299dc6c0d5f47ad863885b26f44d4e40f360777b175e16eb38c66694434005c37e49bdb02cf4497fecbe6d3a5d7df6005da41fed5613d1ac16c303b5f5673c8d3950a7792811aaa6cac15fcc60ac0661888420efad79a860ef6d0c10cb63d916d354be2c8daa7513166a738d7c81fdf8bcc586702e3a95ae628ec0b7a37f873963d9a3ea54e98ef9b916c1bd72b7a0c4be516e938d5dd3144271f200ab2aac93e4015cdafcdd399502d36d0e632e57901970f55d39b4eafabfd76a96f723a0e064c022915ce207cd5fab2ee493bc88b5b1000c716d9ff57733b3dc7ce2c56b0a82aca39d0dbf8da2e97e888eeab790d8f97d9647b81526c3d19140a8a89247c67a5651dcf49b328d5ac414031ed3d39a8ce5b7ea13b650386d3dd0d0a12722f8771045794efea0b27d72e9791492da3702ce000152fefb86092d16da306b9d1765c17dad8abdb1bc59f209e3223cbda5dbf3efa35de18206d1f0f171fe481e64a12274d2226c746654c228f325c76d4e3351d3d949e2500119b2e97c074f542b70ced4fa23c62e01c184b67749fb0ad6bfa8b8d752450dd4c24c222db66940982da6be0a0d1a8d84b611b9e5a6f654410a8ffc748cf55181f077524edc174eaeb5ede656058280bd809c3fb17e9ad746b5d2e7aac63d9450acc4970ce12e783c18d4dd1982d1edd6c6e48bc01219a351dd782dd283235ba0710aeeb59f8f3bf6648fe9841e3d8897212850055452c0a94d99f295148aedc491cda92d7c463bb8de715390399b9b46ab6dd201b78f9fae01e961bae4078e4382316ca1ef4a0ac96be4c2927d65fc134f87360c9332f6c8f570f52a5b269dda0eb6662f9e16e913dfcb6986396449126ef3ca8cafad6c55fb1bf11a1bd460942fb685b6280406d29de048e7bafbb0c1391e434375331ebfaabc6e41ab400519d5d2d3e89ace6608db9b86fd3e108999ff6dab4ec5facf94ce2b106a504b582824ffdccb8513df0dda9b9f70a92c7f1282782d52d55cc02befbab4cf63623cd95192a4032aec651d9b501c96c1883633186b4d2e6acc29747bf789d7c7fae01603f7a9f82d43a91861805a5edb9d097b3e0d9590376df41abf3bf38a500a30e7d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'ha11b4e3712a296dc84348c23f0346fda105d63f91b944f13ffaed8b11660326df673773c90c3ea1ef33e21d2c441e24a152aaa4a238316c4a72b0f321badcd03fe64790f0a1ff365ad619b6ac3702406edfc1f0fa2a486de1ff0425c2011d7bdd5c14d45b4874aba389698fbb687daaf5bd8dfc6a8585ba95c027beed28242d0c271059895ae610d8bd19cff3479f7f3a9f8bd089be0fed62d25830e35969df9077b7c56391397bf51f7497b5b549193d9741b4842c721459544ebb1bb5af247597e9423eae96b018db0bebecf3fa95cec7ddd4044a34b97e46eb1cb94e0a469951a337c28fc36205e0da7e79d1910c53e40321c3326c88e0bb0de592397960e1a2b75323b4975de0746811465c8d10b3ace5ccf3066e76860103df1c549fc9fd2e59ffbe19b49c6876f808ef75cbc54602f5212dbc4ab309108796ec2269d7715bff96e2acb872fb0dc6bb55149e2a0532a809436f51730f758c7ba2ca0879d55f31bc582c85d979b514aa622fef53b1d9bd0df62bea9540ea9e5441ace84117e060fa92896b1d0b15ded29cd33dfed9fb014d1dbf8e349844e8cd690b96773cbc26e89f3e1cb098811c0b5b502ac9b26df9c936a88fdb5555a9807240aef8111305bc0dbb21efe4c0dd8bc9701119c2e7e81690d726e6776d2d2c6f523a585b96ee13dd7a9710bc26227e7fc0308bbf24c0726f686bba3e394b2d49f77cacf5b49879a7280d4ae0547698fac8b2cc93c2535d559684d4ccb04150c0eb1a6ff9ecb3c37faa4c99a270a013e406a1b4ea05038933cf72e61b601b8e4a82e791d6c0a5e4c285db1fa28d2c1d6f2b4ff99eb5db58c3f71c3ea2ff6584b977b4b985c63fa6211f58567fffffd38515c268f6a172bcf7a85a40e25507cb7474067dd19dc7a2f876a2150f0f09175fa75f289019e7dbb6fe386373b0a9b34a8c27cb1adcfab6bb475719611bb642cb67aacd2e2cf0bd251e50f0b91fa12a8fb8230276551b36ff19f91a4ac5c9f936494482be5835b4d35778d1451e5160022aa28f9935f796180f3c7cab6816a7edfa44ffe78b3657b3d4f6aa3e63876804447cfab362586ab6b19985026afbf3e5549e75fc9a8ef56bb2315e9feccc4c5b81a531cf4cff4f48e57bcd196d4663ea72793b06cdcebfc1051da4142374402253998fbee17ca6fdaad6f3c3e26b9ccf7b29608c056ff16f65dd782957d4def9e4e8cff88a409b24963fc7e444238f36c6a5094af269ac07c745b1d828e6eb5932847bc29bfe1150bd375f0ee9cbc07d09b3448376b28d9270087b813a9e223343d1ab069d36de7620e1ad348ace472e5b30be7af094fa61d8b3352f1fe86eb1ebf824efdd7ebc03052ec042b13f56f9ef3f2f6d76a6aae52031fbf45ebefa70886155605344b5d8886cbe17ee281cdf5f4921f313fd019e76b23a7260860763e7543f0fd5e1f10c4d78e61bd09bf1401574329f7077e8dff960ae1235b5d7eb06bb59c6bcd78bf9cf7539e6dd881c420e1342de89f14d7b4de48a5f6eaa07d86f7009157f3c76e683e072f297c28278a659c0017e991077a17edd43a4e6cb8af937cc49b4b24bf03a194c765f33f655c615e39f4505a6566d800a119d56b7954b53cf6a985e246c1c9db0d598c9ec09c996d16b9b51f4a17a9aa17d8a3d6ebb706e19ad17beffaf8242e02ba35352d0ee1b9abd1190b8dab1959e6aeb258a76040c10da33d45c22b3f10956e690cb7d734070166912dcc4d77bd30f24c07d0d5bb819bd612686883f178a0c8ce3ec692f5bb7d0120f4164bdb9aeae8433e753d95fd5e8bf28e44ba15b019b2b1e4f7fcaf1e5998c516dc065fcab292783bec270ff67c6a4d4d339d8c7337aa3d0ae1a3fa8a4e3aa94d71d6a293372885d2fa721704c5c265cffe93c0aa0cf68859d1b1f97d6aba8e05ec22691dad69733d45261aab7c74a600516098bf14db74ad12dffae3f2ca44fdea8245ff5bf84334c92b79924ada54e7acf4fd8c6e8a5c0b70f344cdc495755bd4e53862fffbf02215a2ce2286ac3a991a10c009e87d9bbabbea3d46aa3bb84e37c740fbeea4f26d0ceaae0c9a46ad96ea8dc10c797256fde6e72537de4bbbd3093d1927275f84e5c632d07f800eb2faf1c8964ccdfd52e08ec34ed1262037d43323a7f01dbd3db502908042f9538729a5f4bb2430936ed92b4c11ac2c31048519dca152f60ea6e17321d20270c318e27c13fa1914634755364a97e412309ac6c7aa3d9369de6c33ab93492aa78636faf3b0551a8ceccf771e9278ab1c2097cc0c47ffd27f0ce6475c768941139782324d7363ac71fa45f47de914b6daaf033c2fd1c561814e9168c70608ff7318845ee2c43984ee083e80a58c46434e22c87cb06cec8f7df06cf7d0d21acee78e7b41c20e872cebaa6ca153b2b62806905c12dedd50900e8e5d3b709921e37b98945ee4739533d68d0e348bb0518d67e372134aad70cea98c2e9e173f0e8802182f5fbf49b2144137ca3d114429068df89569c443caaa1db64f404b3b0cf7951cdc9fd3ae1f60c9ec80141015daf06d4a05c08430e29cd7f8656afdab2cc769c8926bed92b1258e2e880ce5626f4170a4174ae520547accbbf0e16de5757d1e282ff364c1a2ffaa2c405cf6c015c1221061d079f7dabe72da0b8fc07caeab956409d92a70eab2594ab79c672423b44a19b57e6520a8655a3199f29b8e50506e4bd3deb43fb9562d602525af9b25881c7e71b37a7408a62b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h65d46c0a712d8b07ca15ab2a8e77737345ece76210e0fa8efdb10c48b95af825197950f231356e01472edd793d786c0b4a4810349108a9338a1c1ebb625b6e4a9fd773bd732aeb23729c8816915e0ab3364a515351036aa891aa95cbe89b14f0becf3150bdda529f81f00ef9ac87ae4fbceacb9098d39525052085764530c7c6211d1685031b604babe2bd5e5892a4b4deefeaaf009a5387fb0d139b686864b556d0fcddfa9d38729b83124cbad741ddd373ddc8e94127a299c38075d08bea4505204a7420b012f6936b00e608fe6eb7366b675a3c500c74b7ef477bbadac11e23108acaed2c9d3429d53d0ed87f4da266545d3c13e4497eab5f693fc4f5123a5985dfa789685791b7780f90d2b9fe6aeeb327bde687589de996b2954b1cb1b7f09e55fed21cd04f071cdde48e9a9c95450557af7c52f6d8b117afbf885a35b82c8c99f52746868ecc046a3c27e712809dedac07932a95e7bde7a36abe7e45a5a857c97d8c4907e87b1a58be1a92bc0541a0cbfbeb1520d1d6f2dace2241b510dfd0776a299c704e8d253a0584911bec59a7e7c35f7356cff18a6d71b88ec315f15487d13effd7cc7b2b2df46b018d91ed636af78acd68e1fcbef278388007dba3512a035c2986a6ed47ae0e9a00594499fabb13eec43cf80eef79a4d197736560dca202c1c38ed9021795df138fe62f5129c22fd7282e74683f8c4433c33c55cf8fd1e64e8afd3352eb560beeff945d6cd58adf0c61f27b014231d0dbd8d5f393ad389dbfbf0469585a3a030368a8483bca701558944be1733cee08cc480a2acfe00182ac8c545338e43970bad50a20bf007dca1429ae7935461b368ffca1cecb060392c3186e7fbe8cceda31c45f9b08122dcd0663c86611f157a0e4a7cc61cd84244f2d0fefea3be3ca7118f5695bfbafc9939da74303cc5fe22532ad491545f1f78f70a41818992ada21429fb569d43c524a5b134f3fbb217653c9a7e8d7c28d3cdbc52c8a534105e16586e945989a65a7ded249f61c61e46d99eb6195d5b582e20672aeb377fd5212964fb0e35e699a9a2ffbbdfdd73c6611bd88e34fb824e574acc098be23c13821adb876d2229b51b1429d70c9f90b40e5ff72862c88e72261a15d0a60aec6b4a1b74d36ec56e985627b49be352ea9260c6ff10468bf7049edd2174ac02cff53b2daec039463953b6150efb4bdbd80c65094a67e39d9c3f6df03ce1b6e98d3cdd1245fb157e207d0d3af3bb90f240ab0d6a653f02243b94eea5cf154fefb96629e9c8f1a9a3bc98c673f0727a11893cd24b76d3a319dc281def10e98a3309e989dded0a511a2c618d77c561a110c351f4288bc0f4b814fcf75192a0272e72a3ddaf0d518cb33f7239b656825ab52bbcc2d7b25819d848f9d5cd189ed24a20032349c713f2880fd9f624bb725f0e1138a62861b82a9a481e90c4c9ae740b5b97e069c19c909f58e5bed9e31e73b7e029176dbdc180be2162e8713310d0ff0f2dd81f2c299f55b4e0f463ec0bc7fc13ec409de04a4a5226b4af744ad2530307f953022c6ff6c91d00ca0a2d9d1116e3b6b7b993ff5ad56155bc8ce8837fbc335a0f45420f7d26b76628a65610ff1327ffabc05c820807623efb0acb44e4ec01cb18b6f5d396babf0e8d753b6fdbbbd829c0b1f721abd7b191f6858ca7c11e8ed851d8b1dca3b9723aad060a5214a4042d88377bf53bb32b5ccc1bc1f18c92d32d617ada92f3cd98c0c52cf09cf177f9da6ad1e5a597067d29772c152e06f6981b7266cf1e9a36619a60d5887d399153b162dd3a4c500e34e2c87eadc3e3b59483269936d52718a55177a4485c8a21b69a8b927de326d145d3ac0453975f24d0e597410a6bda07856f56c8f38e75f5b311ff47aef4918c70313a2c94cd4344c6989b0ab4d4ae5c4bce8ba7673162ea912987453a5059acebb794ca03ecc3c56ff3932f109a299be170f31c092fe6c4e852eea70923b024d876261e48a3a7611b4b2658302ef97d1e796b0ac9fc6d1d05907d7a00e24391b6beabdd017fc2b5cd8bdd9f5ac98fa9957bdadb0e077cc7d0f54704b43ac6c7beeac3ece26dbe2a42b19d06e5bdc9cfb92b26d421589856709783f52652c04b9aa853dd010b7e5cc2c579c404dafefebbb042d4e389f768692010b3b07060a1241278640bd789c2360cabf9728254cbcadda3253d6c314e9386c4dfddddeda63323b99745e594aa858358f34af641aec94626dcd5d0709fcc1a36889e27cddee508c76e788c2c28377f70079c12f6bc5c8cb3004abc5c0ef1f1e094c8b88cc0a27030a40cf5cfd451550aacdc67a51edbeb36a3e7a64e3b6d62b09015b4ec2e5e2a6a20a4c145e980c2409df22ebb6ff954b947d9467bd4da717a8a26f717967e9e48253accbe1f9ff9846a6dcec3c686262c04311234fe24948d58a571929bbacdfeb2de603e86a4f4aff98db0b40f78d62f9bff9aaaf433cd81e1a27e083d26f4bd7ae3249ed1b4e423fd54cf0f81e8759d020b68085444b364f09925849c9d68c80b83b6acce42a97c109a5feb17aad954e6e1d2a3be0240f27ac596c772b20f0c0723fbff4fa2f6ec319747095e44afd90a4c25f869625688e1a0f145c0c4984ba9bfd2bf51f75edd82abc3140080feb7ce9d2c52aeaf9bd38e9ca50a2effb714efd6869e5f4aefd98773a426b4d6be800654794f2c40182767270ac84e20087cf2fe882cce05ee0bcfedfbe8b4dc37ff5eff62eea7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h26dad5480ba076f8475cce63b900b7fc2aaa8ba3f705346a5b1e52a07995c7a99fa45cfb6a2bb1a5d46b43e15550530a9a39869b0a3d537ebb3c1d262765c6f992fce3218ad9add303126f6db7f6448e955cb9ade665879a37f37fed0b898be29758d31da928614ec5aec4dd2521eef4b80b0f363b312aeb317e662145731bafa7987990b057975d1c2c12dc5bb4a2ebae3457157b54dd48143196d3a0679a96593941954a393f5638208ad335da6ba2c6ceaabd7bb1e3d6d402ed4b0b0d578d4788a490b7bd2258fa80bc0f63064ddf693fa510a5e31ea1763aefbfee78e12786b2d31dcb951db9fcf6f6229b9320fe73cef787f98219fb8bb17641cd62e6414083b1c448371eaae5226b180ec588a3dce6bbd2dd7850ae7a670e8e074b1041de7e482a488818b63761d320d5a167243c79cce221a3b7e48af2d6e418dc0bff57f44130b64405879329a028096fbda767388f4fadf9477c1457fbf86e5100f02c544e334edb651eedeaeb346e9dc658590a6b7dd7ae2db786cf1119ccd42b658072d7b77fa3048ddda1d03f3265e240e7698ed3a56a2cca92bccc2261234cc67759c02fc86710097740b74eb3583849b85a3a43baa4a79cd3599abd15c9b955555829fbcd9ff8ff41ab072080393d3f527880366aa363eba95bd2482cc9b2d41ba288f23f5f2debc40527e999978604434ab6e8de5d608f955106b77c228936bb8aaba0367c960300b17f73ef471a9a25c69b4c2f403718dd6cf435e94be7aaa7d34ea55db90cc4e58a9ddb64737acec9e058646b8ce0b5331520d317a8107490bb8d6deb4ccd1484968badea163f863991a64912d63fccdac3c76ef36b689e8c66f95adc8d84bdee5d39a2e35339b7375ee6ef9ebc3cfed9ac2d8aa842c38419835b85d4e1f12a9bcdb9d0a2b3dac4ffd5de5a43f312184150851ea74885b6f32058108f50ad24035e9b6a7fee8ff78e030290708a45202c82f81a4e939b5c86229470411c8bdda67ce0d57e562370f0940266232bb01f4a894889692cab565b7ca45716b96c547f1ec2ac014635e688ffa8763c17a9785de12224a6a181e3e90384bc89a7f1e1f76be410ae0caf77a9bec075d0b7c824ac5830afb18a4e374cbccb4dd41b66c9afd6c4edb98620e9f2a110de1be966af0688e14b2b9797b22ccec822bc737f0e2f62e753430266bd0ea2246a1676a7dc03491198ddacdbe3fee0fa012dfd942ddb1c0c2384c1dd41bb7b20bb0ec62cc7eb095464b694f124c0fab83c63602a40b447730022d21080b78328772492a54b972ed8cd4288200b6c961248e1b8931a7c461d3bfcdbd6a45b19a0fce63ef99474680be9fbd9e2df0379e96d008522b85e61c03b2daf3794e93b4293121dd346dc6c2bdcf9f27c374af234ad1643fea256c54b904063c2934b308e1a15f93192892dc2a95985487d5aeeb01175a8fbc23fafce2ce734486442941a009b3b7006711e61fa9f53c89c27fecf32faa8ed24a70e3c1091b960ea19b4eb2a9e94d2ca2fde1ab93a3b3093216ed4002e0e98de74e8d5089bc3c558e82bed76db5660d1ea0afda7168a53abc96a176ae07893f335726e2461d2c61f1a5dbd146fe54ea11a1adf6082a3d833c9f0c7d2e3297c6cd41718aac544d06d39b2b6b08a3320b0c1210f1a85b2af6edd95aeb667433d166f113caa9de5d2a458ef9b53ce2420bfb35cf66a24d374e6707240741ac78cd43c470c99ba801b2456168a077c7056346e0785f2e3f79d9aa66f58099c3a13ebfee46166160d941fc7d995741bd191a88d416395a6c6299efcba7639054ae1ed3079669e29f8706ec9a6938fafb0c037fdfb7977ff711a80e0d9004f4b0e9fac7e7b27f42a939ee1283d25459c953dd1e07d193ac4363b27cd47d662b2c2a34a53a6988df84e7a737e3f031e6df5f050ef68882057bef7bc5fa22effd74317b73da90e9d314215a0b9a41319c287c4955cbcbe62fd2bcd6396a1f665482f894882fbcd84ce38c9f53f6b5ad14139ff74870ba43a13ae85c9f98c3abbd5d77a89b5f3bb66513d0c0e433cc9976566f69f439c1e4d59384c61f0b661edc978e021f10da825ca2a944dc37a96ef395e0e1fda58b1664966cd37105d787593f0081ac0b4e9e3f05ab8a4105cf7ec3088a3ecfda43a333ba9cea853c1b75cef3b77f96b470d3ea7be2a2b5fedc4e48b8af281e00f11b76e3c593bc147a6ce7c582cad606b124fba3a582d0e91560d7e7433530391d49ecbe04a387376b2945c8ee1929188bc61d4ab2ef1a351fc566104552ac61a6de710444631c5163d0f4dc6d1569b525df2a19584c8b928418430b95b3481c887d57c5ff44b2465091221144c98ba68508c1409e11d18159ff973a4b302e3fdb73de33e5587d9d37dfee4140823b13f75ab66c32160148a9c8ee15030748ab4c2703ee41f3456a66f00903cefd9f5a6e0ee345bed07a8c35ee9a752c1691a3172ec6cb44b712329e2c7ec985671c441c34e8af6a5a66b1e8b2922272645daab172dba38758fb9f3de8ebe7c533302efbb40df6d9e44e2e3f7f5d3f8b5061ea2d7fd317b29dbdc14f41437725f804c6ccd6d20e1542af47d822a0028b366920520183bfac3b32a3607c04f215c64ac5537a4355b6f53a406c967809298c756b468558007e980d18003d56e10a0f0b2787d96dd663bc8f64f747415e446afda7ca384eebcb9812586ed08953c8131049b8464df5de18fd84a36508abc7927;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h10b9fe55ff04c2c167368387801c4553a689bab578951d1bec3f21566a5bd631af02ced46554e42ed4bc62c2f2ace9d151e2fff7467fe70b4410ebd332e28b0aa245ab50009d9dc103e4909abb95b5c80ab88516e5ea592f22d178065a166247214d744a6c191a8b0af021202f1875d89a82a461853aec976e864cdf51ea75b97852f470f483ad7baf5eadf70821b74e98c8b22f0b3c88a37d6354f62977da8759a33075cb9caa795da7d616176c62625ee5825f776262429c31bbfb7f7ab0a3779da1dc453958caa5b45f7084f9039f8d34cabdb31f2bcf1db094a676bab1d1006169e07889059ae4c7e1655219292b2e0dfb16e966d52596781136b19d42c84b88c4c8dcbabaa92ba88e3e161a523bfef009077bb307435959ad940f9ad118c5255246c20965fc0e6c21d8e9bbcfb2d6a3d87a97f20bd47ac1ad8d6c14acec48719bcaded9fdd3cca0be8b16e5412435a97e8fd0a605b4278662f4f54cf5165f1618f29d73ab0ee94f77f2577355fafa3cf95504c5553358c232865b9420e70194020391713fd8fd76ef908338b192a7ecb7db790a74cb140c6ed56f329adee98d03ab85e2a272866bccae06bacb5c43124f264a8a3c64ad4e5e8f3970562ccb2c0a43b4ff35d8922c0aefc51da724c69fbd27d4099fc81e433995ffb82c6554f35fe82d6d05885aa99ce58adaa1e0ddc442f930e40453a526712635828e6561b8752a0ef3327f29935a5ebb0eeccae751d8dd377f8d62b2f70c841b5c6dfa2b06430716f803fa972cf3b310aa66038e65f92807a484cc5ff4aad31c703084c7a33873c07f470e651261b6808459cda2ae5d16160077ec4b4e66c4058dbe0c8568477df7d1e5919162e6f47be255349f98ba244a486f3051eeee57aaeee09a7b2a058baa62a45f502f14063091a400545f05e663500c885824dad9a23cc1dc04fa2b40ad541de4e3bd4ee1f5d38d8535391a2dd1aa521a9eae565473a0e84c16fef57bf0bea054fd6ac1671157dc1abc6b2a87f255331032fe854f9ac2fa3b6d639303694c4f5c6b64b4f8399afc68d95b21207e4e00d36cc55df4fd279a2a962ff0cd00588917030057276e77ab813823c564b43a1a811e3067fdfb0819860c29f52b64d795bf6e1012a117a207c0e34c153d3cf1501f0efdcced266d7b78e4b5f391690ff33560fcc3305ddef10d7d55cf933cf7d3bf753da218a4de217bb7609ac137b82ba5a15a6c79b6ad9557185298c44cba5313a0f41a4869fffc742ef26ca5b6cdfb06910e2b92a1dc15e4e7aa21bf0a7fc6c944c1b10d4c6eb002e1bb86b2c5656dc268656cb840ad515e5b3414dc4b653070dce855488719371f861d63a6dcb44095fd51d68dd40b3e6b2a11fe6463df24ceb0e44f653aa1b08c04aa18978eb2d3e78f2793883ea851487a8a2cef8ff372786bf985d461aef6f42a727f374bd98ae4d36d1a2af871075d04a23f424f7e956119e02f71b5456dc478342d29d4de4b8452a83c0c13b9d1469c4c96c0e1e3cd222cec6bb0e4f5833a4bef71026f3702ef1f46402b9633e0f3ac03aaf961d1781cd12894b9ac6ee2c6d33608f2b8d2a719a59061fea677a21b64455e2459278731249d9eb919b3523d9e9f169fe07a4d2a434aaf5ec93b459c9b4e537397fd92a75f636721bc78475732429055df05e43772a6753c36ee6b7ce67b15208107748721202ea39f9d7c1d8d716c147cb2a17d8dc0c2ddfc824d2336495cdef71594142d3c58e3cf182b18a30a53649f69d21c168b76aeec89709425ffb8614d7d00ff959564599710251590771fe89539ebb2e5f81f68184c7983f815f872ef0a37d3fa0ceadfc304797ce06ec3161ccbae14ee63a997176f840adf8c21e5239c938b7f1d83c3cfaf106e2a949fc38b1b48b98c496a8730c103f0d4289cf447d36d89cc6399b73e58f8fdd9cc3fcfa5020afd7cfa73f2f55c0c56642699c7aeaf10c71578f69c5032b8df4a4e54d48e81dd18de991307d249feb9ac71c7d185f82f6d0f6497dbdbe0d09236c35b33e74695864cdec2548ac8e4d051d5fb96ee26856822c3f34d07c56dfed3014eaea0c74a843c2ae69f630d9a8914487eb564a0d92f4610ead447caf94eb7717455ad884a06f295ae0e98d15344fcb3b9d3fe1df7754beab1e1d3dec05b8edcd20b6ea7ffe5134a5c3bd73963efd93a1b6a80eeea01b0e9fef941829e25670f4984549db9e97b24e8ba3459115cc41b2e8c19269183ac3d3575ace0131a8d882986275b8bd075a242bf3e252304280a954b5f67d34bd2db947ed1d7c329f80f7a6156f0f8275f70e28022f9c1ae8eabde73d6e5db912678c29870cef77f755ff67315b0c0edcf05844548c2b2430c24b57f2effd8edcb10acf331e0d578204f8fe69317bd66a44ed68b036e68a36ff77943b3ffafa1d882db71f0624eb75fbf0153dc15dd2aa2c9caf166b3aa5bd07f759a84452725145e46dc391e497006012a18b858b4a7bf7c238e93292b75bb5db5fd4ad1ec8641d7e974a6277d1c68c73458a272715c45c8ff6874979919db1eefc5208c1d368558a0a5879dd45776900ad8347582f5f2b99b60f342dcec6cbc134b1f82a2f277711e0ae435444433ddeb33dfd06a7e4a51327a0869e68aa8a8a7287648e92caefa4e0eecfc3fab49c0082e24723c6dfd0571c4065ba0fdaee8502a68f2ad036c59e05f7311a2c66e49cfae25416fa0af021c4c708b724fa20630c700504bc6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h1f4ce85645524b848a711ef2e3ae9cb7309ae47a45bcca4a4ce435249cae5c59a6fe39bfc6a0ddb40aae35eecdf9ddf85374147a191f90ef4ae72b7e029d143b79f03ce1d65d59c5f2a27968533578de61d1ace7c6789894e0102b18b50f4dcb1401449be668ab78927dbbd43e6f75c82c720945b7dc79283d31056cce44afe087475261861195ecef73ae8d9261e65b9cf0a270c45e88050d98c720c8267a81970358cac45ac77127b32f13fb3e75031ae5190ae302c2e43ed8af8804b52a2d273da13b16b8bbb5afe7cad64c60246298fb82e5fac7996ca6b059a922ea085527ff2cf709b1f26a1c03b76e8123c7176d0e39dd69e38d2e70900bfc505503bbddeb67574049ac0c985a002a90acfb48666d0606eccca95849dcaf129db05475ca47f8218feca7ace555b4fd6df857203e9440a9139986290cf1a36309716fd6fb5b1a064f1f2452066f6722682bd4c4b776429afb7991d1fa609ce057ec69f3f0c60a65954469c9e738d86ccafc3899f605500d44fae47e16dd6b1a106b87f77f683db731946009db080facde47b4dc98f21765b2043e2714dda38fa4bed820ff0aa092a299b2512494fbc7fe815c8cf615be9a7e47c8d847b60133e50321f3caa9eb53d0d6dfe7b4c464bd6d5de7ae036e2039a1f21ca52faf1104e824f83aba042f66b7a8440d94370eb584377d8197f1ed9715f2517e55f23e48ab954398358d425af4dfd2093a3ca4c92031cf99145baaf7b2751fccdcaf70d04069f619dc17b7107a6b44911248761ff63ed91babfc9726c70e4391b19266f5738d72ac75f883329f0b07754712fab8e029de6bcdf971cf35c76d4576fed4f3f7cd52620cd471fba3c66055f5cabc8a0b2e73141d1dbf26cd5f66ac5dd1f0edee892c968eab35a471e797181e0306b33ae5f923d189f557440a005dd02f02c124570297f7162c98459dc7e73cd8e42e5e2fe90fbdb11ae2d9f66ea276024783bdc0419fee723ec83c03536144e970ac9a49504f2651e9a5efdac6b3a351fc2fa8d1dbc6fc8a39e9e0c5059fc02cb8a05122d4c5f0093a21b5d9ce75f8e77dfe88e42659f9f0cd7972eba6f1eab532047f963f5440702bbed69438eb5df2e1d012dcb824f38b43e2b93c05fa598f0b030b786603b852936a0ac9b72e4b0d97192161c85be5c3dfba7892eb3199bdd3527095cff20edd032139b5f0d94133373fe844fc7a70bd174870259a6bffff48de2296ef41a5c9dd8e3e81aab7bcc99999eca0b7f5e576ec519525f356b48db0b6cd83575b453f6ada77761738480e3acf09453a9ac8df64a9a6cd562c416fa939733f7480f7d94d83054e550463e6cbd5a3ab0eea29d25bf08c0e48a3f99a07f4649b3bd032994010d39d86a38c80998379e71f035efdacfe08eb70894d28a1ccd3985ebfa1cb931c88df3c9c5fe06552161186d617d9e75a9a1bd58df12fc14bc1431f9d5e1744352bb0e0da892726a06fbc91c379e7bbe32141197f5fa08d889dfc93c77bcf3c7d3c2e4dcb4a7600f2d24586bc6551772e4b72e9dd1f8d997a51215bc76b79ae68d60cc1b0911f54a09823f0f14fd98a35df483e68702bab77f8c66b75bcb19a74db8354d6c004d6afc2551371f17f65b3e6aba767d69b11a16375f092bb16787304be897882b7cf95aa351a8756371d11ef6864d2568e9b5fcc13ac267aacc02441cb56ca26d00b9aad1d690ffb9d890822f9e42f6cfd79117e659a639b323ecac5b1a188ce145de8e3a24893bacf7993f6555e2160d7fc075842eba0c304d1a0baa59afc5820303e8d8da6694d5b282765ae7e7b29f398c6635120ad698497d4640023c9d6d16e26333520fdfc7d68fc99451bdf3cbfa6cac6c857e320886132d44248098a0d178afb9e1d6472c3c0b45173e7855378c5a9769fb2f8d78ca1e6ff0b0eebb3f6714f17377d14348773373be53d5800767d2e94f28f2c2fdc708f9dc85f82b26c5689402afd085298dd5cef33f992c971410f7cf32bbc553d1dd45071cf10afc10fb32954323e848847e417d9aed4f3b5fa0738aa5fcc781b705abada5dbd17bb90a279fcc614f7a6102a460cb81cf566e341cdc3e8fa4d4a7143b9602c7fb9d205c553098b659fe6483a232d43222f8de88a7771ba19b4820588155593e13a832c8ac94027713603910be0a26d685f78842de0c2de6b0d73657f3b70d50a3f01cfce72740782b4f87607d390e6b85d876121bdb143f409807c607a9db302e8e69d74d30e90391b3b1af38fd8c1c9535a1b625d0d8ce995c29c843a1165bca86dc3c0dab10787a231901676c490652b805af6d90d8dd3bf73ece5f96a32c2e86ad9c7fa475aa504d2264865e217dedb57bc76fb70bf84eb9c59bdda192f1a44aa18b5ba3b9f867eabd7753e878545e149087168870e5b609a218ef85cac56377ad17451594b04778501ac1d57b2f445d3b7ddbbc3d9325809d4a5cd8dfe1a19fa7ca584fadfd4a9384bfdf6f5ac1582b2124fb2a1b5c8fec0b5c624acc1d81948355556b4f085949131cbb5167eb69cf38791f14872720f4b56b3a5d8756f331f30e12a9b0e28418257749d458abd5d064afbdf8dc7b8d9063199df074d533bb5088091fc9093650efc6d827bdad4562a2bf4c80f05d5d24f19f0a517344b3f3cd9b3fb618819036751f29ca79a30e2568e143f2325e6756985735ba8ff99758af97bb89329c63c1f6eca13199d5c79176436c7e90cea70851fa3e02b6f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h578df4ea9b1119ba5f98fef040b8527285733eac6048627073690706aab08ac7e2cf69d47e45b22c8154c9353b72fce27fa618eaec25878b10b491a5325fa9d0d881363c96225ec24a36a794808c7bb2a1a780c42c38509c5816ebeae6d317b3f5df0c92bea3597200dd7ebee5886cb09b8fc84ae0eeca1bf2f703898142fa0e9a1699ef8101eeb5ebbaceffc104044957aa78e446fb1bd52b40ad2ad8126b66b515b08c5c37eb611545d5452895a1a9ecace10bfa70e0b1ff592af528f9d92d9632a46f224d08472f701cb10ed75bb30f432a4106e64513c6eaa2c15e2fa3cc1857a4cfc5a23cb01b986ac8b1300c71116e952b1f20dd810cc5149e5ca24466266914c68caecb89ab119d7b0c7c54496c0e6abe6caf9638181b8c9d9ea3fb104f743fdd4b974101ac5544b151b66b4a651b99c9f22c7b88561a839bee22522fe5fe3816f1233fae5c01bf169f51e6e14f6f582b2115990e63cda4e4971d512df3d6fdeb29de66b5b1985a23eabb4c6148d97ffb3e904222ae5a764a1f6bc105debcd8e3df39960eb59f1e30029bed34da261852a733b87e551acfe2d5c740edcafef3fc16c0a16474af5b434f180ab8bd511782b51e746534eb62a29b583be5b4ec88e8287baf475e22a7ee72f290ec7952175c4231d94a208ba00258b257428586e9d5f8fd3397db63a2080dd6be083ccaa37d96e98e4710900de375e3689697e1de7a9182cb2a311a38ccaf7f26b9fcc7ff77feaf5ed3e550ab05a683f4124c03d42b76511cfb5535ee4de2470e8e7c8c17f6c48a05efd28147854039041a5f1cd7273e971a5127663a20253ea3bb7b7fb657617a4b9303c21a2a5f5fd29f14cb8356271d6463847520be1fcc084a889dff259f128b7ea2c6eb140cdb986b2ea6e8cd9006cc2d2caadd4b26489d964b97bb2dd1916060989c77d83ca50a17dcf84dcc29dfbf8cea397b62cbf71020134d04956ec3d352f85a3775094dbf0a4a4db2723d4ba5ae91366cf80bd03067af5322b582b6493179c40deced2ac376a0ba913c8a4d5d541b2fb7850c823799ac5390d70a38e685c286ced5edd9934019b087ba66af1e67bedc178703650c23e7bc680149028ae08e8679f41f194acc5d5f92e2fc6abac9ea65bc8e3822b0b2ef7913ec45b9fd379998c6ea8a353c5e4a9857f46e9d68cb9f4f84919ea3cde0c8616531b5284f36cb6694b97db1339d3a135d763bb71ebe53f26d3a1b905b26f8f6d1fa597cc2c213f8adc76bf3d4cc610d13d6e04587fae4b1459f60f0a23cdbcdee143522edca74a98612fcb9867085cc988ae7c5ba3933ba21bedd641685ca5837a7600b61f98307410500a426b6ad56475f1f1b9e4df4ffe944edf4d5f70c567c9a00701b83227251c38e9bda0187aa2c5e17798604bfdb2f883400305517cb6af35471475c7e4ccaf439e059515d660bfa23c70d73964c6991b63e9c66211f6006edc7df31887d0de39ec18912011028e0a95d26343210b858686ee9f1f3aebbe48dd69e2d90e1700b4cc678d04d8eb0ed768524ac8375d2c8b7fde92af1b0a69ce42ea1eabe4bb4d96ea368889f6ea26937b0a389c4247da4c7819febfcae14216fb2284e1b84bf193f06aea540249663547d0ecccdb900cdc97ed5b2672ecdbd1692ab705d94b45582a1973ea0525da247f90b4227bd1c1eb4c4c44eced042f11f76f11009a06fd8ced0aa362f8c6c9c6859efb9803168183fbcdf5ddde6c4652b0013ef73106b4ec1ad92b584f5951ed8d4445e9edb547abc6306ae326ae1e183bfb74fb512a923e06ef44a445f040f938cec300a02929937d8744e98847714b5531e483514fddc68e19ea0a1a56970304471e57c7221b00029d68ccfecc8f2adfa2bd3354decfae585db12fe2e1772cdff37b2da58306e1b9e25ee7dce957f2ae1a54a4a674cdb0996f07ff4a0b9d286230ff4de17d3b19bc7f0990a0988b29b64a3e14ceb9c39337e6ccd56c1ee95e495d80c99c34a06e43d18a85659659ce1167f9cb2e571f324b46336ac68fe3df74795da85419df356d78d64cd2900b48ddbf6c2a6703dff11b06a9599cfc096e978f37ce42b4a698cea9d5d2ebe859f8f18204492783289d592ba4f7161a10dac9a0249c2859a3f0d1acd245bb958bc6de3ddfbd674b666af0738b6a731a33d51bab13b911a5c9b0cad564bb6e1f96c55d07febf45c576a295564208970c9e411e8c914a4f6db111051d0d907d5ae63d9ac8a167754f1ae7226ea0fffb0fb40a843a980961e2fd45d7242cd1f20f9a04a7ad7ca017e7fe1448bef813ee03ac66542fe7523e541a43302e6800e51e8625a2790dbf16c19a87ffe5bd8482196d55a83e9012f2dc3156c39e2ae9ad6b1dc92f4da42bfff983e9521e0e7fd8ee46b32ea7947646c68440cf3e069377672d0e401165cea897622caff3e2dc92fcf1b1366c131c23fcadae59bc2cd1a0bcbbab0b07847973b9bdfead50ece6485675ac6f06d05e82e67929e5f72a3b5ca473ae726a2d5dffdbd99b958e4dc0b413c95b5184914d2da3cc503024d637c329c7725601f154d4d651522040a54fc4d8140a1bb20fc7220f3dc31dcb9e054763690acab70ca00a38461b097930d0595a3465130235c9262387ad10c5c3704c5cb659f614071925d9b6a42824cea9f0f2d6061e652b704086dc512b7b2b41f6c00e27e4873fa111d0d60976adf6a970fa21d8b2b38e4de52456cee07ad3b01d5316c4426faf0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6661fe0982e79d8881ebd9a993b241953bd7570bcabef29c452edb3651bdb0e03bf92e47bc020bd44def7fc5ef857233529ff256007ed04651c03cfae50f97e4f5ff5fe72d18eea97cd69d194aeaa47d01e09e8282199911bccbacc2abf766faac2a79d0aff8117f1b2cac1d32cc05611a3329ab54d7510b3c4cbd6ca9d1fc9e5c7e4abc94fe101c548e078a423b56e5c9d86fdcb69783145ca1e56863dbb220ae9099aba497920e7b07992c00c72269aa5e7fe026e3a90e13f75e386ca3069fae1e5d75f2f74314e8a1b056b7d3bc08fbf03c7cf32c005fa47be186b9b8092bcd882fa399f67cabdc55ef142d6acad70bb0ae59e491c510f8dd86c1b107075ea4b3b082bc85b1c3e58b7bea8f28f53a2f6edad4e454d6782bfb1539d2a268f508e9ef70715cc8ffbf691fb3b41ab07563c4042feedaaf0a0964ffe6b40b127592e2a0840f963805a4ea5663006978de76d7376fd678ef62fe6691c425b0def2883222feb70d06f0bc8fb0dc7526fd200383cf665f095a54627dbadaa9fd65f178f8691d78cdfd558ae10668bd9970abac81848d146ad146063456ab0f1c75bdf17afff68a0a22eeec35d0004b15c148caaf77a32eef3b3373e29021c6015a98f01073eba99eef4feae8302ea9443a305287362b50ac6305f463d6be01b0cca3e4159a95c461d99fe21252305cbe69b63aef337ee59cc1b5324e515861054418949a268a67a7f7f459c92af848c5606b98dce27ce865a8fb79d22567f0a10a3ddbcc1de4b0a2038f58b64d91d0ea2ac3907d2990901ab8170c3202ecfda0b1835004b2bbf0b5e430f21a83201b22c8cdd793ffb14e62e8aa8053539fbb9398008cdab4afd07d6502215eddfae182f42356e2f88ce2f81617a61c22dc1a87df33a3ae787d057f92aab9039d118398c616edf155ef76e72b7bc559b1a55cf16ad31bb3463211b4e53d8f9874bd9cdd90ce61c0f644b99e935f6768bace3d67da3f10576468ac65e283d9b8085fd112537f9099a4d298d996d513e8f5887b26f49c051a2d16d7274664584dbd59092bceca679c8ccc8eb528ce364d6743b7e95e5b8c253bdf0fba3cfc93a306295adeb09e573f1fa22aa574a2b5702499ac3cbeae3867713b65b0a482eea26530ecea979557c7a8d7e2f7deb1a7664d8206a939e33d9ac58db65b2b13bbac3a3ea0ecc7aab0aeea6855e7e4abcac948a6cb3e6de1b29d016d67609f5d0cee2c59308b00b5bb2f68e5ba1928b8f4835f6c9191bbce43d2b95bdaa6735989700b6b472996d90bf65594992d83f93c0a5685dc62d1cf03183b971d8bdb0fe3b44ef6cf45414ba6f2075c973f7bfacc85ff848e5751a85af326c217097c6188bc4ea57e6e64878fddebacaa6c86833715ec4d21cf9c84c0f0d561eca0c03b15ebb8b0caaa6d9b7aafdee40128b9bd5891446e476aa6024bc3af6ef4e9362e5de2ec181df5036fac6a68cf15d38d4696edec3413aaed6667355201612dffafbf14ba8b962c57b83619fe916f78f4575e3482e3da4add3c11f0ef425f34051fdde8a1a9d2e3480200359b52f7350d95277559ad3a1f781b9f84d4ce165a3689625094fc18de4e2007a55ab9376d113f78dcf88792c072a65f88a8416170fe9d246394dcdcd62142f4f70c3ea3c7aef62529d0fc985d6e4fcfa25d243607e83016232cfda55f5cdfcf521c264e8f2659b0e247dfb933dbc3bd5b7046efe5d243d40a20d7a80c31d3fced4ec027ec21c2b38c3246788b17c28c07a5f2a3476653fc44d6571443f51159a8b8f744fc23940820ef048e2f3effea12610ae8aa2acc4addc7a5fd968ff6ba79e8da31b9fca1482c1012ef4f2ec5a63b64c021b09541ec3e050a490705ff8b7bc5f7763087fbc0559ced5538a8b89995401e257d8da1936cd4d18d73c0367ec430216ef6eebfc9abe5b50ec26d96a1a04d9aafb002ff095cad6a9a822630290354b2b14dc1cbe237a706c6db3aff9df2f1ae8343eecac7a72b928d49b9c9c1008c41ec8a3ff21f2a10c50e4e279c061fe14a93d76014de5550731cecce9f2d94e3ea42246a62d9c53ed6ba1ec41f6a36482d13867f3cbe2599c30e3c0f7d944244214dfb3ad8248f0f8d2c1a3152492f0f42c149cbe9eeac636d987af6fce75cdd613cc7023851e6da6028936422bcdd7cdecbfa34cdeeb176b3c44d71326465522ab4ca18e26a857a070ed09929b20d73a99c61e74590bea3382dcfe74aae8998aafaeb505bb7b79af43f34f713a2984a9e6ac6fc8301f691de130ce163c9293f584d2102dc5c37473003601cdbffb6ac1878a197b8b1e3acaf73d8934eb188c28f58dd8912b8d83a79cce0ee9a4757d09fbda2a971658820c6d03feb0bfa73ec0310dd2feec3e81676fa460720b46f01cc5a382d46dda5f86d6de768f986e85642b031886636afe85563de9fcb97832185d00503b866d11f26cd30d84cb5b79babdae9d35314008167c0489c388af4b6b41b30c676270fc359d598a408869d3a74bd09f99b665b0f2fed04a0a5930ac24051a9ea2df62a5bcd1d1f2e78c4703b213db2cab3a8547e830513e65f44c9c30dbcd863beb637c586709c35a1e399cf8dae5513d2a3c17e6cb3a1a385f5d319259ecd44c38cbb94f9140183556a931f506eecdd455575175fd5810112fb3365614172d1ed77ba2140f63978e5a61115f1497bfe11d70038778c1346cefdddd2fd7d69a05add7e1140a47acb57298a7438f32a83ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h5ff39f38c0777c2f5682cc8912de344f278816b87235a60680e19dcdd49efe582bc6648392544169ca20278629deabbaec9648aeb3594f1ff662d028cc998e574eb21561bb63297d0ab70617d04b5ea91696fc9890f74d83c5c9a4d18d144287163a656b2e13f9057b5a83b4706fb4847c928c65a1f085e37cc52ff767bf7e6b05cf65cdf7fed7fb08fb0738948095e1f3a2bd14687ac411225faf2518ab224bc93168e27683844e784f000ed131a7a6fc7fa93ecbc5c7137edb7213393a69d21413aec9c8fd029c098c7eb951131258ee9a173eaf18a365424237d8ed230ac7a0c2a249ca6ee3b7ec0ab5d058d99e4c9446d90155f29cb2958d9244d6425453c07bf96075b43aafa4c70123c44b8a09bd1ce8ad0a13a6e5b18ef983d89853c6a97b07d0955a1e13a998afd9efeb0c35fd90c92c431c682c35ced6e6bc2d62b5ece871c5fe53dd08549eb9e8847c17c8042c84e90bfd89ec8baeba0ba5f1eba57151f7bc1a5e1605d381dd0c696a08dafaf769d73ebb2fec16666190cf37b613f289648378d9613e33871d5bf0ebc9dc7145913502ff4fd4e131f6ddd82edfba88761d92bfaef0c6e371e14ace46891c070ae030fd2048e2da77ef8519aa936edfbf45ce301bf006427ab86996706f499675217c06dd54139f5b2f8c412be79c48d1f3340d3d73754dbac008d66543f1c5db6c37292e41ae3e2b38f2673073884378948167b24f30bb00088847e74bf026bd564d03fb5b09d7d5984afbd09bbe32162fea6f18542a93d9afef79fa78e63564e4407f83a9ca220766f6eb9bbf8a8b935481e4d576d218d4f6536a9770ab46148b7c47977375fc10df4a5783b03cda9a5d848bbc95e1e79dbb170b90739da9b435ddd0bc3ad4a7aadde7f8b409e29472200fe0f6b8bf95a585f67488b321f239a9c87c2e1c72931ce011b0150d4c6a329769fdcbe1641a41c71f388b0cabf207c0ad5734ccb15c2f749b20efa62da9e513437f9e38e67dfeab21c6fe36103aabcb7243a0a1587df125abd5b095d150f44ea6f735331c63451542f1b0150be597c657864f94d4c38f7b7457b5ab007a5fafafc6d9b76619c0257a4502f03fa2754ccb2055342062f166b8236001d3352febe241d5ec2fc4a6a2d52dbd6bf7334bb04ee07a42f30d6455e5e136d673ba111268e56b04f0624d3bc1cd8929bbb9b7e4bd8ad1f425366a46b4ce60ab270f79826518bb4683221265f65a1691f9815be12851b2d34d5ebf5e576d5b35d2fdb10e466570857c90affdd54418188146310247e8ad7e8f8103be5280442ada4afb24e52e97644ab81e008e34f9ecb955d25e84b47cc0dc56d70ab8ee116ad83d4966e24aae28607f3dec6d9d77475b151d3a57035aae8bbe4075f41111869d83899e8d073aa502025392fd2751070c941de429b61fef96d53267bdd9270d6054e887dcb408ce46938237277165b4fa5e43c6bfe0b9e9abb478cd4f56eb75dbeff8863bdcb7a166874e264eaae261a3ee05f13136821ac8fb8d16915e4d744773e06471f161427c835c7faf598280eb8c6893c8ecdd27c549bedecd67eb932b89141e0378f833f668f95cfad949879c4f89d2c3ed30c60c76552e5053520fb311a88e73d9dacf299afab2557cba8d19bba9b6e9b5bd5fa1284eb21eece788f76067c85b22d4be39f9ca3d73da3e49c4ee59bcd6ce812a11168e7ea0d85b80a57a73dc9083ac87bb86dc97de8390e2013751d47021e242cef0c2c44e03ee87b8a50304e2a71f60391742bfb0adced4ecb28a8cf782b2b83c8bbfddcd7ebe9948d4cf828d2ca9181ee0cc07a10888b788be6087a4f748e40ff9b58e5dbca0f44d05643c5af48482b0ac64cdf68b23a78aaf18f3d695de46cf2f6a3d2ef4bfc5639cfb74d3ab5ef5e4b2b7799104125cce884595391f8771712dc6e706f14f6216a9abc742fd169df3d8d67db3a74ebadd9f5444c81bf6f31b5c46225dd7def2fc02b9b74212c7afe251e318bea4ccf2d45984b845b5de6dede2f5c7f6b6c735ef64bc79335b84ad4af1db01d8b81ec48de6b04a483fee08d6078096a848f79b5e5b5c238eda34d4df125eb39d3fc661dfcb414937bd32acbb6c481bfa772f77bc1ae070fe5f69ca952d7152a5aaef639653ad96c1359e5704a788c2c711782301bbb83a5eb407adca584bd74af2d9e42d2ea55efd434f5ac80aab792f3227c314c0516486fa2cce7f70fd4719feeec107404e4f5d07ab18a83ab62a64afbd4e0a1f9dcad0fb9699a07d3877166d58606856a5231a9db705630cf06f1e04e914c0676fc2d7862bd57153f8b5c7ee6118ff5890b6604415064f4a25d4896c9de75cded9b49cd57cfc62600f136df5809b62861ffcd0fdecad879bca70fb542c4ee18e0e3a1450cb5026f0d5485b1696c085bb7d483a5c31f9c45c895f5f1be3ad0e3a1eb14d0e5e9027ac1b0accb41385ca9b92b1b93211471f97581dbbc1885570e7e639d889ce94d3b310977a8e59570e01509801645b6b0410739c5183c63fcf70cbe4dad34ef9e3b744933ece925dedb204a19b6abeb2344063211327d24cdf45033519ece098431ad22950f2c61c65d966921d7047132d19214f3576f4a2ef72adfef64f92ada1c995cfde6183b33d2b4d9ccf94869531e08acbc3ce53020c3ccc6355fc7c5219e5e90c2710220c1785d000ba00a530fde7d596eaeec6327c6bd78feacbe746049ddce72e1e63fe9dd4ca1f2db9f3a0f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h9aa871ac44db07b0f94716aaa8fadb9a5a4cd15c7af57c43837100659f862c68935dcbbc5d6908dda976f8c3af55db9c4e52516fa3dab5b4e5502af45b10df1ec41cf5a9e06c63eb4ac41e3c9d9961447c67cd67871ff6ce42f34efc90ec28bbb6c4692c9d667e1db74d27bb59bd05341246faec9d4fb4f75315806b9f59ba5227eee354d69b7bdaca455694b412c9c1356a2e8a6563667fbfd5a566fc2d09c62572c7e4dd231caa72095a10fef57ca91596b21b99a9c89c5f62d24b3f49dbb535fc63448c31f06b693390309cc509a8028c4f7b09c24899d5df8058f3b29562a30068d98a2d521e76a7eb03444ed8221d153e5d9b5fcdec0cf1f013954a86bf811382cd2bd7f4cc443b1b29937056f39febcbddbff306e0138c97ccdc6fb7efc723cb7d9af428c044d3c653c25ce02df8a2c447c2c68c940f033ea27b823694b67c02bba8e564a662c955a0273c74d6a84844ffff6d62ebb998513b12d45480f6a7bc454f16957dfba7a680798b323af260a1dc642843a08893faaf3afec2b4ec6ac258d65f2c4a7dd0983a365d0e825a541531d177203df8ef60e722b8ad9a51d72e4845b55b0a375f1fd5ea450ed493c1727464dafb0534ede6ab64e1796a0c6482b4703688d280cde779d54a720ed4493d45ee2a1cbdf55a1a4fc408a1e62c0e5ed375d94a184b420a7dc6365251ce3d16c8ca55a0626ecf97c63220faeb7c2ab75e49809f78ce650149c59283ba46718bb6174f70d341382ee3f6345f361fc13f29331def0f6b810ae285b51f880843ff8d067015c5ea8565fd5dc7509531e68349f09f08632c804fa8305a0e5d398443b144f8a9ae6f33f5c22bbe91499334c33473226f8808e1ff42c2972f9b0b3885bad6b863685352eeea7bd5df9c22c1b998de82b676d1c359c4a8d82062fcd7368174331f0c45c6ac11991ba7513dfdc78d9f4a6024c74d53a08e340468311eadf63320fbde24bbbc62442b331f5425cdfc455583cb8975fd6227ca62b5bfdd6b8ffea8a42e5b9857583c508ee4ccaa812cbeee770b65ef9fb729585c7ae19311bec75ef40f77392c4008116968751e1e539461920a7152b8bcab40bce2c3f739958428f8dae99ff5fb888648ff8e5bd4b7629c2697cdbaa6c7d0c0147666e34228ece4fbcba76187a8245435721f7003a8172176e6d06767cf16751d9fb55881c176ef044b0b2327243645a60e919e5985d832aa91240f91e3e05b3ee36493366034a161a2d9352fc2d5560471a2203be0dd641cc077e8159e4d0fcb4748f6533c6b5944e8b33aeadaf119101f14e0674b3bc14609157c38837cd21536a60c287b33de947edeed43b27c418abc320df84bce0bcc6f481cd01a3177d59d9c85a379b9c81257b490e07c6cf56e0892493fa3ca1816d3dde06e52e85eef52b08a918e4d1ce2c4e179a409564725068437af425de23d0a6bab879687b9c5b95c1aeeb87a1e7ddfdc8e18b301dd2edbee55964b5b6a6ed3b7e2fbb52ea9ebb8c12f093de1ab3b9f6d3dfd1cc5cc21f2fe4704ccddb707dd41c2f375cb6c60035bb1f3a571a612458fd1231bfe03ba6162dfc536f205822971dc89cdc490785ccff094370f51279d9e7be52b54b2422089bfbe220290217c1c9c09a5f3dd9a5576c8e9aeb297a1e858500e12654d62233bbe625e8d891c6af69cddb075a08fda33df225bf15b8640e2afa3e9de512de8683f98ab8d814d37181aeb00766c2e81b25875e7dd6718e77a6577cd29fd2d85f5ac49f088ff82c08b88cd04deea836559d480bdd2d8f4699857e386fe76f610b36f2714af308e46e8f423ca9ed9e8b8afe4f7a3a750e2cdc791a20fa40b78b39d0e3ef77d926ac88b066966256dceb95baa3805c8bf3f30d1a8771f79cdd82748d474dc0518664a7f87dd498e6232b3661099e7e8c6de26d3c52b1acf80ab10d9d2437dcfe61df55f7de0edf7c63ebba10d5edc998eace72aecfbaf00e6c6cf1065b58a9fc7f20ba0d5b63a8b95b5b8c2f2d3342aaeed7a5082234edbdf88e81b80759d40cdabd800ff255c1623339705f0fd0e6665382dbb86af4cbc40fdf37ee6c5a067100c8cf391bea3d34fc45aba57a805dbd9fc19504feaf00e398750bd5a1c307741314d17f9182d220bdd736566f0f7ec52bc3b2d2277fcba70754a2e4413e739b37327eb0c94da82fc429baeb10251e19b6c54d3a1bfffcc8602517bc7f7ed808762d079933542d1c19ffa1754f8b342a520a75b2f39c6ebf1b4736fa7780e1c4e056518e373a562f397dbe4be8325a4d11b34d54d88e8dbc2b15629b0839ca60303fced4df274c1e87defc0c6e3519bab5621df2a4bf23a70b8c573f22fc3cc10037cacc5418d05e4ad029ca080b2349688de74597d6a31f75b78e1e8f6050a4c3ec8a04492c7ee48a9c7df8d236e0beae4e792a85bdd53fa6beb0a6dd7bfa3aa6677649dbdf1ffd1f2df9a93a5715945d78895e16cd3b6a59f89ab8c32d4d3d43955495072d34abb5b84fbacc71edf9163fcb1497546c1fff951a2bdfad87c6c0bccc082a75d90ce90fa9f75bdb110e8c646b2c664b514e2cc379ca18e4408dec258884ecbe8ed81530fa5de6faf5d9469318c274cde5a934cfcbfabf98cc74fb9a0685db260e5c9d4cd75eb8da66a959a2b5b6b669b32c2659a55d7f24f9ec50893c831531bf168ac0495818ee7fb4e5fa0e9cbc5525304e126615bd2dea34b3032863f64c6188c9e6676d957f8dbd69e19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf3bcbda600b7b9eab9a90227d5ad9b2aa053d1374743d4a044ad6becb3c71fa0eb10be9885997b181d433011c9e17c809426c5abb41d67512ad9c08bf786c239f3445ab63647f716f079ad62c693930b8402fff8bcd2d140cca0c60cf2b4f5acd4a9c6bea3c994a4f0e64b8f6be981638c5d2be5d39395308f700d59107f6b2c5819516c09c97b646874a4da6a5cbce0d7f3dec5719a94e1f5c0414f0a3977cea5496a89007905d15cc93ea5ed05ac29c9a559a8172179863a8e273218b6bd3f52f604c8c4821ff570e5bce961121ca9f63df848a5a476607e564c9b19a43e489811819ca2d7023d548714029bd746accadfb6ba798ff9eb766ed0016dfa13b0f729da40d610e0280592ec40389b1beb992d859ed034521bc2621d8f5bf9b7d5600a808c8b4a602333b29aa19560dde3f9abb7140ccd93a043d5b6ba788fb7f002f9e563c4c22577dc93e2fe086ba1ed5210cb2c80ed605abd8d11b8d2c14d4d95307ce78708d7535c6a9ba832f5c6cec8b327214f0b992aa53b5a775506b6e7f774d250d2d000e9d4822748bc053b39e0f1db536d11a5838118e063ef01324ac1ef372c60bcf9b00ce8a1d1a2379abc4366946257389248777886f0cac13326a597694d554dc0ad576e6d48292c2e67126b922479b5ac1419819121c7fb6222dba673e796ba8a19b0b2d2240b9141595c376b673769ca49a9e9e83884a3abab1fc25e33b2a13565102d98a19338786f1df0be7548fd9e692f45b70dbdf1783a2c70c945841c954b45a2d0ea7504caf2ffb4ff710dadd6f9bd2012443e549b63f68ebc335c30787fd6f669ee40b061e4cb35adbf8832b7b16613b5d60c2394afd64ce98fb609bae95d88f9dc751d64788399e2875a64463eec3e7f3bea84d71dc316672b895808677c1df8d28a65bf63ee789316bd5bca3dfffeb7c1b52857a0488fc37c35c274968864ad628edcd87ff11a2ac6e211a1a90f48b6d65e285467e7d9f0825809f6193928655e334e94545308e42ae7fa83e6841e696db5970f7184ecc63fe09554b4c5a39f556a3650675f797ff0475f69a02f8707043ab42e973606e05b612c2247fc288e34a77f8e97ee18566d2e87c17a502c3c5a0bdb3b5abc0e75811d9f78d7fb0d59e4030a6f6b264405142b9f9f45522bc5553bbbcc6ad8f37cfb56e892c03959cd239f42cbc42de72da99570a1efbf01ca59c2e78d5c7f33175373891f3ab1f5ee22d375692bdb5ad5cf4d3c50fada65ae878fd2dab89bf10a885def553cc4efbd30209c13044d430536bcc5b40e7e6104fc5220d4120e7d6568c9d20546c4b2c9c986a2c3f1622e06d4fdac07a19e9c57bd62923077749605bda3ee77b42973e75296f09bea5a821b9d41ad5ccf71dea38b4ba1fc562cb5d367ed67fc31b9de5252c89a8ef647be6f2eaf8d5ac26125b5608fdc149aeb6da45f1422583a287408a93f02aa04df456464b0234998f7a9bd21b66cc72c32dbf288418ad25eb929efd1270fd101000d9a72d9fe112d2769a73a211771c1d5bfd37a2f605fe9291ee9c419d086d748b4bb627bebfeb749d5c44e5780b9b5cbb9c45e58a314d9fd1f9fda84f41bef32a7f906f5e3ea088aa8cf05a28b3e7a081593e43badb86ccdd880a459fa0bc8c5600fe091da46ca17c54ec71e37975da3f915ecc61185a72e4b716ca1504a8cc8dfa4a5289cb49a76ff32aa82b9f43efef36c77f74804449be1e6757241ef9dc4c28e72a65319a5b1020c1d0d9040097f7b5054174e86b98db5d08423c3a53de7f753f7c297ae57eefa5509684e411df2b6b3a557ee5fcc7dbacb12867aae49f743bb09c7a53e5449e5444be128002497e3991a4ca527d489239071f246dbb0635e5000ff37ec79981d055e320176521513fb9e47407c4c03b60438e12e3b0604f857dc8e478843f069d889686ba8daedd6a485ff733a3e574f5070f8ea0348bc59a7de2fcbf056c8884a773cb8ff5beb9f563eb40a0708341e2805adf772837cde57375e4d71320a261ed69d29323e028ff3b8477ba914f08ce000e406381fb0b870082f63b981377859232e2306390f2589611d2dbc4b8140c8de0fe8d6667bdfc0b762bc3b11d56bddd3f97596d46cda2dfbb0fa0b1e39fdbe0ecf468f13669a7ccb798fb9c4a4247281ec56522911c029b47876f047c7bdcbed95483d4c1ce8d07be424f473261eb3fee01cf610421d58907a7c9d0595fbbfe70408e60b9f9675521c661fb10dcae1abfbf70f9d31f80eced67533ce6623e995d87d752586b32fbf151148319ceff94b06065439e52c2dc225df26ca8f8b7627ca1a608fb9b781f550acc5985d5a9d13e4ae696a08584873d19af9ec53f6fcbe25eecc642afb59781c80df6688a6623bc0020ad8fd23d6739b3495a95847779a9057845600e27b3c30522e2bbab6e2bbdc9b983c268a914c97bcb6cf7eb2f52956f679b0aaadb778a64e38c95dd29342eafd3689831cffd28543a22c8869ce99cb084bda61711f43d96a46adfe13bd3d07f847a6a677291d0bda3664031a3619e46e547aaefca03ac41d4342bf009b39c70bd4d976c1e2c163197def7c272094818938970e479face91dc4204391a0bc453de4aa3d5328196478648a3c343961a5bf4a938d2368cb16d658b39bfefd1a5eb12672205090feddc2fbf1643f068caaee845b299f8c86c4b52906ce0839b7061fa008aeaba5412de2679379e3e355480b6ea0c6a0750c62644588;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb9f2d08038ffd694a16d0792a1f3cdb16d7869532ff3487432f73b503393f6461f70443e420c4f7b53faf4e55bd5eda11711e514d1489b284eb9cb3d3c30dabf0094f1fc2338671228698d872ffe2839db3147477f0de2ecad06c51a17f8a472ff9f79e0847ae4192151f8b437706a9caf591f8763ac5b418b6ab2995bd545e95ce6072fa6efe1e64c4c5ee36b956da38ab6f095b8b98040e8079a95da6d931314b11c4e9c4d792d7da42a66d21ef6bf6f33a4ba942f1e4bda40919f36961cff0230bcf889aac71034cc8fd230f5c383a3b3cce8832c8a624b7d4bcd75bba881ddcaf32abe05aac5a2f46589ca2f5f6bef1a6043b4ddd58d17f2e61793979a444fa4c91d2fdc316acf7790691b7b3b27eb9a2bdbcc5191fce36ba897c2c0f51b45d5b152ecf09db2000a6dbf84c45d632430ac69c259498258a079b785943c88501df360a669bce22b81314abc2384533aec6450267e58e20d4c0415c9b5d233842aa950c43f5db30219d516f7ba7f0abdf6b20b1e1d74f17d5d32aebe85204e311dd1f24b71f1a220f981c9bef946431e7312d469433923834f320753454beb8e8ba8e3406f40db618765dbdd72c79082ae227bfd0eed115fd0bacd869ffbddff69e3a4f51e5289995354af9858e9d916a5ceee48264bf73f54eb76e73ff56c4413246fb4556651aed4bdca2411af2d52ec20782367a4f958c6d0e9426eafc940e0014da47ac8ac9056d21be5d5137bfddf0ffe55d10899097e0f5cef3be35c0b0a29480e990ef0ae32c87c4f16c6764b76526fcf8e7ba54998d8ea224cd22abb9e4062144f583e2ce2aeb5457ac4f983fbe3e74ed3b7d8862e6342dc09fffd62a02a3d882e8fbc743abb01994a5e61906f7d63dfab449a1ca95fc2879a80872bac96b993ee0e86c90774bf53225e9b08a4afa375fa72650b60ee3caa872169b5da8a2b9aedf00617dc378254f7ecc66328b0e1ba2b7ebe7aa5a1b9d7e5a73f0676964c68097e99b12fd586fe37342f55b01f486bba67e34326fd6ab4b0b3400e40f3dece6ecc33c2f7e932f58909f1b62f1bc7f7ac022be79e12715b3254423f3925b28bda68cadc097331d597b4c21f742ae39acf1ebf9b3da96a8d05a0760fc80ee901590ab325dcc392f7502f335df20984ca8d313421ad852052c69d5abcbe70dcdcb9271d27de1edf350253d86b869c884dd3c9111a3c5b311eb531ca93d01fe9ed5c2df9436110930168c90a464cc2b01626133bad4fe0d2e843b5afa07d59a4fc1a9d7ac9d52dc32a0798dae466a2acad31950dc40f50a816312ca71401f7a39af0444268e81720ee995abfe1dd9debfd024d203867b87fe11c4472d374e2703e360b0db895ca10704bf5751cb7c98afe1235ac71bcb58749b1a57f55c06a1f58a4c8bdfa12356b736f5eef4301ccda302024ff230d76237c6338e6b6f6efa9f753d521700b863c1ba95ce3c15d96e31b742cd414c6f5c7ef0bc6e4391445bca9f3f2bc6c544c1b4cfaa8a5868d756aa770ffa68d28210d7cba9c4762a74148686da951bad0cf5a7376be90d383c6891d29a6a9bd8623286e50c41c786a404d80918d17b745206af6a1945b96ce58bf15a149a03f1187d2e45e4758ebbfa3b2d93f3f7ecaaacad14831039cd769ab2aca631dd57f6ec49af9b96ceb8bc69ed6c351cdb21426ed486e39c50916ceba7d15c62f5f72158b5723644728f7916f71c17e154bf861344bbe8f8e667289cd495255623a5ad6a21b16d225f5fafe7f5a411d14b322e937c2a242bf536e42643c61965fb4bb65e5e521226fe6c88c27c390734d9438321dc8d22382738573440ea163588d569fc31379c696a6ae169e9a610a7733c981201caaef77d92ca0e0b99bd20783e02532d2d2630004aff40ef546e79df9a892d78ad634cb4742c2587ba5bbd595b808d112c0fb926ae53dd16029173e19394af5ae7ee7a2dde38666e06e4724bc8c0991370366c73a37d9313b6543199c2143d3971cda15f751d848c8e52a136d01d74eb9f1b9da6d27d0e09221808e56f0eba6173f0d789a062ff4b916893b5dc4fda026a422cbaffdfc68bf443df668acd9f2851aa7330d79944659b74b4e50064177d9f195e20e2adc0985b6d7ab238cb47aa19478561cd3d79071c315162721c2432a57b37c2953859535fc0e17e060c2e588535ea32bd5b4eb12576935d70cfc630b5525b25e95ad51ac11f8c0784f6cdfe3cc0311516a109aa5c41a28fbb6c74ae172514322c3f173523f25227663575957fdd0dba622ec798959195c52e4f7d21ac5f9fb1e7b7e458a2679f73b74aeb2e0825141cdf7879303af70263d4fe2d93c9d273c8b518fd7ccf33e9294ff56ceed29ec39172986e41eb1bc42c50602f969dbcbab66f0dbbb0a27041f927ee62cc9980adab1f35a49ba32f8399814d6e6a7d71df840b1b0533290efb7b0c1bfc9b537036d99f4fafa2eed6503532ab9bfe9ed7192ed3a87f10536cc56e03aa288005f551b212dac10ff794aa360bec2e53cb8c4ec591287d456803e22c79b7be980606bd357a5c7a1de448135abea5c252a9a21e90fa156ff5cc4726e3df72271ffe33f973d2b210b8b79abd8b4634bfe78ad50f6301706cedd0c1a2e029db62ebf6e0e4c88cb9d5f92f213202c5616554d1f3650d9e823d3613f5cf398f08f4eabeceeddbb05ba3ff80ae2dfe49c682c59a6351b466e962c1e98b71adbc481779c23b27d2d42ae86a00b376958;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h61a7b612a70b6c7f18e507050411f3208268b7b8f5b2c2e514d31405de66c542565e32d51d4f7ad30911180ba08639981eb9be1beb89780cd95847ef47290e46940c023625f3c663cf4d9a16e75c196f31c7e3eefbcc596d6ef19765530be2fc90cc61c875d094942536db9ee4044b4468953dd30a486886a5407c4cb1592b79271f0ed5d41a83f1a7c2690d2b3dd29ed46918fad296f1d664c19f146e276b2a16be11fd08de11744018b7d065da7f166d6fcb3816ac67fe9b9823d220618e2b2eee59828b440050c5ee45ad6274250d5b71506d9e7277fb4ef3f80dce1a3fab7213482fd321d98361c4d83aeaa098c92ce425b8664a642ec3dc925881e57abffbafd5fc5151b2c32da8449696dca7ddda7b797516eea5722bca801daaf8c63b8e34577da3cc2e1fc5f6eea8771fef5c5742b0f20b69af06b7153c565423291e489854e826c3c9493787c9ea53553465025eb99271f7441e02791a8bbcf5496cd241d11e2642c8ee83b354a5c7bd669114676ce27ec97e8b91b42e239e89b88444cb0c7d671dda7ae7c348838393610aa8bdafbf7d1f439bf94eaa6b6a43cd8c9d844fbf4d8a03a2255f6eb2b5d9c0f4ea51dd86f0b28675cbbe88db3ec199cf09e295921067c47502d581b3ec3519d54205a4698c317b4d1a89d59c53c893fc9bb6497a69c330fd831d3e19d315d2f55a4ef4ace7901b04e476d5ab7c6a3ea35da1a16a7155e27be74dbbb2ab382dc8c80b3836280d4ce4b505315602e480a6a431bae57294111bc6bfce7b569410f1e743a1c39d214f4e5760715a4ef740c2884cd2c8f6a89d8544d2284ed5cbdde79db88bee819a2c7ff5ca7f480f700df7f54a749b80670bca23a791f525b5f1c5091b51b9baf31e23dc959b4ff253cd41ab611e411abfb8bf49c6277407b7352fa4bf57eaa5afa1361488c510e8c670e82d78ecd9f1b641faa93e2945e00ffabd34ab5b0dc42015ef13aa5d8bb87ed68a808feabfeb3438c22851a2f0e11976f3da4479b608a0940c75f4b6a09220da8749b6763ddad511191e8d81447d63e1993b7874ad2b7abd9b13a61e745cdcc13cf2cee4d345dc15a2792f65bb8ad9b56dbe0fc9202c715ce28ae64c1518ce229c895947581c431d28ed604849eb01d6a7cc291eb98a0971966b64906e3ab7ebe2f1377202317501bbdb7c8b115555fe09db9fa1d5a5ef56d4a5f4142b1463df4b4e1b42fd8f5d965fa5322fb9c2f46439cfd60d28f59a32242d67fd9c3a93d20bc0182d9f7fd602256d4cb95afdd8c83524f5d3090c206d29f9e0677c3f81f28da99edba002c18dd610830d487fa63e63d98d0c17e6bca18c24aafaf5fe34230008a3069bf3e5ccd00b920644d54cd64a76da8b13e91a67f77cddf513f38139cb217a7025c092665bfc6ae22b2be830bbcd01ca4bafa02ac8fed432bafc04b2d56934ce892d98b428f97250a60466830862336f1a327e78194119826066a99b78cbec2436b6b7defca6badc7151aff1cf89f9e595883b9492e3b1a6ae1ea2c824f004c8475cb035e929426880bde437529e531d9e9b621719ba21bf6967071ffa74fa137066ebe945466db25cb88915c0242b49a472d54b04886471d0b76d7fdad1447b9a847bfd6aac6e9852e06e40acfd3ffc3d8a7ff1f061cc50edcaaa3e3d600b06a16aa24af7c2fcdd6ea841af30792d9b50bd8e02d4dfdbfc99483340e282a4a1e4947e298932a5f68955c9629b08e9ead21b23b1449a0451db51712984cfd5c84c612fe55d04e17fa856e40d73c56d65f77cf8fdfe9c51104f888e2e128c51418865cd53d28bfab8d25d059e959d7cb81830965154abdc639b8e5d052802ef574621d16083b025f1f5305b211ee4a6a3dac90b5e42203f20967aa6ca72b27a1d50565f4b8f2087394ee9269e20f96f4b67a410f77cac454a0427de5113057bc3c8479cc0dd4215a97355f66b5732f2ede8e78971ca66b6740b040d6f9c3d90cee4155b53ddfa5d15a872a77b0bfba5810897e5430206814995831cc75d180eed79db346c3a250b7e59e3817f9e092866d69e910b26f1f2032d299fd34d3e7e3b83c10f13f815cca20b78ee961425785e1491e39605c669a663eafb8c25b2b085f99b0f8df93f10aff04f9862422d873aea77e6d68cebd3595dcfa4da6e7dfe5a523c4a9a0835b704414bdcadcecff2111de9ca50ad8b3e3080dff05e10f3fac154b9e8c607870d8babd877d360e0f6af69b3be0a716b698c6a2dcb6d9acbd9327df4d6b7c94f01d7a687a2ce90948297cb0f9bb56f9b161201bf643e8ab2a8e1ebfb22d144b7413e0a8ebf42370d30f71c0483bd72b8fd5e7ab2ed527fb99a11dcb2ec2a51ab22999be07e167e068369446106bb3b38a28a0e9d49c7b097d510ab55785f4d5383c3949b28f02655ba6232d3e9e3dddea3521d0fdee074271f3d505d8849880db9ea8529141d0778b780acfd191392ed35c45f772aa9aa72af8d469120d2f9fc042096e83f6a5f742bac39fa808e0e4c723e1d0a875083d9a9db5b9240f96c98eaaa392b6420838832ff723d130e46fd6f86eee7685d541bda707a0cc7e82e3042ddd691e58e406d33dee6e4458984c36cc1e7e6ad45fa21fe289819c2ded10bd7f8aee71ede2bdba91d670f4b83853f2d56ee5bba3943198177b72d835235c57e792d8eb8106a2f8043433fee8729a641075ced727a333ab623da22bf1419ee1df0f78ed725dd4f43a85eaf7192e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h3261eab4cf3902ec6eb441e841f62e9e5311fd46770fa369e2b33b412dbbd22415d9b728d461505d25748ffa8777578b65e09612a3d92f3466f7db896bea6793d0a85b13756f010885ffb38a7f95cb1c0d78a3b4543a2ba7806227016ab3fc5f119894269968323b7e8ff548a469def2553835d3ac3c430cce53a219818555be3f36219391ab62dbfebab099e2453e22359e9d8aeaba657f38cc8f17b125a57d80b5eae681def54df5bbe5c5d285d05fc2ca229ae0f961b7f85ade13e3119df137f03263d332b9e0a3df3f131dd0119cea7b7e70b56a6e24de6a13893ef5ef1ac72d4b18ae4e2e6d789bc13513a219d3dfd6b2aad28c5d49b130750853291b451ed6a29130e13aa29ccdf1bdf17e055ecb5c69e3b1ade6c0f53f62fa3f2196068795362719fd49680a3a91728bde3a610a28f9ff995de32342a17952ee67ace43d74f4feb4ff60f92cd0a1eeb49346ec06fb31891c0f87bb71e826e5531c8c798c92da115944319e1e84da6d9fe0dc4b53e695ea9ea9eb077545c95a43ae1a6dd88d17d9f67c4c68ffc46597d8d945c56ecb0c6c2a3131fd09d76dabaa177114a7774d4f9ce7462bb86b2993b979edfb783b7da66c3e3cf7de533d120a59a8a5195a3f0a33da672cf12547693bbf4a0b5f504ad57623877376958d270e4aabcfe8a7c710ac1bc4785f46993150b4410e967822c7c0a7b6ccea14c1b1f530a686de18e4314e793e6e81eb19c2743a1978072b526112af9b06ac96166892bafe56d92a206a3e6315c05d6297b01f18b28b08af1d116cdff9f7edc6ad61db1b71e1cf7b6369b7bc951eb2813edf454d6330664a3544e97437138e3a9718d9f9dbf0a2a9ba76a79848bb0f9de8581af1f7b11e2a9e0ad52bb95bfc6c3dc3d0c0d431b5d84bcda0c548467dc7048fedbc9aefdbe209a3dea3e5cbf62ae486c3e28d8b9f434ec3adbe1c15744d325a7df093c9ae45f98cfecd0854b62caf560c9b0611833ed3e706af9b3ea7e2daae68a9554da6f9340f414109602fa6ce55a2008b011a94ef223cede013c4d541cb999a41c1c4fce0bdb19e4a4d2d720f1f53f3a385e6ea1b1b7b6b5d88695ae64c75aed02d9040b030b2ad6694b6b6e5f7649bcc4c2373c90751add13b3a3d2bc7f0c6612469e63a322cd578ecef8f197a470d4d3919d0ac7e4177a4e0c36a29209fea954714e5dcbdf5e5f0aade1d919c7a4d181f9c620cdc3ee73376bd2cca76396b34a57887ba37abeb8e80bc9953f52f9fe6433db1a68adc632f6c29b86c0c081afc7cebd1b57bf78b0650e4da51f63209bb8012cb4211c3823c29259cc63fcf2d561a8c3613c9daa8bb4fc946d24a109d7029304002bb75b46ec1a861ff80188ac51c104cef17f25ec2eadec5f34472d2d44843e210dc82efbd41cdabe41e48c42cdc08b064b40040441a5d52d5532a0963a09717f18d2e87f0ed0ef24d75affbce9cb7929ef944daa35017275fafda446b04a9c5aa4e778eb58c8c760bad53a1bc37dd8a8101081fa722c8cd0478907e2ece7a7417254242408bdc3aedcb5c36a4f06fb0397da9585a05e71794925861cae54c01178d18da99f8b6297b9d44f064ac01d407a4ff120781d55e5adb3c54f7ffa932b4d9a08d7e92af9f4fcdfdb85d62affc883d663ab0d8e9552fb7bbf326652d56206fc69c4e8756613a7cd5b7a5ddc191e69c08fbc265134bbc5efd9a566a82bee8a662ac58b269fa19d868e49d987fb3f186f7b5f5894c1498698a233d4011be79ad371859ef0cb26df79e0b8952dd85eb0071dca6ab85bc812f4a3b7f8c5030f150b9a95be03dbab2ca3d69536768155219563f7e22602f9bbdadcbcff6e5c48841a6dab1ff3e468ee4dc75ae23fea827b9ff77b8f1a36a7d6e297a248a3faf7d7770f5df6aa0144dd60a0d6a9541184fa63f9db5a71e7b7da869043a88b698a5d4e04f2cf9b400753ac3e2e52ebcffbff2426404cee9177f36c06215f4d219d08ef3e18494da291d5facfed13e5541e67a60fe4e2016d6bd27398190741854364cfbad271deffbd77afb2e83009205b8cfa8a657de6d1fee4bcef00c1f831c5fc0724704c79c6372ceaed8533a33e75f06190d7e22e54ba227061ca29d4a3114f61cecd433c36d2a8cb504b4e3a6ed068c41dc021b1eb714ec86bba6bc7318ec85fd725f80a31d92e25b179f42ff9efb1b4d4df4835fbab2c7c18d5750f08c5ea46414ee9bac62577cdfcb7beba11a225152326e943da452aa14447a820998703d566614f719281c9a163e1dba30a7705dd1f25bd714bf1b8e5320355c129008cb51ccec7ced89330b617b83c42583b49dd3c52917e4d0a6d4e807ad30586f871a71f602bc347ca8dae48fd9b4279119789d2ea67eb1a7d30eea0b1afc7bff2ba053baf4f9d8507dd127d08de81c98b58f48f18036195663e3255ef33c83035763c1e105a99e7ae023dd436d0e54b2e6917d9221d8cb3098495878a699fe8988b0eb59da69327f6f27e388892a16f2668edfa22d4ce322358afc2008282d95ade82dcf79215da12bb028b9161ab94bcf31f931be9fb9c420b99922c6a337da5669dd654a6abe0b18c99098f96547ec4eef19c2549ae9bdc8362827783ed2fcc509e01d362a57e5174af0e56dd104a5c4550654b685510d8539af36b9454c8b178dffdf749f3c9e0bdefef3c5312439b01c9ee27c0516535509290ce84c3d070b5dc1b251f9e80bf5ef61566f70e51c59c1248b0d38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h7b549b0289a593a237155865fee4d2103810787757f5e4cc9663373bbbba4997689de4c14892ac0914bafb20ba21ce526dd5895cca740593088607a66f83b8a8814ba1af7d63a56c42ef444206e1d2b218f18e1f74ad3196459e4f7ff5c30a08977eccf8f963859288db32c6489c1a935854d383038699efb9fc1eae045e6c88f9bcd70115208492738af3285f7cade8a0a5a18dd89610795f797124ef163b52d91cffc34ac5cbdf8bf1c1cece09390f581f024af55d4d527102499bf529528a9898c7017d359917fa6e850d04260b56c5839f4990e01787280a196ad987406f9063fb39020cc8a434869b5eac04a5f3303ee1011003432d5da15a0d56f542a72b258c35bf90e606633a80176d87558e6dbcad85442e4a12bb9affda9013cc0a87d945e8d5d0c976927c66cf0b50da638a89121d134e3bdbe972698760de87a8084feb20b65235fcb77c4e36d94922617c6e8de89836ab11bd636b261fc8165f7cb204ab0ade612f0816f8e3f9b0b5a60948f1db70f70034b7bf923cc016cc6cc1055f779ccb2bf1b48feca902022883ab0aae7af5a7b9fd2aff3a8ff52981a8a5316fe3d19619867858150c716037869657b58c3f93e83183c832411d3bfcbf4262a7b8a8a7fbfe9351bf362d9adfcdb5080101a51a69b33823bbf9412068705b0d268bd5857131d106a227412201d5ed6ad894662cb2c697779a43f33a4e5ed1531e7d713d7ef7179c6f48832befd59cf60a4c230c746ab77c5a99e00404ba66b766a46c3af38f31d7ae0844c5edb3d1dc666a22c73c81373dc712e2b3d998ceca27bb6183896e6cc0ac4e229b003fa292740757040124ee8d20481d5170f8f755437dcd12f13cd0afce615a6564c6a7068bfb5e51b7910e1a46d58b1e393495be521ec99501a9281cd1b4b2058264a0e06ed0d7c1152c813167907a8f9cdb204a70e44af38fcb5dc58d93d2c38f398fa675402e0ec49fbbef0722d9cab02ae1ba4c949cc5bcd16d8805a3883a29f8b8e88345b5974db7e495554935f682301b1bc7927a6b412e6eb8bcb4ff8804d53a32e6de43890dc9fbd492497958fb16ab0023a6a59498f5b1c3dd63dc5f4092d393ac83d70836f147bea4a104b27d9ed2f3d961008aa17477e1592e04880f0938a6c713e5cc0989f889857e9b5639e9e63a2a818285be3fc4601780df258acfdbcba39ffef9322fd398250de8f6090c3efdb7fccc50a1254b6f77421437cb83e7e61fe86b8fc83a17427178e2ce6f75f3b3bedca0b84e5235bf8b1e15498395ca1a1a6196340859eace29b5e71659e2b61a1dd74fb39b0e58696e79614a966639d52529f830a1b4dbc757dae5905def878d41caefd994f3c7a3d0ae7195b4bfa53d03dcd4e90c9524b843e2227eac7c1f8ec91637946691958b425aac7928ed6c4c2d2223503d12bbcdc3ce3bec7549caa8af1c8ccdeb2d68ce809c6344f4bf2733cf2b4421cc6f6483e80df7a27802ba061fa71c6a35cef51107c1e63bc19e218acc4f866a3bca8316f43b2e45dd44e6f38921b8cba17e1829784a471610a8ca710b524e692df3e4124948d2b592c594f72d172663281143cac10055210630a9fac2394eddff4592b7483556a16fff5e12d876a39bc0675f40f2ffbbd7c96d2a7a75d45c2c4d760ffcd393c997a46a98e745c5d0f9700efef3454f935b154d8179de0b21a8ef0e73b7450dc8675a2d93eaa9db30977d7a9bc11b299d5a7fceaacabd7d2950a32ac113a4c88fc8668aa4b8bfc69ec61c2f2084865e913992ba7b68ec788892f37353dc29c99ce352b632c4e1e1e8ef54c1f5725a34a207396fdf37f863a5e80e1504a8cf814437699edf6f79b480b844d3e1363f287b7357e6bdfa8702d964b38f4ed81477344aa989b98c5e818b201a08024a77544b85799abe99994549313f1448dbc0abc0e3de7edafd81865263e1aa53e145988a36e8e1cfea0e454ecdb2f108b86ccbe189322bec3f05b8baa8f0ce6e2f029155ccd285cb093d8d27868e5f022bdb730e54985c742d0f390342dc73649534b64424d39548d7f679acc62027585bee2a7c28581f702f24d2624171269094362ffde3a8773fa275c85b06fa3db8cf7862f7cbe3b0af1e12408516b921acaecd3bccdcd2dc1c68627a1bb84631bba86cb317a886b1763c69e8d3c883d09049bfed3ad320d86e5e8a821e88e7aab1ddb383b1bb68b31a58f2a7be984075804e02a432b7301f1536493f09c1f0c1bb2e4b9b98124a51b570ca3bcc51d332266970268d8719fa6ad6564897b8cdcb12a9ec340a08798df4f9e0cbe563151451aeb86e403ef6f531405ce88ffeb3375fa47ac923b894fb7bba2a1a0689d40cb13c1a4d5859dea150dc0c8a575dd93e4502e7da6b99aa48608544cd62aeea3f2b2f815ab91e8a9d939511d8c09f12d8a7464338f300a20ac0b718be7e63145ffffc20e7cc87addebc52037f32a9dfe6c61193e937aa94e8429622df204812c96b76421a4cc95975a18b7f65adcb5b0834754b9a1ea945e79935fa5bee68e2b241be58eaef8595bda511be43e75ebdad2783544bb6ec0fb2de07ac2724f8a1beed040c774bd77ce7aa5f3bdeaebd8ca7d492731f244c0339a2bc33672e4a0f0a4afa6338abd9d5627f084c0a46dd9d535f459b5af28b3923d491c9f4baec48de85cf02994cf540605e8879b8ce36a0e78fa67050e79985e0f0f28e12c73f336f5ef9661c7d9fb2522c15081dff6c8246;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6a771c3c6891d7bd2c97d5a245aca8fe40772f8b833a1f501db9cf6d418f94f4a503ae92115bd3f74241a8f0d693bff68f1aa06ea418c1cb8c4d41380fa1e49b2461d070711b9fd11b65b23e07e51f50095bc6c6ce7edc334b296fc4b5f8a240046e49250e329bd342489a94504d3606f5401d0ae160169470ebf0210dc87d1fb9a54e3df77ab1356a1e3a710879b93ece3f88575e128c60abcb6724ffec2960422d81a847b14ff72125e27397e70c1d26b6545db5e6b41d96f8d821ce8c6e652973147cd3e1bbfe5229d060a8df6e5376057ce0c8d0a8b1bfe920665ef59f00512453a2e42a8d8b4c62582df827ce5658c6232a22b1513428db5f630b05b14c2bfcdc08a933266f6d12fdf363973376baffa4e431d6df5ac33eb6dd94554025fa8c87bb47be048fa94a02760493c93214515b5d3c41d626e7cc8a4f19508c9646d566d3ac82aa49f29d6feb34aa1bf5d2e05e52921a004f52326afe005580ff7f049b3f7dbbb9fb50793edb2f6cf3455dbeb976d7227178f95863908ad53c271b595976b1c316719d98e84948083e42c9978920900c28b10098c68a6b6f8e11c92ac9ee0b12507b449607e6e64ab3db8aff96f22ce5bd67af31d1997404bc8eae0b246c7a5cbe052347fa405ce9a70409721599c0904bdfa3bb1cb4b287a6214926a1abf4ca88411655f934d167712576fa0a92c9670fc17d0a96a568fcec5480281c8b40b663fdac20c911f924b8587d61356090e6c3059998b891c992e4d9e07c0cd32924a0b2fab88b7b2df486c2d979ccee7ad67a1ea3fcd9741990444a685f2d01cbee3bb9f02d49d2ee71a79d4e022a952a2a1b8486fd63a77fea94d726093490cb8fa166ff47a38a54fc78ad1547484269d61cc9e16db681603865455da4416d83294efbe13d9981a19fbc5d6ffc2ab436bc493d37f09ef657bdb16499c4cbdca6f30f1b3eb258106c7bc3f6bf7b96432d36bab7664944cdc8305bc80213ca8384e0532ddc822ffef88ed7dbec999268ce4ff532fe9a01d4185a1a1e73dafe004400e324996e934b61852b2f47812ffa0a3cb15362ca39a7051e0af9c8ea0dfd10cc21a35b48fbdf4d13287f6371462d0190472ff7da326083de6fad755ae89d5f4696f8a1a31f2157015910bfa90deead8198ca6b2379c2cd416612ffb7f4b1e1866c0d7e0ed9fb39fe2adc7b7c657952c19f148847e04a5eec8f660c0db2bb991a6bce980e45f1253f98eb8cf8c4600312f54c4da5f43553391077ef59db77057207bb67249537f805aee86daf8afc401c5b03e06eb5740520ba038a29436e428246394d3577b76c7c74579d166350edbc4524ffe12af4105094670b0b51b9476a4b18cf53f43f614cef48447e01bc6b0be0bc4f23885809f324c282b6c322668c341a07147e335880925fca6dc5ad8ab3601a6493b469a9d3e90dfe8e4a4e2282aa33d1805de578742f8492be1f7d4200485664b81f4ce8621337abb191036f417f23f971b6004557ce074a0d5b35b5b3b426f1541a0168d8ec364d1920e7be6a210bb31d3946022b551fcaa507baf8a29a81f4c89fc7507255ce015264bdc7640d51375afdcd41c3ee31e7ac7a7ad00fc85af604d9c7b274f91e94da536aa804e89273a782e80f2caf0765682f8f57ac6bb5aaeae4b83e84184d8ccd528612a2a37e9854411722d1d8e17d5385228b7f1512b0806002173234fb173219616f6ef73aef1f23c15890e742d6ad143a4367977cc153ba9d8587db42b47fe494f003fec0cf0e2200cde1d309a3d44b33d30c698a65ac5171a5e566bee3d7ca1657f186b782fedaaea31ed42a0c58368a2aa56ca0ae00fb22663c08fd35994607db6356b37be9d3c6cba304c62a3c38c5d109aedc3fa5878e0891007cf0dd299e6a8c82f973b8aae1bff7002821a37211d9d62ce53b75f84d4d0ea8db8a468672709e81a2bbef09961417302fee48b654ab6361ca54c8121c1fe4afcb81a0e2c4fbabe9e67e85a3adb558b6e6cfe17c418f2283b62029d3265a3392d0d4fbd7b3ddf5750593afd840eea345fb0a171c62f9be47c53160de5176082169d9fdbac9d117da6fa06e4159ac342e775240f81d8fe88be0d0b43a810391c82e8d261276990f7f6f19966f25e4dc77dd453df57fe6a88cffd6930796cebdd346d18ce61c15dc674ff7f629b596b2bd929e36e11605fa31a5c771a98a178e22f62368686c973fdff311819b84fcf01a5552d5248456cd834381e34a14512c63f28c94d472071f77194f80ee803ba5db7118d6bfd8a2f4cb1d0c7974049aac8c1b8066893dd974e7ec5abb59e1c165577b0971477e7afd731b5d11f7555c782d89c9261bbe410927871b8f5b1ceae53c78b6af4d39ef4e4cda5b39bf968ef401473517061fd924f32f314674e1da6c0078f0ed7cb4127787689e178c32811050f1238290dae0b8db5089ac12af1221a4d68a45ce7f0ba9251f2ea859effa483a7a78ddb71a1f58782acba5823aaba7d048b1793c81d6ec8234e16bb50b9d53b8707892aafdf9010ddcc6702382b3ffd9a54636dc39c670a834ea320d9173944edbb79631025a8f639cfa209783fdb852506dee0ce33268ee94fc3eae1e22347697bd98b9029618af9d4f002902db47c35ecdb87a22d9ce2ebca711bebeb098ccda15a7c6ee565ec0e9291259a2880096843baccb2dbe7f30bf5a32db03153aca746b5f46beeab1d3195007562121ed9107db3e4386a8de9f4e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h3b9fb90dfc0b847e0d1e829da1fd8872b79bc3068f29554e6766bee58e8912190b87f087925e0b98ac3c8a466841c0682f20cb88455e0c9a97fcbbc205530981898b23a93bd4d2cd518d6f8e31d6660bd06fc36fb11254af7e4f9cd179d386d3d16146246c4473e63c8b4f9d733b4261c2fa09da004d950954c4e26086b942b894c1d6dd7b0ee3e0cc809a5638dd7dbb74344a8a971730455b3b7cd070ef6223562c0e5a469e8f898d97d4fb8e77b9452f6ba8befda29f0b4535dea1c3748a9591fca1afc22fa6a9835d621a07d57c3433a7440f2e24aacc172b550ea4fe1a18f2a3bbdc0d107c32e8053b15fd3211f2b9cd92a3bd858d73160ea77ea048723568eb4dc3f4260147208df39603e3ff34d3112afcf68877b291726282f2d4a220cb62840bc689890915fbeae33f67e7101eb99524e99076903a3dd5b14617799da9d7367f2e1a1b84fb35e6b53a2cd95bca4303004f56f315e7152c694dbb4b284a4acc12607f9bd4375a33358a7b121896a27c63cdf37556baf79f0d99536a212eb30acc9b42b0e71d80f539db0a4e50b6dd3ae3098ed5ef88ca8e1f2590d66ebf662493181cd758405c76ac0b64a28d3a058b7860bed393d703a748ec3fb356505c00d9b8221091a0da2cb49e622c2cc482baf9e9714a19e638d67254ec5fa5b0725efe57095b186204382340ca18b4de57dbd4635c2fd7155a8f7f181f53efe0b5318a976370698e9ef65447321b4b0fe61673e1605b0b9c21769d5c5691d48a8907f0c36b836ddc952816c7f09d6e13960cc0117731bf199fbacc51f2207b418a3c17b3bf8f9d6147881971b8e8cf4c63f65db063b1aeb966ba0042a7c2593d123fddd8ce15f0c7b4c73c98edfbb2ecf5dfb7dee22ba6916dfa95d95130f07b2d9a7e0f0520aa947d3629c94a4d9dae0eaecf7c1e7481c9f089324bca7ff1c32c7be627ad2443a54f6f204c7da385928e8243311534695cb503d7df6d4088b7a6ca0d5576eae4edf31f2841a3279b2b328f9277bcc922348ddecefce50ff6e43774dc36f6d224cc4b7d77a8bd17c9b68f99acc59a4d40d75ba92116099d13aa359b2f7db994fa671a7daffab7e27a971365e95bc99a723e94ec5425bbdbc3972f50191fc7c63c8cb3118d32896893cd373fb999c5c90c3a9fd32fa3cb1c6bd16d276b476489adf678de235aebc9c63ac00d2b84abf3aab7b4a4642bc3a29d2bf653355345128fed93b0b72666ca677ea8a0eebbdb3bcfd8ab5d9aa70c401856cb8d7e433bd070893cd5790b989e6a03402758824faee392408f827cb6f5dcd625acd1745f576711181d6a7efae69a8963597676165260f2dcddc6a1be91e5b58279aaae09c5fa348afc680b5e0c5cef926f5e494f461a1959eb284295f0d1014c56e67938bba8bd8df9a1e8aa625432deff1800db34a7631880f441544154e4e07fa202cb2bafb3279d5ae738f5b5980994fb0ee339596afd680e850eef4ac9c7d6c57ccf7b0bf5dc068dc2ceefa18ce3a15cbf29e1bb51b6864901d3f37eb58ab35841210954dbd382b83edcc69c381ee8374ed99aba915691b3a2b62e8fe7b0610e9ed302ba91867f19773dd498ac4a22ac911de7dc716dc3b8d34b3b3abe920b9af68b285d08712b169d098fd7a93d3ed5a95bef4e274d647782c4ae8b638736ed99339197c4bb80d3f199ef526adb912bb448bdb394ef022aa3fb3b6e5d7c2230b0f222ef226639af6d5a66c9403546cbaa416ad8e5bd9a2417ddc7011bc029bdb3fa9ffc770bcb985b61e50112b0489d999f637bea79da2cd3b0e02ce571cebdcdac68e5fdb15e7cb511309f3bb7b7d645e9b8974a260dbf914ce104aa12f2edbaac9c4933cca7007db814109cdc3ec062ba1069d5a68a70214d58727b5be09cc50c0a0321333ecaf9de1abe0ed5b2f9453f57b645c8b070b656c51e965a0c4174ca5528eda1ec0aad843a35188c1d7019608631ee43bad3a5f6ac550b3b2c25eb46ab49ac62d6ee7bb946370a282ccb68011edd0d6fb2f54c87cff0efcc11cc0d1981b05e953f2d922dd0491df8b7c1f43be8bda0586b0ea10f0b6676a6725f1b612300c72751a7a80cf90b65a051177106d0c4a86cc4939e81a76dcfc2642a5715e23f9252092c4a75d963cf9875ac3cd516a44868a8f562fb2757d8fcd5c703e2b9b7c0bd91343ee1abdece16e3cccf988698d40f97a6cb486725a3975c8cf8757e8b5019d917268990d0c08873baec94259cd044a5b804fc7357c9b0559bf49efcf94144b2d35a4355711f68fc4ab39450902777f2560bb1c7d1233082e5a99a0c4fd664f3753e93768da67e4f633d05cd2504368e949f96ec24325f36bcbe8426cecc5bffbec9f35e2e53c81793b8d1e1c3d6a77be942455919e11a5c096b3d04cd6af75d3cb7f64ff21b784af7c689ac8d4fddb56c0b688f528f0730bd3e290d4a3ada03e3ad11a78c313f4ef09f162e8e3c2802631c28e6bbf6c40e38120e1254bc57dfe152b0d07b1f21ab10a365a945e3430fbf2d6e5f837daf47ed801b3a6981b09e99ddb08aefdf429f1bb1a6f883ed072c24e0375c7f1572df7989d0c022af4f12de0613a64ef9b15ec0e7fd44f284a486303c50033cad843409c9bdfd48683477622753fd082f82d547764c5d305ac5d2861230ae2e26b1a7467cdc67d0a1d320344b78c5ddc7557c66a2613137db83fa48bb19bae47f5df2a219c747e89d99d5e4eb39618f2a7c04d582fc27de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbd2f13ffdb5d1c896c6353b198d0a7319985d59fdd0705621991ab48c49e6b3434f99d963277946b7fd290cd55d273a13d096c98527c9d6cbedd7fc9d9d3349098bed697de316460a18514e28f4202c054fd0cb08d4bd86f20a54b5bf78c8a35c359648df1190203c3892473a5f1a2a0969e568cddfd566078da095e0d1b0fa8a095c2f832df8a2e11a30c0935c7a58d7afb04c63c0852a8cc8b11f554a9b9daab7e7452c078b22ba1f4906b4363a7b85ba730e4222895570596e9443f10fe45409a0e6725fbc95aa0d9fefb7bec420b2f30fd486bd7d2e860b66b8c17a67351eef089f49f571d060478d064e577c6a7b1771e405ab973773090c6321529ab95a581d17e405889e5138adf55b7d6cdd30f589cab3d6da2c554916704685fa14a10c755f061be4b900578ecb433ee61f115629ad9981f45b4d895006784b658e5b70770537b8a4264b7af3b02157870d45e211663d2ca12bc284e524a624d740d973ab39bef63c9de98d4131896281ae6451bbdd04d67f728b9163ba49261c1b6ef4003a32ebbfc603f635adc4a60ac3e965dc14280e027efaf9fc266e1abb35d778d4cedbc7ec6e139c72fc68adb4a31bb3c4589b853891da0a5615be16dd984ce43af8ef3995876a749fc0a04214579cc7aa00d51bc973f524c8aaa3fd55b6f69ef2e769162b374a89d554d673529a45eba420cb13901e7268e40fecd98f6e1bbe7832737de858aabe235cf3de276135b2d0920e696341ea8f9778ba8b9ca1efffbbcf1fc9326746397466b1491b7180f20ebfde62f5ad75c808a190dba7c6bc0b98744e3846b90e85e5af05f43157900286761c58030a2bd2c025de40db450c388a3d1a7a9e3ac80ca12fdcb3e4f5e15e96e648486f9e0b38ce2f632a4a99e814d88f26aa8e99a615806f4760f99736ce1566c3eae9b102d61b3d71ac46f53db952542c03182dad3cdad2ce9579fa5f392b14581483d84c353f85bcbb58fa79a8bfbc79a9deeb5b294c2c38493f1eb5623f4256e0b7e28ad1ca36122bb50458cae2b2483515109b0ef3a07d15e4e53ce8312f8a5aafbc5295cee2d35221f228af17fef0e614f3a590eab0972d021e73de3dcf18cd083805b857b9b9f63f53fe1324359502e7d5c37cc39e380468852e3b587b78b6fc1b8f7b0248d07f0ffcf61b7e09678d118ce31d0060f3a53733c7385aa89bf0a3ebfa208422e5f3ad05e6886261c0ad23595a624eb3ae005e7a1c1a788f4fdb3836a441cf5ef629f012926f1eb75025918fa9e05f8e24693d2384b7213f3ec0cc1987fe47cbecd5edc1ce62b5493ff62c0aec9ba9372f989bbba10a740d9fceee093ab517e7a7ece4b7e2ff8101962628194aec124584aba3924ffb67bf8145f56b0c0b71f5292ee8b69572b37667a8f024cd22a75072a9024d37d9bb15640a893a4ebcfadb9b8a0c6cb0653a08404caaef432022ed472cd290059e8f107bec59b25347e18c589f88212dc3b6fc1f88472068e4af5fe5ec5a074dea19b0b66b0155f6f83709948a7d28b3a9f7a96580cad5c0a49877871a92b40e0e0f3dcb206f65c800f20aa033598daf6f19a5ec3863922c7a8ada9a20869b9c04c066d1be1b5af22043cbaf116c6c9695fe4cc02ac38115ab29fd43f504606ec825b35cc60bb98765288e945b1025645207ea653c194b1c91c573beb5d2d7429dc9f27978a5c7def3d7680f9318f928cec1d180eed643e07eb40a0ccf1ca989fe7f23045d753554e08a8c8afaf0bcf43775b477d8d3a606c785a3f0c8e20c4d7ee0ed99114d0cf4753272a153dcc392e60867caacdd5a015246684468cfc08d2b4330f81d621792fcdb8c4d032080c56fa6ad2457cb6060d01924b2e4c8d5280006f4649dabe673a849303fed8158930bcd05a531244653de8ec40a4f868ced88478099ae4b9b8613e57194ed726ebf1741be06c6cea35d4cd0c88d6082ef297807da44f893a0384fc3a334ddf2ca21450a320d70d2214bd0edcfc9cb0de5fe58f178664b570243e7c7d9c3280c0b16bc8bc33b3d0ee670669381db08e69ef9042e5e1b814a26e34fbf142c494c6c3bd430bc002fed65b726af65db034fddaca2b537cf60171c10f7a1df09351a7799eb4fe0944bb98d3801a170d8e5237c228ecd314c815d14f474f81ea79bc88405c12aab6c500460c1166c12e90ff740b54ca9696906851a6541248ca44bc831535bc8978225cf96420c477ba5eff8ec50f100b3fe27f018b203513cc6806c97e942a8d63c602d09b8e78330bd078b7e0ce109dcf45e3844cfb16feb49a4c27dfde8f1eecf0b9ae9ffbbc87c74cec5d1184bd7043a14c329fcc877fe00236d5a6f03730cbe0689cf8a3ceb675af5929a7de847cab982e829ceb4ba6f59e8016ede9b0c4a168a1a3b86fd9479ddc2c8f61c0a39c1c29b85c71e02b55a59cc392ea04ea6d93f599f358a908ae9123c8fa115228cefb404f8ab3930327722331b376cb64f37942eb4fc06ffe7ec02974a0e7f19198fc7d361f871d5b41c49d9f9ee4c7a099159c3278c4fb96d3fb1fe8c1fc743db4f451ff8e3a0af3952bc1a9d0de0f4828c532b5f16f9e55faae1471947c9bf0e6a940e65eebf308ba52bead25fa05251403ef56ed75c64889c3fdac855ec69b560002a3cf1bde08587c9497a5df591161858e0fe53b0e7b139a493181d342558723c42233190eff87834613545e6d3020824ad56fa4dbb62401ff8b355890a3b8a4b826714a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hee430b803241ef57f49d36ae86072176ae8de019536c6278d9ab643e20ddc30539fcdba19db8f52fec13667665607fbbfb9d5496f6f9e3c983490fc76d56e6646ad11b0c6720e89e9c068be098222f9a2e0f647b53965048eb5d2decd9da51cbecec5a3d358a63b9a06863336e8da2eec114546174d89543c55c6b54f78d052f03f185ddd6518ee5b1b3133f3e049d403d1b154f2179f74031ce2e4bf546fce79a6d0393568e943b765420f1df4a93d662b99a18db1e5227d5672da9c218a2c001a3d44058a2d053233de4b5687daec35324abbc1b9620de7bf8f4cbeff2f79f0d03c802530ff557cfa6ac9ab89a897de979ed9336672262cd58f742181b1b4967b7879f249aa52aff27c34862ddb5797420ee97e3045e2fd27a5b4eed4f6c098aecc9da7d935c1cfe12650ea85885f1a6294f9902f48badc0a5eb02dca77b84c835f33b897f387588032426a5ca29d32bf76d215b427f128484b37ae25ef6c2435e0aeef80306a7024de41408d3af4877f57927d84a5f9688b47e65bc02eebe1836bc070fda26dedd387d73e84e8f51d7e526f74df018b953a26a376595a18fef963f62cb41a497fd5ad958119b52462a36e499e5cfc5a889ae4b2f317a95eeb559e5c5c214c21d77c6f55151b7d095110727357fc30d29d8f0d53f2159671c8df8f756089686cbaa930e6c940e919d52208184e4c3abcbffba4d481bc4d578b6ce1cee7926d368bb3bfd60a052147f245dbcff48f060a3dc8e883e24163fab4ee9ecee8faa4f1bb1511feecd49b383d452729f644192fad6203d071b9f6ef9aa2760d835d8bc96a44c2d61d1592ea2da1bd9e5497cd4ecb440085f34053d758decd6dbd1ca09ddecf3a892905238a7efc904b54df1b9224c8584d222f7c5e779fc819024da2a57d347ed8c24ce3b7c024ab2a1bf393719834b61f693bec067267a6b7691395bfb07109fc503c6a0bef0429f8e011d15c7b9ccbdf238ae8433798da2b004b6e7b6ff4d8ca6c93145b7bff2ceb337cece0b6b27388ab3fe943642d6b10f38bf0673787514926e81df7e9d81ad59ec98eddb512c29bd54e8c2b1dd6e1bac03fdee8a75c16215204d393ff8689db2dd98d3f8d5f0311a6d9b82ebcf75ce2df228ad886d3513bcf2041b41e01604ef378058c88cc4e4a3ab4b82a87d6850264a149d014eb16a88b8e4a3acd465e9a8455f7b146638f34e9ff08537bac6b3c6b0c4bf9ff32030ee56c904024397c9285997d0b833430efe91807f1e4b1ea3070e5386c7f2a27e6778e039b9f8867318e11234a2f13a955e3ffbd6efa6f939e2307716f30a30a987774ee8799c2d2821ac27e7506e866978edfcc835cb4f94382285715013aea36ab6c4de9fc02688f95ff9beae19432820cce141b25f3f065d177e5b16a050e85fc3f30954765a0f9eb522a74caf5b64246c6c3ac91e705f015efadd1feaa0fa749d9cfbabeddc1b4536ff69cb9b1eed0ce3ea66a3ac93586bcb4f97320d11399171d99c7c6a6801b61d1a8a1b8266881de188b2291d89a4e0b34c9ee8be03503062e00f263c8a7c10ff8188dd8292205be84629b5d96babee3b5811bea7834588831ec85673f2274999db1704f11ebfa3d9e8f1f12ffcd05e451477430386d03aae50ce864aaaa6557d0160a8d41944f5834e708036b312c0462d5d4fc274ecab73a3483b9f9910b0159fcf9d6c2b8fbbe3868af9c3b7716ff0710b352be395499a561102e14d651362c8558f397fec7552639da43f51c88bee2aa585e04bf7bfe1ec1599e3d9b33a7e330a9582569fc4fae472aaa21cc762946fa1433fda0ab80c549d8640556d05e707b43531ee6ca4a0e975e3632dc79495c3619a6f43c61acc072d11dea6e6b9fbe9b8fe1d7f2ea732c7e2a0947697a5f03ec673087a4343d3bffc000fdbb8813d6bedb6ec29922fd8fb46bc923a7628bdfafc3d85227d8a50bad052b3e7d45f10242b97fc3152596728712f5fb809ff565f8258c743bbc909811c780bf15f8e6666dc0979a35d7ca6aec3ecf28d026e65207018194c9829062a30c061599f5b8fca1059da3b89eeadf078b971898f606ca4119aa1353a5529955b4bc945ef1e804d641dd930006fa615912dd169e2c780b836a414d10770093e82cd0adf537aeba3362ccc4825a848727e9c76cda9ebeab1918015f11a672def9fa267d116abcc2098a32a16e18787c3c979522a890233a10c4f7b628147cf4c065c475ee1122f2b93f454ebabf6efa157d4bdb91d63b495d72685a1cdacfdcfaa19b59f0909aa0a0ac4a2176347b649a30ab9a74d243420e6570a7619e00739db7206619018fab6ba2384360c897e8c9e205be04e25b90dcaee1a7ea833173f5f9483065d1a4ee16b1dd9f9031111e49c7c43337e0c497480b1148d93712e10e4242a4a4ec3ce642e2cf4fb6494c8b02362e090efc6fad107b02db8648af635f07e5a7c9955c6141adb52b78b59034c5162827165acff42a0c2378ee39901ecb9cea73db1c879c2ef52f49b45647fb74289d285003e9ce265ed63baeb5c1e5e9d70cae5c66ebbe95af056656041bf35b4b4880f9cb90473d868e32ddb6c279ad0366fc85de553717bcb565ae9b084cfebc6e76196d359acf902e7aa47e0494d22d16faca0341116139e2772b4e29e15dbfd7ca588725fb941a525c2a649efef12db03fda4f215a6b053dfc51945d7c9ee5081c2b1063d36fc65d5acecff63fa8261c85bfa6623ff05a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h5c2f969f57882eaaa094a662ede59e3f78a189c807c8bf5c9b2cde11c7fed49bf54d2389e1c3d84b9ec6c2777763cd9bcf542d00428018f21bcb6dedb6c9895655ee398198c5b29dc862c58943607a399824949045c04b76d3c3fc8619f0416d5f5e5d1103866ecb3310d33bc73ab6c8f8408a2dfa295ef2cd1e87108eec16d93798941a39d6a5dd5b168e9475f64c3cc4ab6bc58cfeba03d03d43a4f9163f36ca5aa138eb75133940ef672312166bab3ed55e34483b702cd45a9fa69b0fe045237209ee20bee5300d6cc004203cd18a1adae679249929ce1fe0db3870dd5e5f65d3ec9f8f48e283eebdf3ddeb75965c5fff2f6dfc395ecc165d336ebca7f24c60ac688607249a8187679443711e84a1d0e4d92a3154b2f0923c015a0172a42b0c3ed777b78fcc05088036055be59aed6d63ec95a3f8c131e14712d893e61611f3e25916ae7d32237260e561f96d4f11e16dc693005dd6c38132baca907eab4cc49e545eba6669504d9cad98fe77e8cb41f34c071fda1c15344d569357533452d6be786f3b49f7d5b190b22f5e9e8ee06fe6545188c061cf090f46752ff3728c9b61d7bf79091db4ffa3303d1ac8aa79b876d6f71442898fd7d87b72297da624312ea576c5f73c29f40861d02295400d17c989060ac93457abb57c8b5b1fe93f0e6bac4e9622aa99ae7eb53950f8244d2e8fc988c11f589706168de609d772ce08df3733e07377e86fe31fe529c658e1eae1e762a4685e7c936f4c3b9dbd0d0e940e5edf716aed03eb55bef5b7e0a4c7ffc19f194e5e232d3d983716576e5d9c69e4213906176763a7248d2fa858c97b108842dc71c1034e161b67d77dd543a292b9cca9091d52b6655a325eca1dab8cce8b08c86986146810e35b47413d70152d76bb177074caf6f04fe4b04c5849d04285aae71d5b0b451b1ddf6f094bd6543effbd8605bc817f91568d647cb93f7035280fa9cc752eb54f2e707ef1fd749a039f4fc6bf8c2581035906bc7948f1b78a956ff09ad0b91c09251ec3e9f6b9ae011bd6dfc556589f5879d64e7bc4b7c1cb11c21302468f9eefd73fe2594c77074f19f5c90cec60a68bec60f0a1b5ef8638167b3c619f3052b7a7568e475853fe5916055543f94d9d7021f7c1c8ebebfac95a60ce88494bb0b60fd0d04e8393c3326b576e937e1d31d697adf40fd35bef535afcf8ab5a511ab330bb93c95f1d39b45c890047afb61220e7e004a62c461f984bf4802cc4b1a75069c30a6438949b6ea972f8bc9179d924706618d8641d272d7ccf6693485fc83dd2ab5399e707d5a52dffd95ec83fa6ed79bafcfed0b0069d37e786ad33057a6867af6917b394480ffdb17d30b204546bc63b2fec10052e5ac3d50b9fc2703608a76a51a404a0b2b157b6fc0ac55dfea775dce148eb4ecbe17b3f844d838038c18c9f82e599f882044d2d8996bdad23f7248fa675058dc9a6eaa5c11fa4f0f8e0e4089fd7575b75c7df97421744aeb39a70b3aada45badfa7fa77970e7cd07dd1f2bc6fc4cd61d56950658a1a8ed8bbc37aba7c6ec526decbf19b84f43d7ad722aed38814240c9a1bc850244701ae7b1166b87dcd8bcd32b60ef3e14fc1c839fbcd96ad0adb03f0652ffa0fd87bce1d407695b78f8f04ff9a58b5df134cfc3887b30fa3b11de7a11b8cdad2271a2b5a06316d461895a8e32296cf81ac543feb659096fa91473184f902872711516bbda3c18ef46ee19864524e2d7872243faa3235991f91aab24da603097ab5cdea2bd87e1c3a2e1e935747bbe04eb934a01590b075b3483604aaf4a8193a1be998bb959f596064581cb1d41eadbe18faad309ff9acec3a255b7dc17da1cc7af877a487e2a4e4c499debd30e23a3f0dfc1f2ad74c7c460efb9b2cca903e93cafff703146530a7d3d2a4c917fa378ee948366591414d6587fb7147af6c8c75b961760e085d9986156c8381accdc9322ab4142c533d7bdabdb2249767620b7bdedc5bb8083bbc9097c00ddadecb27bf46d348cabcdd686baddeb23b4252541ca450e1ffe70b66465e050855f0b8b8aa1bfa510627e5ee891950d3a420345b20a53c0c8002f428285a595b4525b9383cd8e0e9a35bd650d986de37d3337f0291ad92a48e18eeaca0775dd04036c66fc328455db40dd6793eba1b5253b724e4341a9bbde04f566f66a43b9abb994167d9130abffafd7ddb30ab0c5eaed852e3fa798c01d330248503c45b9627c49442e163213261e2e093a4ad9cd724a189ab5d25f646142863cb63f752e49acc6257bdc3e79805575b410b2bf52607fec29b9d0627e3a268554e460a992fc4295260fbc2c2768ebda8cdd343251a960d5237a11d42f3a1b30eb73b85e85d1a1de5fe11bc10262339a797c362f9410f30dd3349e0317ede2a024ea9d9b9502290cecc271991b8439270d5a285df06dd837581092d204bc9be1e372543009eae616b38d5dbecb04bfc3318296cfdf38bdc3f3e8cfa2f6a3e0167d74c9896a97abedec720ef67e7e1987517ccb6ed0d10ec7387421a253513e584f0173c5b3d2b4780f2fcf1b800d7feb15cb76ee17d4745d2ee3209f2f4a28fb1afabbd8970f18663d55cf9ef32d51a436835686990ff51d34c8c32385f669dab429a8ec3aa751b01f03443307479c1c0bbd2198ae936f7a8dd4eefff745a2700437a2282896ceb292c5ae34cf3ebee076c15d6531568ab4e71d712ea4b13faea0b5addca352cdd04365eae5a93f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h616aaeb6032aaaa2d18fea7d4f60dd2b4866eddc7ada2af03a55bcf17c4e7a265fc9c779208472298f09e649ef352af9b586b4ee6ece8abe07233a06171bc13944fe599c884b54ea5fb5c104ca57a3327f96c18645c83d860b0d2f0663d5c530c1b8bb01851e25997839b561a5f81acfebd04697ccf8fb5d564dd52824dea0eb4be52711cecce8da2e7067829abee0344e6789b87b97f1976d6e0352811defdf48232f254c3911c4dc6f61651d05a34af74013853832d0f33c9411d9f19c257946e01bd2406d53776c8c686aa90f9e1293827f4728e8d794d25259123d0764f0b007a5b653536aa0e1bc896feb05be03d1f838a8c04e18fe6e42e04aed2ffafafa12467702571cb02e63853de5fbd98f221ed874a22c4fe84dd277cba4957d1a3fd3e049e58eef54318cfbbe0fccc22143fdef29d2baf7f03dba0861bbe03c8509a28555bede329672d52522a3ca716fb6259215f9b9d0ef2965f227ffb9fe48db36d1f980a1bb9557296d65ae78b9c6a8e44e3ce40c9b74f0751ad6e9d6ec6da95171d8b0469256a19c4faba73de53cf301173a701277d35217214dbf300af02ae8e2dbc31faf08ef978a3c5f358ecf87391911ae74b98594bb6dc3e630f8fef44767c92243f403667157e7b92c256d2f40c2a0fb352587fb1904ed36573428f5f22a03dfab3582f9e407e4285442254662705ae94bd1ca1a8481126d8d7ba5f2e42eea4dbfe242c4061e5f3f888a9fc578590bd7b22ab59fc9b4767ae50485bb04045d055160186e93a50ebd4b83db88a1c2bb7c16a98ccc7a9cf72e73ee0483aceeaaced5a75abfb81dd84892812f31e089718dba51b7f0d2c4a7b5219c4576c093151b1c54e81276277b3b8de79b6980d03774034e49cdec2c3720659068ad18010f516f7b41c9edae4e010e08848ed0123a147cd8047e833a47f5be27d05c34f659b55e6958ac27fa1e8f9d2f559c4548fd672a32385ae309c4e02db865418bbb1bd2c1e044d81a13da814e4c6721559ef186c339b7a0e46acacbd79d4873406a935fdf7f9f98696e431b63d3218e599fa3db79f55989f68045e38cb1e0fd43187871798bb2950f908ffa13bd0dca373d31dacbe0ad546c013ac0deeaa4f3e20dca2bba7348bb3ea26aa1bed71f681593b54d89f2f3d11fc1c3b14208e12f62f8e1873c6bb977599135f9ee4f6123c93560578cf9f5c616e80159c180ef00368d1e467f5596ac22902948bf62c4abb72f759948ea0f41744c3ec77cc30794081154e613ebb8d301ed7019ff1daa41b86000cf6e2d030fd7f7b4ca5d886f11d919d6dfc4c038f7361be6321303f9193b3003e316715ba2971cb695d32f66112df56e5604cc4f28a7ddf041c26799a3b63c54ed82efbee330fb80c2d18390e4a2c25771fa14da7b5fef23227117b13343fdc5fde819929d14d66886545946a6610e30926c2de6a5c3e5e3647c410fc96dabcf3ce7dd154d3c75dfd3e2cccb8eaac15907b95b3de029a6d0dea1bbac377ad2135597ca046df7e0e95727688fc2f72c0d8996fe43c3a86bd0fd22bf976cc80bdbe334e7e11e47e55476d92440b303c881479e7f485ac2eae7503efbe1cca3a23b5c7553d485477a8cfbc3d78bea2ac88d5d2d0281657844a8daef94cef3252d32b808ef7106430858b181caa2a174f6e065d602386844c0477c5adb25d94ef2d092c7f47be6f33cd802c56186aa817b1296fab7460009309800fc0688880e4ad3595b3956d67599db5a9de3467aa77766f3373d66235f276edf8c52f160d1c9c69ce3f7b61c45874f329216a6b0662325f64c6b5c0ba37980ab3738363698cc13c7aa1520c60a6afc05f23b193705bcf32fba66c488c946937c20752b84470e56ed3cf583ac02a1bbaea07b68baba01b349846efe09b06fa01f8a1bb53a400f2ae962305b55c9ebbe3527212830fe2e5d133f8cc10ea53283906c29aace4459232ef9f3ec7373cfdce92077fa2bac3534d323494a8a393141932adde98f600e4b5d00c88b3ebf5d6cefd84ff986841fced904fac54f882222d5ee01c717a9412803d47c2fc5fb589da0c48265a9e3bdf7c6ed785b8d5f07a1904d013842cdd7ce2efbcf439a25baea6d452a56c5cda688c8398cd096e6d1315ec7534791d6a59f858dd12982f2a810c4ca7eda2312a07752e056861cb4eef14322d2262c2543801aad33862571da7f65dded098349f80aaac17b2a02a60b9e63f30b6c2d616ab78dcfbe3ee9002eb5e9201590fb9b0a1adc3238a57e2031ea8acbf87e04697461273750e1764ce959de53d82da07519be79fadff696c77187ea4573f7072467e2396aed5096859fe6dd7a70b6b1c96244e3e056ee0937fea7309ed3568d17200f4c036149f370bbf79e1a650147d639a02cf5b879783fcf3c5747fa8d3a3471dc7ec29c4d968d7db8539d55d07a52fbfdc7ce66695390c4fddef98f680f1ba6860499bde05e20bcbb01cc74c1dfe4ddda2f1c074870d319f4f39fbc128a5e260c0e5ec943d8ef9efe359c9ed82fabb2e32dd89078b0aa89b840a026bd7a7653f0b37623d41a2ab81cd63a23378b968ce9dc69b59d3e78b038c29484782569f1c2f774c14dfb820693c94dd76c73434b79e3c601226304544dd19d1bf40c7233a27b9914b16bffe9212899e360dfbb6aeccb292f5be8cb5596b8572646b640a8053485b9ab8248bffd2e74bb9a11df4ca05baebf397434d5528d33b769cedfe8264919021f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hc7d66193502e6d2597539c11ddac0b903b38ad57eb12887dfa34f5d517e425dd352b7bc9ccdc5600ea55c03c11d3c97316d37e4be49ff3a77383dbfb536d1616e390ea3388e2e905534cf63f677bcf9adc343a0f86dc7017ebed74282355a5c3fb2cdb26c2fe178354c28b0828af574769392d21f9c013b2f79c839248467d44818b230fa65aa0c39f80bf25ee9a585b4a58a4369ee2c333cb084ee744e7a0129d4ce2b50bdcc37b5f34efbd2a5fbee3693952b41866e24412227db1b96efdd937823fcd8dc6097a3b34d95c5a3e4f70f9c6d231815f21e5ddafa14199e8e90bb882eec07c56f7a9ce8115fc7a781f207ca0e6c48ebb65212a1abd5ed790cdc69568af7898cf0d60513c9c8a2c8619033eb679fcda3e12d2d10ddaf7c18f7a3e6fbcfd094a5040eb69c029e872b5dace44828cf2a5612957c7c83001ff7fc805353beb23dc036cea9af9d521a4df3fe91a74855616f964fa98003411b9f6ed97493b685ef894d933cf637ff9d5262628a2398ae731996dda56efe2fc3a1d22720929bf4cab5aa1cdd0a8499221e25cda98ab26ab82f487dcd1297080645cfb67c38a26067656da90e9dae3065978db11951b92e266fe57873236e0b4e9357302c734466fcdc99e974c79a4496ca1f21e1e85ba351df1223fac8c21541b4c87ebbf0e23aa4679f39550990437d00cb20e741fa96bdec8c403f6a42996592704cde4fc2d1d247e75328e8c2c33c8dca66a7f179562b06abb635f518434ba4fc5626a442728f4ddacb632f63671505ca6a406a484940879f5cc666abdfd7ade842fc62d7d636bf3965bdca35a3e7790b1141849153a7cc10b062fc0f3f274e5486e58f7513bdca6cf2aa0e1f293f20270f39327ad8215fdcda8b32ec7b1f584c3fb88682d667f1ace467abb22b7514514f4f3b1c793ddbf21cc08c362c4da06642e8b7b6311c86756b56bc2e3290047057084809df9bd4338d4dd9e459914543eb06a17c29c18d11002fe20d3e7714bc34e15e8a4732e6f8fcb052f845a5fddf36ac9ec44f34f69d37fce7e0b9b64fb58e834dc0543fa85c4c5d44854a1dc672a62532d457024290b0535794f841760bed420b68eb80048b74fb6c9adeae76daec9591535b055940158f2d71e05137544e910ce78149be9ea9d6337fe3c365665539e43af72d66f657c0730c1d0564104335c4dcf041b6151a4020ec4a45c79aebf12967d0bba4c1a19da0dd8be84c3101ca01b4e23c37e2bf072451e73874de2c5e7ef6511600adbf7396d6fc2856341700d084e8378c850228983c89f75344a5d8b99cb5bfc8bfbcebf59993e6edf3a54dd685493f9c4d0432cf53a36bb1b77fd61feffd3d2348b1f5c5379561bfb9a3b2dba15cdf986b4fe371ca6763393510dbdc2727db0103c71d3c6bcd6ebb2fa658397f4d49e9c8f8cc854af9345285f62ea07c847fe344acbd9e98cf918a420ee3e34851f42e9d07dbb2ae7ee89ce8f6c9e81aa52dcf699a6bc9847ba1f3f6bd5bcb939d8381b44d1a467a6773c82a58836439147e1b3a9a5f10a755e48622bd4e3bbbed1c599a3d2168c3fa99d42ed03242d7df3bb6f30a44e54f8a50334cef06ff341b6ce006b7372f99c846c0c0831e433b14cd334a145252998e12cc2004226f177bca6b73b33b278c84d7aa2c021d0eea4eeae9c8b986b159bc953a9e7d0a90e95ce5b26fbe01e0168a7c08f82f1ac478ddc42481ca32845e60d13dec0d379b4c7c3255acf194678a7f54784a1afacedcc588a6ff3320c4c8d95057a74e55c28140241e5dc80b776e61615bc86b127078658d2ac098c20b210ec5c6899854c3f66f99b7cb5fb1074aa41af3054625490f30ab7290280fd735ca58aa270d73617d7e7d51d539bf2b6471f166cb423276dcd453a9fd2384ae31e2c8782563d0a185778c05302b97315c66cab810abee63d37b8a0b8e6c6c8189b97c70ec67e8ecf6d0f11aef6f3e024960c4c29dbe57a9dd849e389eedcc1afa77fa57550c65243045d24cefd4edc30b11a5c39a30fa20b280bebbae48d5998c7fd7716576dde7a14c55deb99e27508fa5ec177701d7247189c4647809dda5a983cf19367a5bb5049ad4ab2e118ba448c16607b723670546f4e54d41599d37d3cbc0b9cc86bf4d7ea1a15a559f048c8b23b14d15842cd0232a7262ac35dd39bdcd48fc54e9388f55a1282e6640b298c441f725150238a14ecc3bbac40e4b629a27ec2c0606f8e8e3273ca25a2d4f9cbe0c10029bcbbae6ceb9f66cfacee1e029e954c20fb7f57aacbc9002137fb23d9a1e35fcc228373df51602fff8e08bbc112a52050340216a12ae305aa09936f84cf8a4985378fb03721c5b50de9863592e124a7c3ec5271b9b53d57ba386d763abb5328d1bf8b79ddff4c8a993e2a80827a1b6cd74a0e86bedb54922c41dd136f7f04a89a3a5cc01d0ce8a347d50f6e57dd23ed636f42a68c698aac2a3b03fc59642d5d9e03e0cb6b8d0fa790910a8987d1994eb0f5647837f4c6e2780e84b6b408d08cc5171dfd33ce0f64eaa27979e8c6ab21f672600c8b8795540ec93323295fbcf62337e192d3b5001a8c006df3712be6823e967c9940eb057a030793dea9ec1c522be9bd4bb3d6a9299dcd9d72e8bcc251cbb1aaa4777c6089a0166e297d0961cb811436eb3858f40e611036d7cbe2a64f12c31926aae0097a9b976fff7d72e82e28aef6c74cbf67fe8c23748d2c5f95cb3acd2d5e38ae857865ccc1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he5c17bfc82b13a3d76c61f60db4bbb7d8bea641497cbc2296845969d76eb77617a6bb68e04f98d40826341e79a224be95869c07802144f44c2c5e5e879fd4d9ec644531fb95e971d0b41d923112f6004176caeba856970029481419dfd6a72d4cabe3cb7f6d1ac6665ae8f441c7f387adfcbf44380b81760f2f180074606e0db9541085fbb204c5986e1581d85db81da92f880712db8f67e7e7dd37eb68b9ba2c43e909c2da669e993dbc90fa6031d24c4625f2a2bc79164bf86dc924c87885ea2dc2ab545a8188351ba0f24cce183030b36f38d6a73d0017d8414b3b573f7d24f9ed0bdcd5c035deb8e0b7a0bc1c6602acb53824caa96f6506897fbdb56d33d054666e3afdd6e796ac64997d7f03d454b20a712bdaac18ef016699098b9447a3371ef8beac446b0726345178e16dab983af839e7739fc69f18c23530bc4bfedc10120b8218a3066ab081053fb9b571f88d9728da7d329820a1542ee660986c26c895ae8329a3f67226576b154f6a8071cda18152a2675b759928ab355f7df799607f6cd452353f69cac0745b73f3829df6f024f09cd0990b201baacac819cbc0088f64582462ac02b3ae49331d2f998843746147bd92b7fdc371b8433e345155396049e99a1c96e60d4baa8c9debffe7c1e1576c76e71d6f1a969c695e8c6d9c9731e64421e3df1f91cd9bc8e543c19af463b0fd82b28f4628fbe026b8e701b9ea39f86bfaf1f8acbadbdc56ddc5ed1d9773c81c201bdae0bf099af4565ed5de525d8dccb0d954575b182c911979a05274ad39ac8d433fe79af6bab779b212562b15527a28fc6844fe7956f133d4664d92d5eaf2881b0e2d519a5a63b81c15f905577fccf9a49ba244052da3659b0198dacf8923bfd03a8f0504fca3e73c6630954a8ab70f2def868671ebfbfa416a853cdbcb76ed5eb6a5c543dc92e388742845a2aabcab057f2aabd7a5ee129209b34f7a76ca950d071c4e439b3ee6ded7adb65966ad3b5dfc67b4ca3f455d7f7e6a8d79b138f9368ca475e2844b59113e8f56bd86aba7613feaa3d32c81b99325a4b07b970f80810895e5a537d562391d4d866c6add5e8b6524b031163a02887338b5db8143e303446b4d94462514b541374d3d776fbdc75d153adb14a0b5ba1df494a6e9200fd4a20ea41c442284194cf03102b74ff189ae26c812968503892e58b329c5d65ec65a08d3eb18327782c544936ea2c22b9210bcade2a746b7a609260f00c0a9251d0341e802ce02bac6ba1133c70cd5c73a4340a9d1308ffcd2fe363405f885291ef5a40be1d50d61289fd61bb70dc4f89f49db685fb7f145f337776c35e5ded727c61b0fc2b26dddaf5c9d0ae29385a57bf4d2aca8638f579689a49eff7f04b6b2cbcb5e853cc330513c553c8b401007798d40ee615faf4856987174b4989d66519fa4d6b7064d07c77d1b9879abea635184cabfcfb3291922d0541bae9a9839e71eebe6075c4fa29052095a032baaec036e7108ae6b0e49b50f98d1412177ea8bda43c11912ef1a6629f5fcb8f066232987e05e3b8405e020ec6889a1794ae0e2dcbc67954ce8b57caafb995d583d74b97501e09fa38c67416daa28e6d27e8569e617a5ac680ad1d347d7fb3b4de6cbf99ab6513a6ecdce19c307d95a8fc5a19f8f861c0689a331b7b8683aac4b40411bba9a9e69887891de8a8e09520de26c63530bbc9c29691799ba96b0bd8925ff596574efa3a3221a94dc530dc0ef65921f6873eec629dfaca2112cb2083a0b84fd789fe45d1933a030cf62802057bb87871f32340d8b70ffbbf34935c78e1e71b98e7de7992120343bf4b48705e9dc418f21c5f271f577c749e64f9514e2eda2b58e3c5ca46b38cfecf8ed70a04da40c159cc31a426a73b9fbb26ae428bdfc328d0923c07651111638eacf12b337f655b0351f99fd3ea10ee1d5b41522c8c0947adf799f13f82c52600dbce5d75c29ca21d52d76728f6260278975d992d72343e5375280186fea8bd28789e12446819c698114102322265c9701c2d64e395e2283dee81b6a13db3cb16cc00543f3783340bafe98a1cadebfddb21809a10fe013cbd434843aa734e140d3b58709f8d84f39e3283882817e00eed423e6050aa8596a85168c39096917176dc2a878f704194cbba9dfec3c991c6408846c4656003afc0d53b2f7d79d0391693d35e5e857dcc9a532b0c869f045e629cb8e4c032a817de8a673cada3a86f36c902159acab1a88f9517e8a370ad6e845d7414b5c7f4a856558bcebdb5687b31dc5a8d885581ae2ec6d00975c5a1cbd8d07277ad8f213f04f9fd85e0cbebf9890b7973546c25de2d5071e26a4b726aa5193c00f450454f1796edd0e97fed57b17616a994ee7a9925f080234e877233a6b7ea04526ca76411d4b2695807f72030451bd373148bfcf15d6927d7ee5fb4e91bd3ea3bbaec46f59e7ecc04c3f659bcfd274ef383cf14c44c1f22b7bd6565f8df5920e296b11fc8c977a0109c06aef674c200ffba4da4852040be926e78ef46624093a3fa72fd7174731f52845591e162b244c84845052ce383e43dbd79a93c5f866dec60470f2a3285a6f8794809d9f6209cb397a9e5563b79b300e50e670f88d831b0a21a008453617d67f488c8724cb60cad0d61b1fd5eb3b43d6f936d43077e185ea58ab42c5f563af9b10fa0fa28602a2521c24a0b01d53d8fd824e505fc06fa2304bc25a340782bf65fde6120ad20a82f2c4fff78c8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hdc23a9cff9eb466379dc4dd5feb13400523547bc84337a9fb0f81806209d730d85bc403ab9acd521d219bf387d2e9ed9847cf144e06093f5ef400bebe924e15af9817840672fca9b86b12bb2d376f1db6a0920c1482129f73abeb7ef08236014c5387d3e395ad209854083733ed7725a5d5622158e5ce16dbfe562a7e37b0e56a5f8b6573db5d629b14a8ec4e74705a44145bfdcc6ae92bfc6476fb9c3f0842a05da52551dcac0c85250a1af4bbea273c31ac92ce9a49c1589359e5e19b6ea27780d77c0681d62a96b2525b35712bbf9e64a0d0d9a34b3c1deb2ce63c1bdca399412054808884945452454e8adf9e543e6742a84ba0f78288df51d962c4a4d8e84b1b71835bd8e835948ef02902b9631a7d6108b7f21b92114b98019a17a6fa8cc6144b5028ad38b5174c47d153403324f783878b2a8f293a38718d5af022405d934c76ddbddc27a3a50b5f1f5ecae3e19252985f115667334a2b1793d4ff345d5042ecd9731112e608b1f6e420a27f8a7b4268b1da4641b2e94e1f7b5253115ab6ecf1047281c9614e5e5b05d124856828d72e41dc2c3ea868cfd22f87d2549e59ed18c309b2e5a4b48634664c32655933d7c51800298de9719380ac1686f7eba2906865477af94b3ea761660f279f598369f7243af0635c304ef85b1f8fd18772aabffb6a6f6c0924df6afc6ef0260bbca8f583e512d64912beef89fd39982b95c5bffeca2135a4386363adae5eeeac294d2eba67913d68500cd6b17a0d33509fa71ee631f82504ea3db61cc6f10438a6108cf87f18856bbc160ee1df1ec23bbad703dc2ad91c19363ea2a197255a9d82806bec6622a4d017b6ac4edad5a6c941abdcb3127a652b3fcd4279375c101df599a69feaff42017f7939d5f62366710927a23d2012a3d5306570d626c0e1e8f8038c1375118ce59e5c114d8163d1e52ae857ae6193728cfc36425ed6346abd4818a36eb2de1a80777508d23906bcb8b7a7889989ccaf1f9e8e449c76ee54703b4b40222199ac3d10d595cf6e0fbab682bf3d8355b91a157b126d3c102515f988df03d9cfaedea8b930e1725d547c68b5040fe63decf5afeb999d909c6eca1f3adc69c1f78b7d2baa0875c2cb6a5e9b377fb9fb31be29087a5a9869877d4b24f88fed62bfd0c510c2df2a7ee83d9752b00e7685c70e85e79262955b8872373ba6836229de074a135c82f5b2f991ecec4767eef014b0b01b8bf62d0f81f19919ec6c4f8848229a59e33526accf49830f5f0a90f73319c3a27fcd9d341a43b24ddab2879c890325d004709c409222c5d36aed35453103f55742d3dc96a014899b4000899f63f50fab4c805356cc14619e3727ed061430d52aa2c8ece330c6e1e6cea350d546c972964194307ff5ee161131f191af3fbc9d1abcdf1d0fa5acf5059a29a55728a1552c71720ca2293f8c617fcffe3a86f92626a7c5b718172f7ebabb094872d281de432627d8c731f876be5b21b635bd0b950154197ff1fbb5d1dcb7a68312f1a5ce7441e815b540fa8b3e629a6a8c47cd5055d4d455fd29336b67b63d54e76689f037d7cd37541d0683a86c57631d2f8228de109153ae7ac4cfdedc3acca1645892113d3f1156f90d55c576d2e153686d2e08e6ff56773227f5d2c00e4ff0d9660a5ee3e38702846e846008ff34cce40a807f915a31c34df03429527edf260344109a46074d269f0bf9b5320e05c031e9ddc93ce59736905af11493dee1917dda23304c2be53c587cc7fe03db069247f25a7dac1aa8385c2007dbe3f5fb057acd3b054777b26079fac6456abf6a7a11cb96a5c9a69065055690769164c2f7d7df470fa2a37e1fcc240888af6a8f96aeea1f63bdaac76ef1fb965c4b166f52660cb806256fc1273852333f67403f06e15c1db807664f2ef1e8a3b9fce415e6b417bdda1461f02a1cad6a984584c7034fbfb2c63a799e8bf2c5651129c176e01353e9e21b44746045b58d6b189931fc60cc31f1cbd4c0cf167e3d1bc02a9503d98a93d76c0f185e552973392444e5ee5f5c78aa59ced41511743e6f0450f36b6f475e8b63a86bc084f8b541e7ebd1106767c6219ac0589032cda6ee3d0685fb02970a5cb1103525459b3299d7ba6f8bfa12cf9e0f24f6f38badab3aa7eb58fb9e76175852f5113599f2454bb4bdaaf36779b08b677e78244b20884b295334701282779512e2b305a334859aa9021bec5320913b1eda55b3f9f6b1e2fb3ad17f89ac97cd8c6a0d57958652946e42b7df45a135543d8c1404fca4911c1e291aa8ab80f1c16aa4d8d7f6bd048041ee5f488c41edd8f50de6be1daf23fd0f1c552979ca51e286df0092d87fb7f8f82cc3977f790c163d36abb0a3b11509a417e4912731c02552f8183f7ac9b1079a0a2d3730991d180f1045831a7bacc47bbbb94fdafd34527ced66fd48232cef61442a165ee8a185c7ea17ab1883eef4c97877d21361b67d977920f104b8ac0abe8add79137347a7ac2839adf223579f815d3a2f0e88b3adb8370d48cf95dc8d4c36a85787a62491e4341aa8cde276baa2cf1cf888be6a6c0868bf321cb4070d1d7ac74a36323aa4c91b85e5bc831288432c0527b610fa2da7c4659ff361adc4eade0d950b4f059dff9a57edf1c12d2b9b8e7bf2709941d6994f1f8c6258916276e668fb1232992199e23a4dfd6d14924d911862521d27b0b6b671234dba0a203d3d6dda521be2064d34d1a7c73678c76bd5e519bc32428;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hdc59443f79d88a8d2a31f994fc0a11d53f7bb05485f84dadb25735aae3044cc44e444df89ac648434aace0bb00f40e2574a7f4cdbae804eeeba9a201daa7941786c41d94b04c41188e30dee56c8e4c05f1215e610ad59d40f871de2bf7047052cfbf0c7ba5b2ae0217f4bc32bd61c0b5a15f1c51cc85720baa995f929629a48180ddbd8dbd41d0fd53916833dd69f4b32175d985461f2eec83e3a022714fa02e2c6f88220f980531448b04a17dbdd64cd859a23326059a480a6f88066bab5e073c2fd45c1975e7b848f7bc473d227cd9c37be6d8d8ac7fae28cde5a24a0a88bc7833b9eaadcf28f00dbd9804e12a23653afcfc16ed55058efee176f191c351372afd804dc4b995112caf0546c5c069bfae045619a94c8cd25929c0b0ce15ebf5319fae63a6778bb37d8fc7425f8ab659d74756f8ea8c417a1f81e85a307a748c82c94fd0d72712707fe1c7696914a827d155cc3ed6e933f44e364e59cf0e515701444e99dcfad62bdb83dfd354701d3277c59c043179cf7bbcfc7107fa426e4588c5a436996411839a2fd1bb7f8cb7555b9751d37c6448a47dee3622d3a84b0053c906c8fbcab3f6796e353f298d1baa82cbc599bb9dff3b085c724a095fe7d014d35a4862e50fdfb730080041a9608814e79ba19b9fb2877168e9d6383c24312086c13841b637e29c33fff59495a8f0b069fcd3762fb9329ccf2ce3a9eeebe868a6f90cd3a448ddb9f004f1c7da142246ceab1c85043e20d19460ae2e862b084a477d6766e4f07f2df5caa29994f6816f69617a7adfda49c138573c556b739fb0314051143e233f7f1f05a54da8a4832f811b31baa914ad0ef0d505b2f18b1fe244a808b7dece05da22e90216968f3e864bcf31319a0c6dcde8b827c991456b63486574ec4ea9715a327a22aa04b86970e4edb79beeb8770bc719299c01734a27456e961ee7d6eefe75feb396b1d3b278a0d75ac2f731f57075cfe3a766fd5c2d30c049ff15ee084298f7355afeb0053f04298fd57c4a8314630cd55505fadbf73df9dffd65b1ac00cc8488e8ab320f8461a828539c3301c14d32f7067119752ce98583f197f5bf18c20647538fcf9dd6dd58f564e479542efe55681272dc4f9455a48295812044e4134f850e8bbf4e8189d3fb2bf9ac65be6757d2a0a82f22ab68571214d73d5013b5d00ee9a1f2ff91bbac7a003aa3a19da14d6c818056cb493bc4bb2fe4cc7a00d6df71885fafa7601d96962049353e5a355bfd4aafa3d879868bbfc3796d7ebc48513a22082663600f913abb65fcacd4260b3bd38bfecad6cd307c69e8a1cab50c0c609dfde3fd1bf0e03b6444e5b1cc6f9cf03a190771307e7ee1cd6def34ada78ddd6ed5afff6321840efa575ed99739f50630c2f506a8c7c58894b5c363cbcff7365835375aa402f93968412670b7e91d5c0785503758fe4c51ae42cc5259f4f63b9606a4935a3e47f5f2526ba09c2606d99ccdb9a9c9e39862575bbcede1590935588a58b9479154d88786a0f24c8f954e09c2d5e285a79f8b5ba64f3b52bf178be9f46143ce1f01d9f2e5b3d5d8f9c5a99d481fdb31c1c0d64275a0fccc960282085c492d5426e1554e03b35949d09f7a534d26810557b3c192a6441a570306e52229ec107a549d482406fa9b6fbd66fec868a15178c312660ba9908f7bc922a84a15ae552f3d86c0ad99adc99798833df0d2aa0827d7dac9187dd0f104bebb29668bf8f0d0c337a916d6b3d2127195fcbe9ed6283f94d9e09f596c38aad0a9afe1c0004143a8d94d74d3405895b949a67ac6740da6b203bcd270bb0e31446ece64da38c7b15d9f4c09de80ef2117f8f6feb32e1631f4903a464ed840bf5d43a0dd76d2284334828155de8838703629ea95f62fc47c5056182f5af6cbd8a8443fdc64668230f9880ffe2b4a5e8c4d5a92fc81cae6dd6cdbc34aaddb293985c4ee6047a9063ea81d10d56cb4d59c6e599ce1cb8f4e8d55707297fc86ec27f26cb9ed313de7abc8bd5d88861d723f6e4effbd80a178de96be5df93e37aa3c179d74a0a615873639478c3dd5b3e5b61178e91f8828407e784b257efc1658b3d06796c47b96836d1e1aae170200578523e9aa3eb4b8214b0a17d4091ea307813fccb0561ebc305237e89f8598289285badf7f0e8b12776c668fbb001ad764da570571af790346aa29b0e38b86f4a3906bd9c1053ecd15a7700f9b590a86b670279639784ff357f896c53fb5a767ce07177973f4decaa72a00a92afd711e9ac2cd8a702bd2c90b5c03a9d8c619e1856186cf1d024166485c51ea6ccd017419569fb9759d5ea6c8b145563b8b84440368dfe81ba83290897ede714f94825bf1fc21a174f539e7d5cbcc02864fb762da8f47c4375db185820e7fd3b7bc93d7391bce354984e35390456b39988046b86e3706419a2c4017d673586b8b9f1830e4a2934401c81720fefac12c15b9498f381951968e60d5c9852a51f7db3a392bdfc0904f2675c0697bfc7071983ec21da57df9c84370b0c59505668ed152edd7d8516a1e9321dfb90ee7dc86ecbfff3a446f73d62ca574503712871af75e42e5f213c8aef0aab686ec5d2ccfc43e35829660e76de005f71266c0bcbe512b058d280f48f4fa5e1acc2b8a36ce63b91ac79bb515f601c0b0a7620737870747326d286b4e8375f4c715f67494e028ad84fb228ede6634c53216047c168975bea87c719dbc19da1167ca73c80cfc2e7520719e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hd84086299572e73cb74e83c858a7a90a73244eedaffe56c8055edb25d61fc51fd88ce6992cb7b022928e0dcd4eb7ab4c5109aa43da03eb3f6701bd5bc18193407f497a5c474758ec816acb0508df5f4305ba5135e7d4e056888e8f38c933d3ea0d95f985a6af874390d41322da000211227bf6ed0a8e4a9ba2fdbcd38ce986bb56f2707b05e5037f78bb8f51717880120650ddfb88d0744fdd462e9eedce51a652148d34254005f39a2562fa2371b3af8d33a89f1bb7d212bb69d38d91f4cd3220f09ccce98979c830cc24547bb76b89ae957d50c15f33715e22de4ebdc35c04e523830328418093d78f8f6449314486bd430322ea3c32a283e38237df654f191e08479fb3c40b7164b3f937c20ab9ce517d809019f39b8ecdbd16b990d28d3114a1b7454bdeb4aed8419f0a0867dfb5c9366bf5e851ec08c8c6f312e65a2ad67603b592319ef2737851ed198b0875f7876cb1de30e2ff25f321c3cd30ee87bed4d8e1d2263d53f4387d29dcc3ac3e484573c69a97784cefa2516467af8f0f763fba1aa7d8dae09b319ca70d0f49f49b14d9075e6f156ab2853b934e13de38a2f1c61121a005c74c512b6990f834902bbe706be3f1be0d85b4bd5ca941f43ec667075f6c998bb46180fbecc404395ef5553f759c05d82815734cd66376608f3da7eb904c9788261db6117b902b9139c94efe64469e0258a33dc73ca48630ade664d488fc3a71d9cfa4773de3d98817cae415ee8e560c5bd97356cc083c17d815c9f3f68ac4cf77d6dbe047b3ae3769bf22973ed30cb9c51b2ca3e670bc07b512483d40f3cc399974fe2da017cfcccb2cfc12cfb948b7c63f97c4cf475b8d5cb894b66cb0f94b962f809cc11c86f141856774a772ae4f5bb56b87105b5a20520e03e9c444572ec75f5abf47226d41b45e971ae604786a617fc9d05ce5c5125edf66004c8b2ccff80c5e238d4dc9f2e4664c2de2428e96ae219913b137aa05dfe3a5401a58da5248518137db5ee240fa01fc38719b4474aa09f7fdeb0cbaef2a02d3973acb8942e75c0c0e868237f44dc87431ecc01e60e1c8a55ff56d44a48bf491abb8f0102182b31d8eb1a13f7c32f06421f419951dea7a850149a678cae740b262b44eedaad1f68867af578a19d9074d533b82d0efc9a52e6707ea5524a07f93e0919ebe66150f87fcab949f1e8694b3f01614169475149874b5e4e77d34f8b5e089cb7a3982eeb5b6549a083e4346bd61074fd1f050c2bbd0908442f43a1cb23c4130cf67735667744b7f3313a3cf28dc187de576f72067fb22e6252d1b768c5481ddd39e81ac9084a3d2969376702924ae5e1d546ec3df6b8c8f9eed0592ca0453fdc9fa24b00826ef7134f0f1f72f6c4f9f0ab1e6b6eec5f201db45991b825e0cb8acd263886c2df5a339c5768bf5f7176db3260409e98daacfe040df24fc75cc2a303fb4c659b9094ae0119fa0a373b7b1db6fdbfaa35d4a14bde91e656fbc48791f318a7c5773c142f1a7a11a34d3b831973d56b5c4daf59816f08cc8b8b9657699fb0e8f10387e0c0a5a706e9f34be5d4879a1ad0a71daaa9d8bf90fe37f84c3fbb55f7976d1faf435517c03fb4c243d8333a7b0679e2a5bb07fe64c1e4706cace6babfe8f8a238b0df81321df05dbd3580a4d1997dc4bcd7ead36e8fbd4a1c36bdb668c2386e2608ba00b28efb1ed8e9ccb7c99457ff8313edb424d9585eb6aa19a880e2be22a2d9a0378a8ada323349289e90d132e2c6f99f3a0381ac5223a58b2c6d8cadac803ee5905548a3c6b6dec4b2bc53d1ddb9dd6ca4aa885ef9c30381b84256c6f07d30422122f3fa73dd5bcdd294592f7113573e7a97b3faafd84c6c60c84cb2a02edf91c17e83747e02220fa5ef723a1b92250bbafb2b69368218cbe5f84766a023a0efafe8f87a0514c2412a31535e962a36a05eb47e0fa976d62c963d1a250b213c447bc1034690d84e505dbbf477e26fb5b3d150b7f29d33a3af78cc9f5978f8bdacb76f6d1b58e2ae68bcd2d4fa4c48572c824a78ca49c73233ff72d4832ca559bf205fbc1fa2ef2173ebc1679923c49c35d8a0ecae86a390415851ffe81b9b7b9096624783b5404a58fe7ece8bcabed46bc8e3c3c3a1f30c747dc601ff01547db888335b9ecba9ff11be8e624366ab08ecc5cfbea1782a72657d9e7036c7d38e0476f04e25ccf38711dc7675855537323f76c787be7ab0bd7581cead041c8dc2dc92fae3eb02e64ae08388d8a4b50a13d77eed1d004db76d29ce62da20635ad973c89cc5302633b272bd79433292b4a4220a647d28e78017f0b4f55a4b4e08331dfc61839b33d603046685659aacfae52eb583bda1bb59a3a082621f696966c29bd3c5f0fd8b5643af8e6cef0620ecd0f9ab6d1fc9e1a3408f329e9b39fdc896c59e6466e3f3f9480a964672ac848778713e74a73c0fbcd1473f5eff3b2d7f09ec715d27d7aa189e0f2839996c039a88747ebad9a7b77680eb8aed490aa6ada160b616288bb8b0782ce1aa6e9c6f0adb55bd21fb56d228cbf612d73248db5c7a0e17d7b75c4d505085c70849ab3fef01e056503891dc33b7b6d237c179368881c83563c8083c858663ee34da7bc39fce703c563203826931238632a8131edeacb4c14a42ad51cdb35f9def05fa7277064167281b342b130b3bebe1766a56bc9b5b56393d6274e04e4bf377558d00bcb2ad9d5d2691d4926976e1f5a05be41bf3b9cdf33beb837541b9b0593;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hd6912893a2fbe3842950ffc05e07e1363847b9e056d3462fcc93ca7a6fdac4ba7bc18c25f115186fd6a184c8f8012c00b4d6412a126a426727d6e2cf7f62d7f1fb1e64c403f2199f9b1f48d032227b2114cb39bc7f050d6c4764b01283d3b00f9e8e0c82eeb4f07cf8c16eee5bac0e1e267e8051a1c5f516e030327550eeb2335152dc18f6f0f7cad931aac46a143567fc72ed5c07ec3ec9a452e80ed1bc9fe169a65dee96684773b341e68a746bf14fbfacb35fce25f434023fdec70afc245e5d1c4ea38f376afd74e56998e0c6c404275857d6e508e4e6bcd27026ce0c6b9742bf4bc6ff22a99650c99e48001dbf2f7578d06130fd4587f0371f94b5124506bf6788f2d0069f50848198350284d5aec880f0826244888cfc9d9305cfbcfbd96fe1c53a4a5921ee341a3f37e23212e947a09a45339464860b9c1caefbc014c1f978cfdf542c5a91270afb9d754c98444147dc57e911f0151bb86288971f42d2344dc6269f59aa9cad3f94021b9617fe334fe0d563112f3ecdf9d1bc968af05a8d1d29e52d729d3e57bc491dc48a7331571c4e3a72b3c20e8b09504611012242c261fd36cfc1ab7f7c533743a204230ddd9c6f4ab7711ea9a7c5233b180e86dfcd8a3f85af5f232b2af75a1c663c8fe39e797aa07f144658798bc5d6592821153eeb66494d2d29879e0308f1b9487146ded8eb8f098ab2500767a49dde049162eb34137e02be3d061bf24ab2d0ff0e5f23c4ad47aab464bca00abd0fa93db72dac84c9e86fdcd934414171327976b073bdd33fda2e8d831d1a810fc0f60d76eef063566f7e6d911143bce03b2bf0b84619dbad290ee1e614ee72641ece377f02f3fc872a002db5c733c4fb153c6d58ec5f798235b39fd90ec15cf9f5040276da4c9df7e8d93d6ab38bc9106439cedaf9f94407dd169a9bc97a420fe984cb3f436e77dbdd9f9c065e8047b4ff757c8fbb3ce7924466d652b7396be4b84556938068c3f95b84f30bd7a11dc6323f2d7afefb7c4c3f5df752ced9cee7db6c8e8cf94eb19e4e6998cc41325dfabb72b9e3aa16b0d5229542f5006b1cd851e79fa30f256ba509988a454c4774fcdc43256f41e5eeedb217ed2ce07b603fac445fa4fd3c0b385da600d17fff959820e997fa130ca212f0d3eb45c794bb8987443e4d5a8d16d11319e76edf616e0f49a0f9ca32b8eb434b169be44b086b6a6c68623a65e9842c98599dd3219790ab566388d922983aa985b15449010ab663ab2fb476a181b02211b4ef5b8dda000b3090aab13376128e137fcfe7b4fa688d9d8edfe39edd2383be6e0f5b17bbf82805571a7e521098a998bd50533e7a8e0bf722beb7d37bb474cec5e2fc78502e3d02d7a925700997bb1555203b483eb5fdbfa18b6938ac5d2ac2d5daca915bd01f0ef431bd345c7ac19a3c3be75a230ef8f5b799cf2c4cd68c54a2ffdb848499765ab259089b3a3460fe0c33b15ca97fbd6d97c3fb4ec909c92747c062058a8b64454646b58ed964733cdeb1ee230438bf22458f087a68799a63025f3030e5d667c98f281fc40c3e35e58d51a31275344316843238e7d8c54d311cad10095ec6f2620c85b00633dc27514879299156ff36bad783bb7749e4ec32c4b9b2a61b0ab8a0581bcebb12ee82c5b49dfec0c5aad84c708595b98aca080aeda3f36d6355467a8d365cb5629f6cc5672c878748c6c3441d6b1f6a3f96cfec01c633d04377138b310cc6be3e86d8269fcb43d8f2a5ad64c9b0308c6ca1d1f123f3c5566dada747dd2250943ce7ee30d1c92f247287cc978dd81ea4f677f206066ac402468ca9f3d749e2f33d48124b561731fef2ca6f53fd1f8145dbd4afeeff1181cd48f1096d7d9f7d1ce9f3f9520fc82b644d1a8a451b2192c168316428dc95775f916c1b960d851d691d996e78984f82a027bbc6657f32239076ff8a4de1685923a0b665a0e9b0441af2573f1a75814b852473f8a807696e69bbea11366657d79be0fe7ebb3cb8d1dd14a38b297c7ccb421f11155e58ab1650c79ff503bf67a8a2a42a528b90029662e36f40b395fe3bc4490af3a0963473124a34c94c96293e5685753b665a6888131f921d44f265303e8eb158fc402bd3bc184c104ecab2e5d03db4f69e0622e9631d065a1c1a79bcc560863e2f0ad1ca435065af1ec403926c86eb3de64a8c69ee0ac89bb2536f65f10a4ffeb124fb5b02ae6ecc842a7c4254d4ce16bed8b46054647df48649c928e5f614c226577d15bebdb77ea8a52bd617e02575dd3cd70ba87f3ee2a5d8d3a36cd08d534686905e2e1edadfc0f4245f8661e8959cd902a4b36118634c2679b0b753b68bf0cc97a8d3dcf1873651cd0bfbb2ac1ed822da3e4ac451fc0b78c355ecbf7c434509815e33cc7c825349fa1728aa28a99dd860755d8098d1274d6438288458614670d77aaac6d9c361a410a458d454648511a411e62f50a2a5f8bf9f1b9cf80678942c8a1e1a40a00745d08e99e4f57c42b23dde871f923afacc0143e8d6c19afa645cc204f7a7b714d7e251bb1fa2ef46cc0f7b4b538fab1028d7f7b929b97ebfb4ae20d2b0fc20afc8595aff47277895ec031917c3d404631de2e6109242d95548ec605620c9ef3346867ea94f8c70a14f7b3c32e062298dcfab420146fe204ca8b5d9cc2cee06cf2caf43d98f6301a5a4e9228009d512434a0adc36576ecc342a5cc97033b5448428106169c31e34dd6669fe413a326e490f02addb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb4804f67b1223246e5ee30cfb2ddb658bc7fa07c96086c1a9be39925606b8f3917a6e6049d505e4fba6d21006d251fdc987e6d4168b6571d67b151591f102aa6d02a43056cd8fac5a2f838e1d9be0f7c4f9e17320ef2e4745f619166b7b103e7afc086929738a09571eb9fef7412cfea9cbe78c76aa402724354900d71a6a62bd1796e86a85bd931c58a912435386af0f7fa158e5a9c3df5c509f08f4517ba929e0a23fcc9a0de7458e6b38c2975a6153bb542d897dc03033a66783772eaf79ed52d16aad56d508e7deb40dba98b0570d8386d52e7c6a1d2c61288264dacb7646ed79a9059ca0362e3e235070a3e4a1156d238c506c971977440dae62f3152c29790e8283c69be29d000c06500a880787767f858f7ac03972914f8cd47c48749bc79a33cd928c4e63c766a2ed4314e739726e4e72c8abde2c72c497b79a43220613cd096973a414f081e75d34abc24828a59d0efbabbcf3ab2b382ea279eb1cdfe54efdba2b3b36efc6b91131757da0210b738fb523c361b05a6dca6996bf970318237125bcdde102bd796ad7c19d97b92e0ca9ea83e5dd854c0784ae264226dd5b5db35c6a9512b8df184f5ca29e84f8f82fdc45cfaf0692d03065330a14a3270c90af44976953d4dafbb9f8c5228605d18356976aa79bb8768d2e698e8507dcfaec42390765b5769771264056d551043c2c91a9523652e42af5ba3618a89ec50df5b7bf554a0786fa64a0388c1b775e371c1270c640cf4a0841b610fd860afeb835b7c1cac3e23297c166d237c3aa1ceee3a708ac31b14aa20a49e62155ef2d9f85ef849026e5341998c6f249317a47f28b8255464ccf32e768e9d63aa1dc6f2d2d4165cf9795742c1813256da59929a6da8af63702c99383508096d68be3518456f8067845dc6493de68cdcef65c108c07ebb05b2791784e1d4328f31ff9ff37c02e0b478cecc331f9dd80e912949ddafd3b0c716b53d6f74835573758509bbe2effe1ff8715071b2ce06f5b9b82feed155fc20c234f2b934abc7faf38f16d4f51fa42cae8828e8649780b0752c27dff41cd4f6bb6e7a56e330e6b5a3465a28f7c07616bf0f23793b795acf107ef3f363eea4b9e9aa1e3fa693af8e2d437a08044644ecdb9f9cbd845fbf282a18acdce7dda2197e29f82ee75ff0a4eb2c7a3aa6d7914040eb8d783139479a2c40ccef2cb5cce51d786c8a0a672d7c28e437c28038ff371edc3753be400d098134e180082bd503e9723971c1abffcf85f1d019d1b3170d4c98350a2d6500a2da2bd5e30b82245d8123ac5585d119e36f166f921184c3833e96eb6266534c90c79a6e1fa34c7f66298e32b3895daa1ef339c4d4c7e3d719f5d4c0876f7e77cbdb4d53a648b6ce4e13012940620a79f1f57fd4f1a57915b51a72e06acbae9dcbd77c30b2893a873a7a31c03c3d9724b5b0da0b2f1a65ea45e9e55ed0c2e84351656be819b9a9d54d7040edc09727e9eca175ef49255c1af2e1e5cdd6a61f1d498b9f69493b73e75e47785e7579b385d123790d72440135a4095f78c4e63039cd27aed94957e01a146b7de4d77b71076eb6dc7fdb4407934c4e3b3361f14907d7038345245e743056e5dbcf0086977b862aa3960af6579c836a7fdf6bc6e18a94dfd3dd93a9212f5ec361772996778c761551a173d4f757855cd882bb54a307af07cb4831afb65dc59ace15b5eb734a524aca0d825e3fe180cef1381c0006378bdafd138085f783568009ad6fefe87f0a1122b17b934d930e31dcc97dc81db7c9060b3825290453ea5de646862905d89f73170117af3fd540ebf5b69aa431d77759141613f89c1ec3d06658ba33b83ba0fbfd4732cc5dd1060a33522c0bc601322dff0285ea677b4e7cc0d28c1e80469778ae0b01f72563eb25ca539db8955931551a709440844336ae086bb766eab1a3a44084879f71950f1a8561befb4d552be01f89ede5d16e5226ea0e8758c6db0a96d0b6139689abd96b2f028633a794c370fb625e1e3b59221ae3dff517dfcfa0c28a39bbf0595f162cb594ca81b93544828dc26cfd66ed32a7c78c563ced3f209ef750aa9d17e909fc97846671de979b88b3e4e41c860563b17785713f67d5f42a33ff9c3b22e3fe904a66e53b2ba0efd549fbb322362c76391ef480d758467760181a966fa1ed9d84c93f663c1c2cad09aec604fe805aade4792dfdda2e70aa5ff4ad4598e272cb2fd23b500a48494688ba90a7a44ee257f6858027978e7fe535f795bfb4c4c96c271a27b302592d7d3bfa2d46543c27b6d8fd83821a36605c02e98cb361c831538a74f3a1f626f758109f909a17a34ab79b1d1eb9f9ad9489d9b6daa3f3009cefa1ba4f39596fac4afc25f0630ded0bdac27d05d98423e25efcb89d49e5729fb8d99e317a1241789b9801f89ec53fa6d0110a7c537d5c3494e3ebe5a00a0c7565773f58256ad27de805544013f0b39d3346995503349178cc79a857d7e4c6e0a6bef9da40e2101c0551b2a445c62606b4687bba241c99768bebce6d77f2305155a2da63681c448bc908891aae0b0f990f15cc872a3b485c95263b9b529823f76f57029528000a3be786714ff21d724d8d151c04fdf1ce2745d87fb1d9782e75bf50627da6b44ec7c2f4d8354711f5c7017caa837087da781544c1e32bce24fafce037deedc281629d7b0b28f4baea3e333923cfdf9a35c542c70a14878a3be0f7e053421ccf810310c07c53cba5f2682e9b521a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h20ab606e76b63fc92ae0914589868e86ad5e5b9f0a9510c91ac4dbc219c28f21feb2c1847c1298deb3ca37baf15843f28e6f42cba613ecb97874486804d97128e996862f7ad9b632da77c60c14a75152cf001f1be77953d894f88d12e818e9d32f67b52e250cb9d164106b960fe0e70c17b398cbb7461cab3929cdd7f79a8c2908ba1f6f30d394a553586a88b989558736b0475687ac8fdcbbdfb4e59cb1809df6c2d8d83a2770043321c12b47cee14a461e7882423fb58c772b630b89a693adcfbac31a3fb78fcfe17bd99b9ed87186dd2e680d93b17f67ff4acd3a741b8fd0a25b0d74f0beaa1da6d66fd7392e8e8d9525c3e996cc281265730e8b6b77b413890fb2908eeb3fb5fff48cbf997214edf870a381a08a08528831a68f50ca982e86eacdf601ac44eee12f2ea663bfd223fec958c333d4b5e76244dea5fd01090f6d5252a2f682a9171b701b18ab77792c64c91476bd93e16580ee87dc8e62ac23ecaeee323baf5bd3780573fbc6dabe3a847f98d369085256c8883f37f5977400f237da2d8a7bd75b541dafdcd54d291d1fafe3c909988a17724c8dc42bf5bf4a2ac598bbb884a0c3898da9ac7ef47cb7a951d544e735dd6d63b86e4cb73fc695a14e555ac40e72b4355b9f9adcc2d02b86da172655e1378ba6586fba40df804bcd77e723dbcf277148bef0b06f7538f8387a5b49d825ed4be4900c13f5de01d851a3d68523e4ec2bec59e046105ef007ecfd2f16ecda21bd9b79812b2153fcf7e4c79f6cfe33bf95ded101719befc62375435b05265f833bd1fb19d5118aab47b61f067db21e97f299b54382b158a568ce0671ca96983f3dcbf3621b393f3cdc3914a7b56146b49f4d9e893327c73c7b7a41e576f7e63efc208ea6db953d103222ddd414c5cbc47907e855f6a08874bef3af2ef10af70d51e7e8a93e704a11f3928e483e9073620e4c28cde60c55ebe0ca218e5fb16802981a4ffc2e43cbb7caee68c70b415e996d26c74fc3dd1671059cad848540421a29059c716fd17e156bd8d507bfce427b1802fb053bd19f75207cd3e350041ec339fd53ace8cdf63fc7f131fe81287786c5c55831334b12d91ff478702e309aaedd92281ff733385725562e0e0bb8d2103ae52fa5dbbc65d82539477bc9e2744e77a68869b0e95241f260a8419d1320acd0c14ffcc20adb3a6bea49fd9facab9f1d6bfb568c1bc5e5c840a67a60a57a558631b9f91c43574b33d9ade62438cb3dd6f39e643095fe68209e7726517061df32ddfe53cf696d66a91c102623fcda96fbabb9afdc69a6b2c3c7e62a7c84472cc5e27fbe1e76c37566b36276407f3f2b14c35cd54899b74c25de660fbdbfa33ef2a2c92de22cbcc0421d781b484a029449b53965ede0e88e28a9548066cd567530e31d5945ea767eb4e3963237f311c1761112078e59d51a7a516294975050e341280790c48b459ecbd1b461e4877e91d386a46cf526cc5c3d8bfe992de4897ba4d165ac5f8bc5ca423e3d0fe96808aebd4e3c31b3cff46e51f1dfcdd560d4d5a60be20e06b6653a058571650305e3ed404cdf5737004dd3a197a3b87513d677bb205d1d2ffce6022df1dcc196382cc2f2ab03ebc8cbac8374a0fa5b115d281e8bffbd6e52ef204c4ec972b26124ec65bcbb87d5e52a4ce134f1af06c5f68c08e194198b6c1e60bc24690aaa00007dddf91d6a202d74bda02810cfb68ade363d19a366417bdbd4a0705d05a63b86a0227f815a721f0ad7ab25826a050b4c9597ca444266bd14d13b1a8d90cebe56a156403b79b6016773b02efb55c7e6fd8e1c1475e531ede413e4838cda8fa92681ef16c86b82652e327705ba3588a53dae3e33780f087c3c1aaaea58372deef438e08accb13b799bccbda504485de814a36663287844fc7cfb765a272c4da3b737bc596b03ec96e5a402afcc76e410b84384b7e7f8d41fcb35bc41c89cf504c2d75ae847d3fe88791a7b84598262ddf55852a6580e47b28983c3c9b21fbd07270ac55af27bcacba7753599acd1731e3a9266cd95c83efc375a4dcf1c41fb5f7e4c926a2669cffbaaded9b6d67618f96860a067051b8a4ad1ef33bdc3d72cb27d173e142507c25cbf7fadcf501933f3c8f3525277dedc90a50526bdd810f7b3746bd2f289a59e329d616e9e378f96933461fcd14c82c27af1a3407069bd19fc2b7197a5a24041ddc287572cf4face8d2556e27843cb9baa88dad2abe981451a5357018da7fcd77286d032178bbf4661fd4f1424a38dba9a7a9f09a3b541eb8feb3cf1d42d0b93fea30f038f61cabdc7251ea1cb61ee2d02298a7c3bf958e43b5904a49d935ac9fa75dac6ae177916cb7edeb8efeaf2c048075521b4e644a797824e7ef38ad35a6a8ee400e76392be2769cfcce186bb7abc4935964b7c246c4562acdd3adb57ee36a47c18ef449c605335f1fae91e6ac62044b5ceec061596b1e2809baa52a5d7391f789f10c7f54df4f3104b79e6049e3341984c8a1e3908e003c937078971c1172cb593b468946dcbe3f7bbf77802a0d38363a38f5b1f9326241fa394bd02cf65278a904ecc0f05505aeaad3e73dd1b9818f83fce1a2825fa469274a03cba531f90a3ee2d19a7401c2f762462a9492c7515917b09965c59638147baf4cc8ef66232fedf7d5a3b9d3be0405658e7a9d00af4cc6685966fdde20884a3d9175715765eeb9988221b26e596e087ec90696497f0f4a554095a68e05ecb18c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'ha39150d70389fac57968f1fe83a0151c32932abaae2530ed0e9f314ff362f3797c83801d6bc7d3eb819c2fbaa79ac86824cec4d5240e7bc6fbfb393bea814900d93e5d59ff47100ce442c359f9a2d9ced0a72be336438c23d3ec365ec06eea6fb3ff6ebc1c44df45d296590c268b920eed812a5a3c0e18078053b125e52c3f37ff26325bfdde30d3c32cf78cd8ce89ae59aa113c7bd5a3b4a017a56f180b67f022baafeecdcb0ffea20b2905ad472e90805a92875c0a69bf30e35deeb4ae4ea10bbad5aadf88ed12e9cb50a77d218a96664d1812fb4f567683046ea9ec772d5a1d28bd75acf19d42981bc610764e15888f03b72dd7e94fbc4c49760478bd1329ffa394aee5e8d08fdbad060e3abbbe4925ebc0e847705e49d6468eeab9dc7fc664cd9a439301779283cf1b31f4fb33fa3dbaf81d7ba3deeeb457d7156a934406e0de0b2b0a0e46acdd7c982205ba2a058f5543352595c6af7b7218aeb63063e9449784a4914934eb51e00b67d21119725e432c5e834d1f87361c7a4dd320832c55f60185eff9132960328a4bee60fb710384740c276c989af6edb5a0570f19971fa9db6228aaf0df68158ccbe6a774d6a3c11bb86e033c06a91093a1c2d4844de5f8db02a06bb933aa3bb977fabd98ec4c92a5330d8aba2318dd6f2a3da6b48f9e1ea981145ea60afab75c752b60b6d87c2b04f956d295459da6004c99629247a8efecc0da4bb37678bb58bcbf2dc6873b7e83148a617988a8365721e01a711863bbb77a8e6e57c028fd723356a407c4b6c818165488f857ec3528c0cdf6bb815e8b114360f8b288ec32dbe42d5efe2cb9c5cbb8500b6a1b5637a2b23a0ae4ff50e65c8fcbc6baf498e9eb329e2a21a5e219269f1d0cfcc6b423c14073e9f3ca80f8eaa084d81cd61b3ef9ebb40ca7b57bea12f5704c262ba85b441dbca5d1909f575c14ee20080fd5e9944e73ce64099fbc0a8ebae948d310a78166b85651696ed3a75439c6cda8dd15b5f8025be4c07d78f6d995c82ce2463db34aceaf9a5f4321967abc344d52b202bb65bd27cf3acd65818494657310ae9907deafe4a37e7a7a3597b6bddb2a04c2616bf46a0f3b426a7ead66751bd112cb5a7ce3bc99bbce78c6548d44f192badcefa2f988282e846a2a78342057d8e0d395c3f8a34936a8966e333a0b2d0154eb7d87e0c6bbbb0f343d1bb94c4e73d90ec92bd63376f996320a13f712b221c9f162d50e94e76e926c53b443094106f1c04536ed0cd046015ea3bbbb2ab91a735235a1315f682402495fabf9aed942c7f0eb27603e3c145c935f5e53bbd92dbcd1a02afe49945948fb3f2fd716f1895f0d67e2dbc4cfa63d5a5d973556e81f0d665b6c96fae44c088743f39937e55531fae2d1e955f23b1160c3ecd7118c5f41d135ccce9351ef0fe9f7d7ad408ed072b5f09266b4abb5d20c574edec6655242add302576dbd689807c2fe89ac584efafd019a3977ac2e4f66e69ccf19bec8d3620e34ce5e34e7f3097f87df37b6a4a025eca3701c50a6b47aef517e214212200b8b8cee70d39e7655b1f5b2b28af47580cba7c28935d414654469cbd073693fb415ee1c9be987b24833936f972253876044790182c5035d2909725e79591e29c89385cca2536d0d67a006bcb849b6322bf910735586b87dea3c54e2942de72a7f001cc5a3c207522a4f4d5f23786296bb246538fd4a2f3aafd8f2d5ba6f1805c05c37f94f723bc72d52deb13db3cdf72719f245f7be2fe65f4853c7f55133caafee45d99702e40c3f53416799c169b6330d0d85afd042a54972a2e12755f87e104eb25da3ad1eb8e4d6303e3155526f06d6f0b0830aad63f87188b9205402b3868cbb118ae9a82c253308b5b346247812dcd799fe49230e343a8775b068e15ef1baafb7d390e6d8c89bfc7220905d83fe6a8d1989b63843ba21ee2d07adfead0ced3926d8df1a703c0e43128b92ecc39723b7bb7fc37d3e6c0ea32df08264b79add2f89cabb6330b1cbe7ed8f079b94dbb953ff427835c842fac25fad124c44aa0a98332e631721824d8faa56ca9da1d5c3c5649c4f799213dca9ac756bdac897967f6b6c0d3b073bba80e221232f82237428496b92a9cb9c32e62623f1e4864a95a60c7005697daa64f6b8f79cd26e9860e68030dd268172209565e3fcce763b1870a187255fd6b617b7e8c36aba2889b23885f4e00bcee9de46d6c94d88533de3bd16f83a32a3f837f7a40303554a3a95ad76d4f8d87806308940c9d8645254b313f3332d59eb28fa7929196bb6d1c29b715034f6a3bbec5292beb4815dc62c5bbe313b44fc101a9ccce4f16540ada5bb6521882ccaeed84e705a6aa6ef6df0f4426e782709e28a1f99b2aa4fd9c1bb4ab39a1cbd0691fe63b844c22315e325b90bd5ff202dbc58bf4e8b32f7bb4369773132b2396f27d3a5257a854711687b39348f143bc91c7dd3ad545d7c7e3ad8eef6ef67898a510d5dacda54149e4eb5b0ba99affddf0f11a8996785078a7bcc300870ca0d196d2d1fcf7d3301838cd1d2f81a1ac70d38d645f0b9ceba6737215cda12141aaf8be31787ffe8cce9a6bf48cf06b1e2c6262b7086966bdcd7651438dbbaedb5dfd3efe78ceb1543476a80e81ef272e4a3cf691014859bbd81453ab2fa31dbbb1ff472501a7fffff5c27eda0578f21797a28e9ecbaf01989f23320012061c9cd76ba4a260ca50285e7e78d84c94130ff9ce4be76aaca489b8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h33ba9ecfc4e470370e5c471b449df3b7bad2375e87f3bb97e645701d9305c3a6b280e4773114b85380945d71331de6bf16cb677cc10bbd995e8f21aad301a4009b9a60e94443e262787ca0c30a42f07d54ca132f01784ee4dd14b7201c9fa22eaff66a25cb64194f00d6e50c2dffcce524c9a044ebf80480c41239d841328423537e5f22359997db7c510d8a9084e02975274dbb0f5699fb5d0b9ba371507e41763a2c9cd7a326a95d7f0bead51feaf17ab947bd51e8bf201f5dde481322b2adbea9ee437f29d99fa2a0a6f905592ba9d6e924669b98f90b201eb3bb9ad25b8dc50d503105be133a08ef46b2aace0b2db175a0aa71bcef50a9ef4683e2fdc90c58fc1146e7dc11e84076d84158baf533cc889bafdef3ebaa711feae552f96b87658b87549e2d97134cba8f015773807718e5c4fa501963b00cd2beb1ab5813b1579771f3909898772e4713c9d45136d955ebb2a64a4f69b23e1141ecbac8fdfea69c371320662c25ef85ab6f6cbc99c95f24db9b07cfbcfcf9df20d5ecda55148095e9e2d622d569d8e6056c74ab08ecfa9a3d7296cb0b7dd689e36fe5cedfbcc417184be0ccac484e3b963554e1db108a9e8eb7147f20e323359b848ff44cd5d6d0e41543f3bde4355cc51776c09895272d8f3d56a0b30eb27db250263711af7e99328de2e0fa0af38b61481da6609350e464f908654be9c60dcbd451f7ba4a8e7c2afe5811077359d5d509f6db1339fadcaa9afa0c8c07a387c65086a694bc90fd9fd4d12dccaecad6240eaacebbfe306e2884ea21e22f71b334fdf39f5a33e2f50d0b4e4c1ea720b3609d7803ac177fd99805f9008323c6e834cd784fa3b34a90d044e59d65dd543ff249b2a9ed978f0b561c5c0531c6f9fcc2f8f901fb339ab8b981ba683cfe944d1ad62cfc52d39ebefaedbb19c271e9cd2bfc0d5da421bd4a98836688c8c6255adb910b605904f57b9a0f8468048a4219cdd30be44b824593968c8a798716cbf7ece27000876d3e5c1303e2fc2f19edaabe1bc289332891608591d7a6229adf0471f06650a6feaaaf1e063d62b1579cfa1d42a33e3b54df108567f1454070b53959fdd1dd33dc603752fe3b1699f57d187617eaa72d2ac93669d952693010b26d50c723e7560200ec7bcda1314d9056d8a892d6d928198862f2c99757a62645cf608c424af9a74e4e708ea1e0bb5ff3c8069e3bd12cc44504b02cdc67147473a18f4aa115f7db77fced5ed7182883900e9dd3521a5c90e4671cc524f530afd975c5d57ff03f17411f5fa4d339cd449d4920fd4b8778d99e90b6352a7e9bb502f64bed456d42bc70a005accf92d38d4556fd5044a6040ab7883b75a1f67d625ca3cf9659998cfb0f844098963a3dd6ba1923f567d0b4a51972a12d2928b9420a551c04815af40894adbd04896d24b9e1ae972ab57876a6cad81dd4206a424a2ee9b9806e6fbdc63ce8cd84561f4fca421a013a1aeb38b8172a14904736fb02cae432123e560dbecf43c074e7f0e9576e50f6c0ff5e53c7c0a52ef26b42036d86e23e2775fae60709e1158b8720bd2b74b92e618ec12b0b57a24141cbc3d639896b1ae03c3dcef093f1ccabc94272344e63035621184b23e0188e5642f637ebb20ed89a0e880ebe00b184db7c3dd2992977f366337ff963c9cdf70de0b145b5d775b4eba2159138b9c04fe978703b2d87c0951e8b08caeabf30b523ad706424865b1142dcfed46f2a057d2ba5104441974b44bab294d92ebd7d58d5a1a20b233665ca1782aa16e83df8c1e3dd241b7437d701eac491ebe3bd2f5cd9027167932e868607c8959616eeb2b825f0e18d62adcdbb9059ee322ea5f174959c98b4f256d42f58b895eb0260007b17b4907c8c6158ca07dfa69ad9ee58bbe6a713c41a30259e96aa65f5e26aaafaf6f88808bebadeff3eebf86f5ee818ae6012404180dd41727e35a640e42aec2cf136cdf98df85e8174983ab97192b8790cfbffe733dcb874e08e6e211827614ae14a4820d1d0e7904743c6817745b0ce558b42d3fdc40d7f4fc529da468a53103c139d6752548cf0ef1d6eedf430d493be0122527a7c9ea6c83b441296a20e9570f9337b3cc14ba81ca97817243034403505f7abd3fcf14da45a9d821267141776a994dc183ae61bafff4dee6235e2e9baf5b28aef630ffc8f231b1ab7e062705dc7988ba2c15b3c84e4c74d193e6a3c78d970f7f66ea0cf9fc42e8cffab1d1e51f26e64763e5dea7f557fb38d6ca491f84bc1a4315bf1dcae87156fcff9ea1a15a16321b0436b11b72092ad172ff42495aa133ff5c061760f0075a565311434e7965906bcb1f986e60360bd786e153d655bd7265166de982a8dbbf8f64118948baa1e1a99bfda2e387c3fe9bc2bcaad2f8fcd3f0b43cf65de9bf1f42407805eec1cf41c61c1e0f48ab44ca4cbf9b9ddd159f192e19971f75ec53fb91e1d195a2ac9353c0fc6279aeafe5144afa54c60d3bfcfc8b62433602456a92d12b8b90dcf29f4f1fbecd9192986f46239b4619221ff4fa438a995cd88e11f983bfa4acc134ed6816403c062f5fa270a5d303d50c80f3a48f0639c4c700f3a47095ba2e328605995eb1be326ef69495ab8317efd6c3e70b480544809c1abc9c96cd8cb5352b9b4748043b4b40a5ff60c4a701f11a182d8952c652557446af478a1a31c0494f02a08adcac9f8baf53ab0ec2eec859c0113a2c1a4609a92e13c499a8358da1b76030883;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h4b8cad47e1e4fe1e3e5dadc87aca85370d0e7ef9032a3c42277990a688237f7e504e77d033384c122e97ac9e915babb4da0e8c8ce2720361db63f7c9e95851a3e22b5ab03791d18c1ff9e65e6d01f1c51e9a2821e35e2fd0396c3625c90172557accbfaf5ba3737b317709491b8e6d53e21c4b70610d7fc4d966124a9f73e5706defc81d15eb2a3dab9a51263a87c5dfdbc3bff0b170092a5458b1725e2297c5bc4a8767b184a012f8680646e6f4b892db66ae655be8bc8c1b010ef9f33e16db42350a97c0ed94f287c4f84cda8a4650716e1d02d452431c7d4fc424d20c1aad51f47fdf7f5abe77658b77ea72ecb95c7264c5bf78b222f0c2bb16752c2ff57c265dacc555c93f5df5b1940aeec893a47c4fc70d97855c51bb6c20858651c990435044c04dd73811ff05cb755ae8aa805c5b61acd913dadeb3ad5b2435371f0445d57f8e7298a8599c6fd88ce814cfb21168647ed11f596c8cd5162db1fad70b1d845371be2d38eb0d7e0ecb62fcc2c42b617056962492f06b7cb7ae3f01ad4974053194e6f11979e0290c8412bf1eb306c11309aa1416ba778f0875b8f85462a3db6db3f67c58ae8477e2a8a2f3110a1275b3fbd0984757ccaff133963cf7ebb162fe6f976291b4619c93ac8c880647335b180c1ae1e335c2d44701553218a2f6a22eab6069e4b7f2e477085d79ab19dc26ecf521a325837590ff4f78912280a4fd7c59d678bfca9a11770d09c7e48e864ff86bde7b5841b7c264d0d47a103d68df1234fd4ab90c03ed8632d25be82e2be291541ccde58c53262fbc975345385567e6b6cff35870a87713095456134f2458b383b3d8983d66306153ac4e8b7db49a030cee71cb4b2fa736f16e629ef09c78adf9d49292cbcf84dac7b826371e1adf034ee6ba7f9347d9a69a2e7818d0f533a7b62f2a602fbe1574cfecce7723faaa7a541a90b8aa411fd111c1e46ff93a3aceec94faa05f2021a611c3c171169cd78b70d3316cf776d8fd53216e70442b4738c3f6aa685d3b06aa314502459f8b1513210121c385412e383ba0447b6ddb1c5ab571c6f9031a84e5fd72aaf3e67ead091a19b17cbe9c56268dc9d1bd026aed48c4d3792d8aa19962c5100d5b459b580489cd3b5f88fd7d656f0b8b5a924f9b7157ed22a077daadb8472732fcd1de0468745acd1b23b438af3a20793da205bbb3f3c2ef0494ff7a89b60907a66818507d128f698ef9aa41a7d8be839d6793f9cee486c949601c4f6b98b61e43a56aa2bfbba86871c3649fa131017dab76d3a0298486d8c78a359ce65240bd79daba20a038a51bbf5dc069478e2b55eb4b81d458de42c411aeed49de0828197fae309eb6ebabfbcb9ba8aea05828de38271326b2f0da3f74ca6d211759634fe714998d71eb42dafa2a532f30e0022dae58347b0079b871a9593f1f88365daf9f570cbe3fe22a93b9a0778c1fff4f163968f7a23e37bb270224da85376935daa7ea48e466f382e87bcdd6e52cff20ec228e80a05c83643f512765b7dbd99fd735e6d3073cfbeda89826918d42bd4880b01c48aa86c196a769d5d21ca09b8ab875f9fe71f50d8840bd038f9113a7d461a01595bde8655078253d80dbdda432e8096890b4fbd067aff819555380195ab49adeb706ee94a3781e726bdea3ff30b6799328e165cefde412e190049b87fb32ab836207f98f140534180d8fb6d6954aefe8bae2b2030dfea07b147de0f3a136b51001e06e7e9b58ea5d1e3fc4baa3ce321f4f2a45d1b1d15ffabc27ee656c24c40b93926fb9f161bb0fb3a466fbb96cc9978e6884375b8cce1079248d00ae04e842d2a44059de4a3f62f5932b2cd228b1d836f31553d6491239dcbc9061c9b43ceb2ebc5fe0abfc7886c2bb11328ff029e4ecd36bf0417c8cd21e6db8854602e2ba9d4c1fdd471ae4854d2744c83b43209058a4a263254a7d501116b2bfee68ce15361b01b8369294ea51ead99a2f31592f6a9f8210f5e7ac93aee5f8d169a8bbcf549d3760ce41e3a966eb8a81c82fb2febfa735f7de78073d95c4cb1b1c5f785152da7d27a979e28d0ca89235aee0beee1741528eeab6478665c1f6a6efaf1927ae037f464d7ea75ed00780791812736a36945938d789a35261902087a7f643cd8fec557563667592050b54a9f2adbfd5b575d6208522a3c4eb2b7ab6bf268dc484ff204945457bed66268d20eef6aa288a3294b5ea882b50fe20b21ad39c3cceac4598d3c5ee6ea992e48effb44d3f2b31346fd2cb19502bb32268cccfd1a1f6b744b7b74d49277be17bdc7fc4dd66f2722e08dd9c7529b3b94cf3655447948bfb77decd4f89ec05ffc9bc004a6ab865cf029b245f2284282a02ae1660feecb0f6d7a3ad4126e91c6ca357ed48cbc6af3f09913ce97d488afbf6cc3ee8f5f4eb52a92f2db9c0e65ac4913ccc1b4e5b09f25e052f78a87eb6647590e3493d378caea9a7bb3fa7a0bcffabb1fcfb5c844c2225a197cda8ce34ec38064ce714d65e92036d00cc4cdad0f546defb59a9390f954c7b6a48d40c9bdf8a359b06597e447e9f19aa2acc68b6cc24eb82bebca9a07e1e71a3e4c3478f6515b77ac00113466ee0a722411b09412a69bd670ddfacc84a204919750c33c7d4713699596fc27ea950787fbc5431a8bbb2210190d8ab43d56858d3be0a7ba6426d9a5ae657f8c5979671a6d43f07767663a3a47e9dd01c86156e05300e1d08a92bd70a728f4de6cbb8554ba5c9b53;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h8a1b3425773b2ef971adba3ca0f4dd591e3e553fe9319055f1fdf812dfca80c65c815772cf5ccb462ce2324611eb0d745e1d06c2191a60f906a022bf891b22fac8ccedbc27401d9bd806bfb746bc1399f53baf69330c8b555b70e302dc21ef5082c58152de72fdcaea2d82a4d6a2b01afefb476cda1549e5388239efc3a69099d6ccf3b1f8bea9f2ef1c581c79ed6bb9585e447d4b97a9c99337bbeb44a04c5991315569d1a6610710738afeb904655a50c9b1ebbe4725f507b78640541178da393e4cb378ff2c42d11dae34a6ac607cad566c80b6b47830364d60ef7cd699ac7aa77c30f2d905c88fe8c965597d279af578cc524b19820dee3b54bc54ca4556097d8a5861252ec52446d47cc5fd0e2f19f67ff8bf680f1771e3edd5f3a103801091a33153f19a770f9e5e8235047399f5adbc702dfc74dd28d9d9416e54a65de95475598f2a01ce0a91788555772fcdafad170fd74666ba8c8b8b536d34b7915ede6e839617a69199a574e33d542ca0499ea42bd64da148bea05f80b5a1de3b37632bd921a80f6b4a62d447283654e1892d6f7b5429be5f618f56e610bfc5fbfad188c37910d4d655d1ea6431be630b4f3614c4f407dd5d31c80aba012a63d70e9cd3757c71ac0c33005e7dc517d7bb3b5576d825d15f79c1adc687e6b9c5ddf352020f88ac98066049aed6defdacd74326bfa595e63056b131161bb19f82c654ba3f1639b1b2ef18cc4c565798f2e42ed607905da467f93da3119266c66413eb245904bda5cfaa229a7ce934048a7b7fdc4295ecf99b5b4c78d12307794867d803f576d5798544a21427c7356efc7695b3329775754b84fb55fea5355296e5734cb1372760c3a64418a4811d2c0d0ca3f50b00c2ca68f07658e3a040416a39c85ed86ad8744f0662241824e79db59d5f328de9eb27fd6c03d16b323ded651fd4db917ddcdd9632980984e59cf7db1c72ecfc2597d35a94a5d2d0d9e9c6062e778d23e52fd2454ab360278027226db6eb679c0c73992c4fb73e2b9a4d9e8955b6157bce96ce449226c58b37a1a6f463e172c780c1b6c7ff8014e75e7673c8406b5f518edc5a1618cac2d7d444d77fa11e03d39883a82fd1e30b4756acb605e2dcbdf797ac3326ca219dd1787d0b178e248301df23c1348223666519b7c7774a42f71ffa8654ca6454c12495f7f2a0ba3f6d554ff301e2f6a7295fcbb8f50e3e0c6f69f1ddfb88430be8ba863dbde476aa60abb8b11bd706b27035d66b2fe746e8234ff9a545a78b7b1b82111cca0698fe75bc91be96318d442e6e4ae502dae4f62a0d0fb5918d1215a6e593b9fd0c32080a94864415d5f31040966cf1a86bf2aaaddeb23ca721f1e3979f93ef3017b2c73f060b7ec5edaf5f00165d0c94a99c67e704d05d60f74fb6c95a2b2f7c7bd38822cbe677e9e6a73b7e12f751b1b9a91f2cdf3dc2c20bec24d2d5640be2a11de7585bfb13a67d3167d1e5832efb491e75d77ff27c9e8b31ccf363c232f6fdfaa1d7b71a8533b260320aa750700c3543eb92c4a6f024a543eb2836f281ae45d1cceed51175c5fd81c3e9207601d7af03cf756eab060bb5edcedcc5549b278d6ca6201329449ba6bcdbc359c7d0ccc26c1e0712c0a56db0bc2ed89361da09899e20d5c6df20e2b20db075c3076f6f40c2907a87837c60600bbe0cfd03198b09013933f4ebc0c7878501f1d7c91e303743b98eaba9bbc979b64a4c8efaea3d5f1212855b4c97fc74b4668067a646b2e4580fe6c7dd1e61e48d36c47a9cb21d7edbcc447cd240062c423399ecca40fcdf18d29e82c40fc75909dfecfb6e315222e0632d7e737e4a21f8fdf72394be49b7e73c31bc1185d80999309342dd12c3e758e7aa3ff30c4597927b4f2d2eb9f8bf4f2e6f18d5650313a865376a2ed564db37366f779f00f4fa6877025a41b323a92e9402257ef8a5ce73b01b75bdc52b543e31fc63caa7d5d761ca78fb6ad30eb6f1a8d439fd06f01ee5fd335ef90bf19b2bedf65baccbde2f585fd2522a2e2168c8e3d841ee0f4e85fccd388c3c2e59899306fa6a2e0e3d29b6d51285efcbeda7f70a2a5e0599ca7aaf7c93ff67de5260f6f1821b8bcb63f3188ad650799a07345b7a1ac75610c280a520e73baf2fa1987ad42d70f372bd72826a956208504830b58f39eab93695b3124302b384b6610213fc256f3ec2826bf1fcc17ce09c3e8022821661a1934483333b98e35e54793039719197307ac885b3e74b2259d5cc3bd48b8e62aeb652c9a9d99b076e4ad9cd09c250bbb61ccbf6a8c97ad391de4bcd143e851c723b8ee9efc0e0c6346a15ce3a494b5a742e0c35d624c9fe26092cabf071927d38e4bb3bc71555b9e38e11819a5d8e65d003980fb8f9ad1fc2a0c5598b4d81424119a888b27c6bbdc5ff45f9a603b299ce306d35f5d6f29960f3fcf48db4d689ed560cc1b655bbaaeec13e9ee32b5ce486e60ac45002b2450fa802677c6d15f1f0d3e4e05ed547c2451063ccf77583db524ddd1b590c897effd9f7494ffbac7ea3f326d293bb8d8ca9ec642278e8543bca7b4153bd44b85537ecef6d3b5754cafba962ba98487d5f1808108c326922615712322f01423b4ed54571c27e6f59a3c9241e1e51532d9778238cef57b6fef25bc2e8738bccf5aad2f36fffe26ae431847b4f14615ae6efdbfebbca9cc3cbccf123f6d9eea88abe77e1e0045d9f2c384aba9d4caac1df9837b0a709aeb47cec456d8dd71f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf657741e3c0bad1fffb9bd1b2ef474c0ff53b83f424e595456adb1d9d03935e5191aad5fa23ef77bbdc37a59ab4f2b3a19a731a6f2bec911b19c034999405bd38259d6b014f21978598bdc25ff893d4e2bf8392273e48390e30d3e190938dc7bef6539fae78be547d30e0249b4848a66fd314379f55136c949417d7ddc5d8b56e455ba40e76593fe67d064b4981dde43e16d6f63255086415ac0ca9dafeb14b94bc184f69c9db78dbcf144f21671925fe03a8f4285ebe5f1abfd1c24366393cca7af9de8944c3eb8f698af3e789bae82e541c6446591da30a5bdd6fa0e48040748a8113a41201b31497f9181ff545daa78ef68e05939b2935de00e88cce18ac0fe5bec5c541ad674424d214490249d9f4187f3e2bf4272f0aeb35e0ab0f257708f9a82b626f4fd031bfe0ec97d09316fd2cc9a9800cba1dd5448f6ba3376594bf9d5b6468a6e5506eb010a4151c76ec62eb252e5d78ab625c7338b7bf9132f5bca6bb637cda21bb1e1940a2005d3521ef1358cbc78ad7d2f80285e5fdb2edeaa11aee802504e279a05ba56ca884d96ca6cc8b372f643592492258f85c4ad43a6dd9e0268be52d6788433a155543b279b442ef70832426ed4e51183f302407483250c30d8721f7672f5a10a02a78dddf597851c70d250523e871e3c2bdbe0eee259db802924b8740716d12cc876f37cbf59e5e8cea6f3cffbec646cd4781eef8ca7cb5286400069d2b1bc2997c5733e2d555e44306546123434f96471f7edf36608efe2debc5ae82be1900c883f4221fed79a314b52fb80eddf4a57b95a87e3b77f443f95b2d695638cd805b0cb0a088401f7e2bc423edf4001a167e1379e97b05192311b5e308c574caf32a6b8170af3e123f907a850c81c32f0317c8fe39c961dcca9a8bfaf28df107df191e6130cda836d4f1ceaffd807fe78557fe9162a72d287a112cc14e74d61e5931562f2062814edcb65c447d33ad991d18c8a7ef08d8d6950a689cb37da209b696094199c71dcde55a2f52c8d722d56a0f2064c18c95f177490b75b072a24b109343166ddd6722e7afabb091d2ae62bd9390450adc4ff78c41dfb7570264ed221ab7400096929c2037bfce120c64fa3e0a6d9135722b91453d380b305a6b28a984f93e15d828bc62fe4d44704290c825c99217aa5780a89e54fa6bc1d09993b811beb012f1f2c80400f163d3ca5ab15419b0eb765a1e5adc7fe9a90a94d6aab0cb32832eb91ba35223c8be1cb28171899eedea5657f0124318b839b1b745b4abdcebb033c746440a78f6af6cf4f690f35b3b6c5482e34f595de01836c99f3be2f17d3fa85c360e683eeafd9e1a3a493b3738f757b257b3056c9b1cb9f27970182451c079da556bcd2815ec10be00862c21bb0c78a03524b10b90cbdf626f6bd9f7ed66b15031e110825cca7925abcc01051912ef5da9f856c9b90d6571518ae5d2d9d3d519ff597d0f58749dda4bae4239c54b481f2f436e1c896514845e3e5907a677f6c692f76033850621bb40ae4fb90485be21677233d2cb30a38292b91af5b613047ef30153e784db7ff10c8fb30092793f541845581cd4f1210e2fbda520c4c64cb1e0b999e91d2cf9443bfcf652461f0e285a9051ece93635adee1c91eb1352e5437aa9dc5b5057d256d9054b84f8e7ed7fb329b80466c6478580991ebd54b537759541de4d191f273cb7c5950aa58328ec1c3a7ddd4296fe368c16a8963eccfed653d32fe92d85c7b338b521ad23a602a9be7b9f8a23900151ba0edced16ed5813e646bd9547cf0f19da395011cf6da6afc0ff17843a15c9732eb1a644560aa60de01fd43509b1c89b59edd2af9c52dfe3b0bfd90b1aaddab9eb1be312164ea46e69dea562f43deafa0f911be3d456d7de40f94911fc335b7ad8efa6b15bcfe921eb8012e3aab83c8a084b7417c65891047e9747ed3c49f90741e34a206e9752b6efc35a8fbe52504db003903bffa5fecc94c5e2846dccb01d64c7142ac006260aa72203b70af59ed53f75fd0f361664a16ee19b78d7bd4007b110e3ed536d6c72fc160f139118d62a36d082e3d98da1e95ce56c5df920b089390846e0602704e15c74ffa9d83ec3edbe94b13bf977344e9001fa550b3af22b685b9ca0e0f8660fb2cd017e9e84da0ca3ad995c5e0c0731be931063c52c7be8f2b109a9e55d5202d56e5ebd29638f9f3cf03ab8483cf7db63091f596a9d6fb64c60e7f0be4a39d17c261c246b7921c763e3fe16f7ad77f19dfaf27fc1278143c2c6d35eeee1d2fc39a483ec632e8afd094ba9280d9af6d0881698c8a71b34f862965d5c5c93c0b1e2b0689e121c7faf54138cb9acb0bac9754eed8fb105ab2ac508c083ed27e5054d9c77e79f26d9ddec339175355de07ab3256534b6d99cdc817a5dc0d4b9b0d7f526e7c085ac45d36ab31821e670117976ac28deea49ecb56fc3aabe48fe46b0bdc761189dc4d4767d4229fb1b6b86be01f6c45c9d2464bc37531934d22db3d5535f271d8aa27f8a3f391f88f320ac9650dd8e08e2597e51ab4e692bbe02a5997d920b38ce96d0e9eaf1b0739254f16f8c11828593812a4bac14cd5d6fa0f0d78b6a00cf9ef4953e4358c3327b2f2459773187bdafae91a37e7460f3bc7352538151d3c297a2d08f64aee6e40fdf885630bf7f9e677b3bc2a04949aa7973c0cefa49a173ab05f28694923a14840590bb3257cd19196ad01142caf9373147e616f251bde0b510e6511;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h7505649de55f14368da9e2a416145f821c27712de711c15b70d58ac807d156ebebcfe95faf03a1299a1d481329b5342e7badfe54d2081c6595bb0325e43109e677120252ddfee467e252770f9c83df7d2a755f3e89c2c2b75784e653938b731feeedb6d7a05b62e329e750ad1784bdbab9ca561080ac8938c6d05f0cae0d64a5e976484c3db66e86cd5667fe2c38de0e7c6db8824f3b2e9711b3dfe008a4a01e8f49745504ddf429083d13eea4e26a14b5c84e4bc445d0caf2cae63eb66a891eb599bc363e0c110ed4bd4496d07b3f8b1624dbaab2399eccd53d94f5cf588fb6f08f4dfbdee3263f5d2d61ac9e04cc74335d84209532578b345e3d2179abd620e0388fa999500b71cdf8339d4307deed986262c82ec1b8fb7b887c19ae0ccb72beba5d3dce24442478d0eafda5439985fdb97ec40b0ffd2812d6d21738f0758e1ff7e0bb6dbbc7da8a97c39a6c507537bdd00ac4793c6e7203e2de121d3912d9f7003f697a2ac5b6bfc65f33799f528a132e15e8596d49af56fd70311b303628cf5cf93ec12665ad589e478a46f6ecda449580314f06b4db751d482b20bc4565643fcf449f9d669baadc093e02d117746ca8be37bd796e371eabdd13a9a5a6d74cad8e6682d731370a9751b3f2b94f6bbd279efc0bc43d4d7668c8f9ec393ff67151abcb2918ac102a079473f517ead174e3e064c515fc9e75fa121effa464cf8ca44bc8ecf41f74a53f54148823e90e5391218d7511a30b1b28afbfd180bc6656db21b53ab6de4d8f414b65a2f5b2d17343de9106722e713b7f3a0ee0b324b5b462fa8d8c9ef7270eb4672e843d38348a0db2fff1f443fbb5964724366ad11b10ff42fe19a8a5014926468e39014eaf82ee7070cebd2b0ca2b31fa5b9244ae5a48783427fe85476edb487844fbcc061d31484afdd34456dc05aca610ab6c8c20509c1ffa4b6a3e5a3dfef347a2a88ee5a380a3335672c988ed59759de55e76d0b4950e706c40efe5b24f124077efc3333a85cc418138ca86b9617fd9deb980b6dbd61d1587e54927e526f2b16ec7cbe653c7220408cf0e534382644e09a56963cc558fd2fefe74a92190c0ba6b57de9b3e7131c077f5d73fc6ae784d5b16b75db2c890bf214d82fcd74a1bd15288220ce87b175ef1bb9e8eb3f9f36ab532d084ab4b917de231940f457c89cc49cfb6b50d20f5e27f3d4a1dcee74aef76fcbf498f3649bfacd239c3fadedb374ec9ad9b49e71a35648ade28ef0a261e92af736236fb5cd5c6e69acfb16f6321580eeca86e9774e52ca27bba00c8b7ba40ab927039da2ff6b9a56e287979806425e330001fc0421ec9d065c715e520e065cb7ef911d91423db206cb469af52e2f53bbef00062897e89671efd9898eba8409bac1cdb376330c22783df12283f2d8300db3f568ce5bce6763d0f1adddf86f2217028c06f877df5d03786ae8df42c3ddf93e9459b14bc1e14c07cdc05a3e2c4a21e86a679c65e2653d55d0e8eb5155d324807b8943393292ca9fa197a6ebb764e705c61f82de84d745066248860097e5f2b9c389766a92a67efe6dd7d7834c1de776e4b5f0084c6d1e886b8d359b4de9a28cabddcd39c42a6811316b5619c9bead260bd1ed828969b9c8f1c733b6f3ff1942799da4b9c20ab1fcedecd6da0140ab1df7f0db04ea5c624df1ac68ee0ed8c938022d59a8aa238d4a3f5ff0476999c0c3b539b5238f5ccbc3e3228797df7e1446d29654760c1b7cb34bafcd8144c8de08fcf12e66cea9c81e7ecefbd5520340f5eb4b6d88e19babe04836379969368b61b6cfaf479f2ff413ce36fb3b05b559ee3dc387c7b34ee26f6a5ba4bf604dc843f30f99ce670f0ca3640171903b96ff0507ac2b416edbc86f070db0c59f86bef6de5ea8ace19c183b981024ab1bc35facdbf6ec1c964070304e9e360c57c5bbc64e6ea5423cfd70db9eed0ae68f26a6bde775bed93343241b8a019300d6b911b8f4765309e62b0a218538906828e6c6d10701218d862740811fdf966ca6f8fcc2a5e702ff814afccbcef3bbb599cf12bd0f3cb35f3ee555c7b9ef6c9ecb3a1b6b0b4384b94dc40869e732818f2626a7ad24f9a53d03592d8a17e01ddce50f502f367dfe9b111ecabee6bd7b120aed0b1b4135461b2358457b54512fb724b9c58676e5b4dc277de1afe58be63d79e94ea0c0441abaa5fe56368df149f28a7b2a4190cf0ef72891fd671c62f99f6e6c7583b26d9559b822faaa3b22484d8c17981e0fac39b389980236680b594159cfbf301a3d394688294c21857f2d9b4a880322e0b16927e816764c4bf91f329183642db5c07b6b59c46d362a51a3c07bced04c51ff431f468576c214432f4697c914a2227038be00e65a2066d207ce125be264069db58eac7c587a4db10518c8c3b01dbe75219edfeca4af9f1e31f2f88550918556ca69e336e1490fee03ae04c7f8eb0d617cc880c800c306b09455b5dd9f6a1966e5f84d11a6c737c0d240d78a75fd7e993de24b9944910f1478aee69dab016fab56c010d03c9de3c07e125e238373a20816811b6b8551c2dd92b49ccaacd7a744a05cb2dca783b87e2a7ba2b321329f860497a61195e31d4a3027c66ad6173f9c32f21586e73d23180e7d2d0afcd40ae9c9b99594bdc8a9351e76c1716bc982cf485bf972b444000260b0468597a6f5d4f269d4baa411c1b6d9165c2b0d7f421f0c73db50bfbe308c12ff495fc052d996f8ffdb82df32;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h720330d025e0cc22c0852d6225bb03aaaa0853fc54657fced17b9d4f56f023e35996ad43683ef7a26bd902ede5dbcd9a510fe5ae59ac677a910678b6c35a1e4d21220047d29a25df7a0f1dad9fb8038dc84036f09a5ef0a646676e7cdac0bd63c1a6047ca2cabb47691760bf4cc100e7ec5f1c0b15b3fc3a4b319928436776c42ed50d7127dfdffe9092f2d3efdc2c07a7eaa9fe7a7391686dc90c3b051d14873ac5a33d9886b76b8447a98593f6d79bfed55917ec9838b592d07499e7c9b0eeca000d41eb23336344d4be87d659a243ac979a59249e19f041177894b2cb97607a78cffba3ef17fbac030b231cc73388c76f18f0cdebac07f1ad45f47c764ba0daf1af2f2f51c15f5e0c963a656351ac906a06eb57ed863babc194d1dd96bfeb2081e59d0e0060158c7bb843a37525af45b98331e6cbb9d2d5e397fd5971726772d761b51007d906b8113bd22105ff743ee90df1eb5d513014b4f492cbbdc4ff90a8606ffa2ca5d8cdce85dbad22171f13b7ac5476e755461990a32f0774c9ef0733a212413111bfed71e808439491ba248b0923b9e3c82c23b745e8d85c9b08968893e63eeb4cff3b511006565827740a6618e4aba2ab2340317869e449fa211f4ea2a9a83822d909473bee7a4038541d05443d26941c1db4e079abb2e9c243fe98b13938fa7686d1e584437d3bc4baade4450b10462b057d9f0c2760712cf6c47537c5814355147c9c778696cf16102f4a699a1b0d9c342bd8154267a865a9526c0950b32d5867ecc68ac8c0ac82a7eb2ffc30f5ebb1f35063daf7a3aadc3c07abdb0e900220b4d181b88b3dae7b9b43dd7f7dfcb6a60aba5e0d9889a419b2d1d2fe891b0557bbdcc3a1d24c2ad327c90205253076456f88518399905db92bf64f75880f6e3bb99bedce16200607a16f00f8e222c3541d11334642445460388cb5467099bebeb1d0e1ce540fcba4296d949db21a27ed7a06818466e3200638bcc056227523fba715ac10430c9d6a5bef5ebb29a5075830ae87826312c9dbb873756ec7b9d0174ea9000f89b28e223cae53f0e7f77c57af6264d8f46d8e2cace4790196f65338550de1cdc7a1d665ad3faf7b84e5d5aa4b969a3eb7bee604116c5d2d94aab98be939733b2a1f41c2048b56d20a2916a26163912fc160e467a53bdc019691b89160c6c5dd8943f9976a1ffcae4226ac21d912da2230c994e7e0d6630c19a53c4ef6edadb4e0bc3039fc28ea6e67ac5f40af9d806e6d9447992867b63f793a043f25136d14df3aa47ed186dc37d2e2c41adeaaef79d8ed8f2b683af9815191344606f57b142719771c8b979fddc13af198ad52ab2139ebca74455a79b2f81d5468afda2989d78aacf28f9916eaacf83667147a1fc9ba1c9d9971308c5316fb7fd373681d4860f4ffa1a8be527b4265e79d6ced6aee012ec90ed1a38902f72ae11a3ec26c41e8e1fb2a29d8e900cbc02164ee028e210caa6ec2439c38dc02b466907bd056a38959b21df426d68fcbe06b180f70462a96f885ed5928023dcb9e6a8daa42b39f07d40051eea29c1dce4ff9b4c0acaebb299e6a6499d8faf8017f26263bf69156c037f197a5092b4ce89f32d4e7716948986908cc72139581a608b45aab5725a35e8bfe321e0ee4d039fa4825d46271f3a4e0a59990ec111bd080ce82bf30d3950ec0934722a3848afede7cdf863530122f31cb7a2cb8e216fe98f1a5b97b33e4b5219dd9232924af976a71aafb1f0a668cecc183b4f24cc11be3870fc965f7bc5f8cc4136fd653e977fc9ff5fd1feda2147cc1b8cbd7c7dfa330d6b0647a247b00022c78299771cb2a294d8a3d7427c58d4851e9b42acc39d3d22a1daff30d4f848295cea1325f0c45a7e85db8b39c4b4c706c8dae733344dd0d89f0bbae67f5f85d0b88afaf4ded0cbd1a96164efb65f3e91e8071832246624eed8440342c40737aa88839431c1c9adb436386d723b17581c459a9e197d024203a01b91105f6636d6f5f196a7f5665a071c2164184ce782f34731f08cdf5b3b8241cd2f81b541e77e3b53b10bb1c0c604fdec60df0d745aa21f635cec866a09952c9ac524aeac7fe87f79a978d0aa05ad5469bebbc6efbd1fdce516dc7a141b10454975c8ad9e30c7fae1967c2d714284d90e679fe71441f4ab0744583585abf4b3391c39c9f1dd3094c7170f5ac8f78edcd77e2d7c38568b7293daf22481943ad3c02da01602e470a5f020bf28cfc9cc8a9baa41ef253160e1458fe41619536f8fe1cf0343a190e0d99ff2111908897212ebd4af9adbf60caf89f02c9d393998fee9ed30a0dfa768b14a3ab84c1a32132df79e3516a626711ce5972d2f87c6ca56f89ebb4daa4ec7be7df50c52a449357595a99a9b82b90f78888b246483608bfe341050b608fcd761d6d7f32c12238f5cad72c402f07eb3a70c16a179fb9289c2b843dadd2afadd91a491f281285a3f4e47fe20ed1210ec1f12c45763788f50dc3eddb853d24e9515ea6ca4edfed7dfd23bc03385a63042505fe15cf3a2768f6efa6e249a059b320250d50838a8acb53cafce12e11a66941b957ef36c613a4b190a63103d156a71bdcdd0b81d664e3e1c7b2064088bf0839fbed83d3db446e2e1c2a7a1d34c1fefb8c5d25da045f22fb5d96baff7b6bf812cf7d15b6efc037226317384105146114af1f1b5bd92e0fb3194e27f2d60cc5ff0b3d6a48b072adadb850a47ba888cfbd6f6974de724b5c6177d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'habde9efde3d5feb9aa2a709cf82348385324d56aca3d983a4d4ae0428e1069082e17fc29c23e0f8b5972b8bea279fded50cbb52e8526f86448f2e183d81121b5f4b8666235aac43ce2974b43685b1e74fd3325bb8d7d4ad6ab4f80a94134b81618111ade3a7bc3c447f779d56b25c0c615817b4c38aade66eaf261d447a41ed5099ec7aaac910417a349f1e93a7c90afdbab12fe1746fe29a0b117fb55e443af52199e31f7c0ab3395133d65f147e6a3be282e869f07a08d91c36fe1cf4443ef428411d0c6c3e26331b3552ceaf1a9a674c2969189eeb3c9934d465ff6f1c2fe7a78e548bcc57a24578082cf2af4e9cedd2044ba18f0c6f8e251571291a75b043b6289f5651d6c56c5e2589d7001cc280767e6304bd7789490c7047a409a1a4911da9d98ad4e22c06371e60db32e02baae78c0f117a98b75730289f18686dd5121ffae8cd762ad722f3de1cf6923c2d8c771d1241044b221e8580abf6955ef76a92afa84e3ddbc99f8a8fd522285d3661c5a1b3f41f702d20f78abb7617d68a7d0c3076ca37608bb16398f578b49d8df73a9e822cfa44b6296da83db7779a6db376ef0a67e7aa85ab1d25597d01a325cf00b1d7937fe16cef45dd4171cc86bb92e48c512fc3adb45abbc0a79fef1983388550e52e740c7438a7f1adbcbcdda0f40520e8173241eb2743eeef76eb92234b61c2c8e84879decd9bf954a7794f3bddb637de811428d6acd2e57e1e759cc6739fc6f254851e3eea31a400d14b174c2c81520908cfb234ac7e0abb8bdc3c2dae065a875cb34007893b748fdb1ab8f1d43f74715ddad0476b924bdb04bb80e26323061a5abdcda03049f575cb6b028ec111485eb120c13a6c5f23014483391e54d26f6912d2684bc2837256ddb4ea21ca3457017099300c9a59246d099b05503f42f625e3db15ebf6e77640c8cbfb46f3c47d9349b180eb4b3d96fc541e94a85981d2dccefc6ae174adb0606f361f62f9e82ed1b843e506088576737ac282c2f9d053edd6bf73c0caadaf31406f53a97ee3031e2d663786c39cb033a3b0a05c7f03b29ba92ad91d5c081e18647b6c4e7b7663f6cf5168c8c9e217f0e3d64e6a3be182bd407fa2196eca47546185fc1e3114b1862db23e920695036af240dfc3fc4fb77904613689c9de372f52f724a0f73e2320da6e3ed7c18c92da60112e0bc85e395a6e45a18324de9ad1d0e71e4772d441e749d6f7bedbc5ba6248db144b9066037db74c06cfc95422910384c0bfe5409df0087b35bc1adb8d9cbb95f48fa59b4eb047b091a9bb803b0ed05035c5d76970e3dfda738c7ac239c2b506619abfcec3cdaa185b364afe03fa50bd36294a7b2efc17781d20eb7e946d5fe5fff4c3ba84fbe7ca7eab1984da5b91aa38b2d290bde401d013a365777c2e695b155b64fc9deeb46eb25559843fce28fb7545818c6b81804fbd246f3d8d0c3cb7e79783c5040e89b3d9ba737a22eefee5345bf886aef7d9917c1f56089cf8a844c29650f3742f0c24012987a742ce42133ca87b662e69f34078b975451849b0200076837fcc06cfe6bbbbdae7dc2b1f5d77dcf22867d80378f56ec0e370d3871cb56609878f225f605b61bee5aa482e0bbaeb6670fc41759e3f366cb218b31a2a7c9797f787f8c1f63451f30e6f37f18363f22606026f1f79fca9521217f9b0fde98ab376f99e0bd35ee3dbc8fe32ed8ccfd989147ce4df3bc72eac64bea878bf8f9c1dbaf63bc03dcb68b9313052311104b97f07873b36515c4edf98dbc61a39f615dd559c635a58bc89aa693ae20838a52b1f82dd57eb24f7aa878b6931c44cbc391b96ea62fef556187a2aef8795b5d6b5e2ce985412f644f11a467caa96bc9e465947ae92c7b8e69ba58b73876f9355398f08bc99ba2e34bc140aa085a8d90d1ddf7bacb017f104f088cc4281a31bed3ceb5e7db8a2b34dc2ae7495bcc1b4e5b56136e956dfac2d70334984027a0b5de1a42d23417054a1eb3afc37ee72316ee2df304f190d5375a52ba305521e41e08e795e0bbc25f15ddf32fafe0176858563d2d5795f9b696d6511d28f6475899fb286abfc5e3fd6867cad2630ebe6f6545c9573685961170f237e8ace3713336dc589ae31d5528209c9cd2821f91df950b6142ebc95bfac37c2cf308c765eb527cd9217e6d39255d78e7a885bf23b734dd4dae38817ead7082e1fe254217cba4b1a5aa45550b4ebe480cdd0a9cf053ae7f416153ac3ab3747eb4a34d06ef604ed0ffb5547ab0c10464fb81aa4a109016f55258e3c1270da6fde242da9c180fceeb08b79d274943daabfbc0dbe6aa9928d97f68d4b56387861385e44ce41ab96bbf59dc96fbd86515596e14822977e74d0f7df451ff146211add1905a529cd3343e9069fbf7fdfa4c9f41063ade3769ef1582f3e70e8689c25ff8722d0d81bba0213006f4f02f5b3fcdf05e62ed5af833194cdc79e6a5f922b73e0de80c3f8fe27404de9f6d69ea88a420804aab77636b81bda1aaa851731635af14610fef83eaef1e0b79de424d766dadba130ca65a73f122e8f90ec559e5e6850c5945fd30e35f10c7286ae5b5b449e1ea2fe6fa63d5378552954cfd082d76d30f75eba783c8b620160b74868317b07844033578d2a685955f30b8a44e1c19deb3b8235d877a883480292dcc91cb91280d378ff539d419b79c7ff2c2a9abd2a786694045b58c2f3fc29139d10c2124e3a0e1551ca22ab2fd35b041bab3d543bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hdbb40d9c03339ee894562787a40294049559891f9d39ee5cfad15483e29ca62dac64da8e73a3fe553b7dcd3e667cdc8aeeb98c82a6eee67f231411eacc5bb44e222220f7e71ed56977c62199e85bf7d4c9fa1dac149fbdf6e0eb0d4f8ef21136cb5f7d28d9ecf8ff8cb61280d317c0bd03e9ffebb8f756a69d3f978aa00564e8b43ea30680545f11c9c72810d80046b7a6e3d7db901a712d379dd29e4539e611f06102622dcae6afe8c490a14ac1b95709fd567f14be52957ad7ff0f052ae9ae2a6ec60e5abc417b918f3ba3351ac1efb621b338094b31ed29be6a60b3fa8f6ade6afc45509534125da22d52c7519f0d1ee0fb70b64c38c38dc1c9a2044c325401d656ed23abfe2c98838823102ca2abea065d8ac49d24bfcce97652b1072a5e352b9206f81e168643ed6fc929f928c10a3f616ca8b73b1d3409d635dc35eb5bdc2644df4bfdfc88cbd6f043920103d139787d1ed4a7e969104755b20a14776721e459aceea507dddaf7d6c44cca85beb072fd4642f0443c8e892616fdee494b25238518431cc59199ce6e5fb5741315927807a6060ab32b5634859c4ea4c0a73d8b8f8c337cd1bb8a7e137e6e385aeb0f1fa1203d5758dcfe49433ce64214363569604afc9ae540b4ec0aa316c0867242b58b9611254bb588445ba4f95d0ff65ef13079e9cb99a26dfe03afe81c50e9afa477bb2f56a222f14bd21d2f25c12366b4642d49d684e76ba2a91bfceb9fe3ccf7dbb7970405e079491a6c1bdec51810c140304d44c666cbe87b1eacf2ec1ffe9ce4fd8e24526a99823f965cd96d01229fe81276f4910b685a3e3857e150b01a2ea0390060ac4d4c66ce5eeccf97e5171668e2b95e4b47e9160d5d5d72733cb8368a0834c7cd629f459301f6f1a5f8998e4046be6e5e2d697aacbe4971c5f6e377e994ff1e5ce6b530e4bd10f164b0cb091697b60d0e41bf38ba3819d4132b9529a23ca70bc15d4e9182d68851579a0e85100b3e7a5d64ab3a62542f0b9db1dcd7fccec87715793cb987d0ea322e7bef7efbacee573cddeb6df3e34af3ed6945cdd6654598f5433eb657352c6bd579733e132ae04a9067329d25ea6178ce6c5a1b02ddb697dd09d6d05c10253e2edf5ff28df2dbef72a1beec06e5af896965e25dc137198d816f7bbec2fb5bda72af0a1866daf5c994ec9aac2006672175d1c7fb8beb8cf63522e9a5676d2fb0877e2c8e5c5440e6ab295f8609740903fcfd950292f333b162d8dfefde8064baec7bb58102fe56cdcfef12607e8e2e9bbcdde154ee02288c55917eb6e9b583d588c3a78ef4ebd70338b66223ff3035372f2e09ffc94559ebc0275f9aec978da3ca90e60db33dc3086b59fb0beb3a626eccfaf39667d05428a49f37ca59843372f0ab0414762768e535b55503a9243a0109d5ca84743337d86681d0195540c77114278a53a62656b25ee1cffae4b76fbc57b4f4019ff4366fdaa3608bd82a2b10f4cb8a2844d2924c5db261de1793456193f6a78b500135a898a2825b34eaf648805c1a7e0b54a6ef1919bf121235e9aa3f01b6b574caf3e0f59c8b0c8aa8c0169c26a4709d9c172031dd66d99027fceb25b698960eb651d1a38d523a67630da0e9091aa6ce84a0d8dc13b3ee81461cf5d3bda2b8499c2c4dafad3a1f1fb91992ebb825953138cb36496a62ddbfc80975972bf7e6c61a5c294dbb1663be128913ae485c8c8ac8bb11c64952c2b69abb9d3ee32f3ab32b621d5228b6e4ec42681042a51dee92dd4364575ac08ccb3ea605489c31f7a45f423280e73643f4432d8adccc8cff149ab4942bee4be0af06944391c575a9f72259b8385a432e91933bb1a12db4fb335598d1894bb34282a7c36c2f2aa2f76bae4356282af35c5c562adeddfad1172849d63fe0742407766c311c8bd66fcad7e63dbbafaba7ebf39cbfe8e3448f263acba5345448913be375f5b7b8b5b895ed0065aa8fa97d5819ab3734de28bf7dd5d5bcd464706e5993e071f5abc7d24ee8904271f5f2608aa140c17ec04295b3c100d66714dbc29702ef5484802b7a05f834b81e3bad2c55628bd13ccd1ca1e8b24ae7cf9d12f6decb5d30c36b1c98f866cfc5714a21eadade77d376d4b2cc3c3e1748ecc5f671918ab74e16e548c4cd3665841f43ea913a118fb9417bb55d10b2fd21c592829339c9dd6d947a74305dda989d9e7eaeb131e3486c342c9998b8f9b778d4108209c54fe88815f65e59d833f68525e93c82d0e0fc7dac923f8c5f58ffb5f9753f9130f7a206827c9ce9f2ee52d49cbc3c5922486690136e8e87a15f39a5fed60a07accdbc254741d877bc9d7ab380cf0044d9da3b47dd8fdbba647315dab2e79478ff3ed801a32139ebd080e5dd2283dd8fc30f4913d87a34874b4bdbbd5de51ec10421320e232f1aeb1ab360ada8c745e65d0e0cda51ad83d3b37fcff011580cdb00a040f9a068c42d02d06d5ec270db1a3505166f9184aa8c490d1440eb0bfeda18b9863d9897c92de1e7d868a2cbf6649f79a796a680f2a6ed95c014534db05b925608c3b8a9e497afc265e630cb64246a65fdc8f3d77495487a1a379c37702b75c0a515f5b39a400ec074d6d9469d469b98cdd407579f9033b1a4ee2d2d9e55ad91990bdf4cff7d92fffcfbdc92d7979f4ec4e979d5dbbee41a629b8a93ce475aefe74beddba30767fa8da2211eed54049f5d0e8e2c49cd6f41b2026cba928e8a16ff1c808d96a988d1771aa9e8ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h7550d9e0283c333625bedbb8ea8bf073a74c8b18dfbd20234c63e5121454690d73f3582aa5b65e2257a6b8f3ea3bb2846904d0ec961d2205343a3fd896f3e0a73139b70fa507afa4aa95750d26030f25bae6e9ad8041b4f9d4ba2135a00657de4d5c245bd7a9c057d893cea8f480b57bd3543f19a7d77f816de0e91ffb87fad81cc01d569f0ceee7e9bfb0c5cf1eb6d81264bee7fe4b39b084bc6251beab369272345a1002d6d3c66705f60221c9bc94f225f4c2d7b0720ff77123d4c669a5855689da71f5bc52128e5693be23d0181e3a5cdc92afebc86361899d17784a08a64318403173e95dc2dfbb2c4ed9fdd3d9fcf129a709bf23f44f71721cdd7a9a6deea4ff34446df0ea4c97e50e393e1daea4c3a0e597583d52fe5dd13c76b16365e89f52cdb752fef4a346526ff02253eec5ca49f05285dd958285ee6cd708b5da62247a744d35b1b4d932fdc981bc4343ae5c14575a224ca110a20bd2e5ce071c63654bf53b2601e478c6192730235c22d4cc0296c6cebf007abb7367f0c92522a6242b38a3013cd254b629292586aab275f1f06be4023237cb1ea0872ea72bfe9fb9da50b1690503f3a4909e8f95668167b2bd0c1e0b46dadc08561ee0527373761566718b69fd4e421fb7e77b7b0ba683e6e6493e112aa69b0489b3e3ddce2f375b95675f9bcbb54251342df2a189b2060c6f5e0b77e07647a47a2a3be9079cb8e0e15365afdf86cbbf10e19afb585a1f6952b2d54a8f469d6f65cca409008a6206ac9cfe0f0417c73862f61ee9e19ce659fec9fc2b09f1cb216b8ba6f8fa28014b52080ae8aa1fb112464a0b840c0f136f43a02cc62bd947dc43f6ff676fe3800d047c7e759062a7ce7ddbda6d2b2708808e93deef38aabdc73fb3816a171df54843d1f9891f6d9223db5614079d628a7f648005929131213e4cd7a39bcbfe9b6cc455b6ec34426370d4111e3104e9e3f7553d2d1c0e64e2d90145c6332f587dab717e03439a0966f474bc9589dedeefc4e78cf2e5f2414b00323a006d24baa6b7877d78b017e52abae3c8da2159460824a397c8eedfc90fadb845c094c89a3d23df7f66a8b0656a4deb2477e57dbd0825cca183ee93c9b5d1a5afa5ffeb8a6e7a48a41e172adbc90a76aab570e469e89f66c2f72641342eeb2f64051c7ac320726ac0b1ea8dc88e0185b70ef072660650e3b00776e646cc167a82bb62eb5c40107d537d127f517e23afe454d660182c6c92ff4049dfa05b37e5b908415d52bde06939980a0612456c270da2d922bd370a764f8303773620f74a47799e7e108a5d3049bffc0a1f26c202ab65bbd1b23c2b5107b111e97e91d52fc26186603289fa1584ca38c93ee1ae01f1ca64bb45428ddcde096c92c71434818298d787c9a391f02ee0f618916c9d6aadb25e95157c95822646dbee741f4020be75a283701bb9f543b46dc14b8da4fe709ce178947f7ce08634cb6369aa2ae6c4dc383f0df279b3870e6e1093f8b967a39180a0ceae0768a03dc9ef2e0ca847410edff541a0a4b8a8685da52ed383be2635ffe73badb77ea972aeed96aaf58ed1d6b0994dafbeb894546dbd88f5dcd4dcf1938fd12d5af732eb10db1d6c98db97e34c172f2558a83bc72863e3edf986f38862ca3bf253f632c52d45726fe334d38c71b59bac836d095cdddeee09f6a32b9d6d2625c3ba2892840424ef8cce9cabb40d27a23d64757623dc672dc1af91606a0399c372f635c7904af8b93da16041f14c848741351c2d5c38cc6831a1f562eccb61221cb481e0d22bffcfc711010686636cb2c8a6310824cbfd3ffeb650c42056487aa5025c213ded03283d4135812ae1269052e43bdaf2318a36f984ab69df014765ae9e7663e464d8eded106b7e3e24b0d8afcdc769c789967bf3dd0f8010a7acdc05d918f238853ba0e23b450e5966dc5cb50d66c9ce524d1771799252117229de1d5c02f1821eada0920c97165d8e1126bb6dba5f81a1c594a9a0473d2ec9f2ea2cffa10ff0caa9f8e5993ba5a510afc8dd1885639479871f46717935fdd64bc78040aa7f334dcb89565262551fb1de00d756bee5f5c6de48d20497fd3bc073448df921f41c14180c3d5fbda5c3b6aea07c6716b6cb2ef952d3564787e20e8672957b6e3342c3c46bafaa4146bf4f730441e94e8bb4c4c9e83f2573140bebfc29a276c68cdbfea599f837f307d172135c5cb37c2dfccbdc6d33eacaaf75fd9e70d30263385793bc5083e9c64bb26016d7491da41df41cb9d0371698de0eccad6c76540ed7817e9746d9d191edc4b33f79b504b93cd8858916924674e358aa7505115c901eaa6133893527a8d09889642906c93b490972ad49f650aa71214120e5b745e2daa2020f1275a4496091dc80f22f2452ba9fd5c6dfa2658d327be1e508fb87bb6c378c7b51b2ffba3ef126855bb9bccf3425728f631fc2842faa9f26a5a26257056aa55d5560e78b3ff0901f4f2ad6183ddae83602f945a775f8b1d0683ebd3ed20ea316db7b466cacc7d5dd193bf04f0c1b134b05a5069f28289784dd5bf8c3efd641cdbb813f66a9b1ffd96e50e2d1572f720eda3633ec77c5b101b05a22cbb87216dbb5d662892724dd2bb9190bcb1cbecbafb6eb0e37c70a8e6452c096ca61b19893c59716edafbde681fc4d4df1fda30c5b46b56cf0037ea7216f69ba093a39d409dd77d5a7ce4421b5d1dbed248802eb60110043204de29235f10945c530101bad91;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h400ba77954a3f1fae084547ea34a8c084290472f2d5b3435ab02fec8b819b3cec8064d1da8291d94e3668a8f62674278164c7ba6260273352f042d16753833368ad15935bbd3cd5e8e52cfb574b804dcfc480be7a06e44dfdaf8ff544cb3121e6750662c704796f51bd7218055dc4a2711e0a814026a8fac49857565569c6ae2d5ba4952bfba395313c9f3375b5fc3ea24b929f80ce7d1476cfc9b613325bbadcba07b1c4021019a3e5ac49c8c165c0445a7ad3e5dcf71dcda4b7affbfd3b38bf83d95625f425718a58f6a7d03f90fbdc74883fd91c2bde9fd55f868ac865c178b6ad48d7683a8ce30273be64ea240428ae0e3fcbc04b4e4e87cd19a1bf892b62798293a87d9ae70e083fca9cedf7bc7a197024146f28c916f8fd4f170a2c2f2d02d7a95ad932b2e14d4f6636c14e5e177c0b871a6062aca859ffa9256c88dea06dae5a949ce2d141c1e8a7cf792da672f14e1abb67dfd726f617f126657d5fce36fc67388496825e558a210d5f311eae707eb60ea92347ab660f2bde0292d45db5b5f2db45a74aa53fa6e93533360166fbf368f03da41584c8ed7f7b7c35979d54b03deaceaeb632162616df91a09a39c33c596fd8ef2787469ef2b1ffb5e61212afa5402be07ae175ec1f6085b040fe890316532cedca2ba4e8618c3f6042cddd5ca6612ef2e4f078f404019d7a0d99ce902b97c64f3faeab9d3fc7cd33e10fe541c02b2c3ec4a7236c017afc20a3d04c21d7574a07aaef88ed95aa29e47195e7d6e96eea18b0024554da77d547c1bc38ce05291975a037ba122cbfdb50071f510c88b328086e86e1f846b091e054dfa30723a555ba592495bd87c3691f87a24f25bb44da07db27aa6fb78db0c7e164ead7d3c936026d59311328cc9ab41a62c6f0ec74c26f91e9f43ee9710f6d0abfc83669a11262e0cb5f135b3ff8df8e30ffa1b1730aee8c96ab981bb3f263eef5a789b5e65fdbc3044d7349faad6dd33afd1aad0bc6c055121b1f68c3f779480b28c8003b5f4d50bbd6bd02e487edafb60195e567f3dddb7cf8a77f62fff97d354dd1ae8131ca20be2a9f36d8820884461ff3a16059e3de3be0af1bf6bed77f0e29e70587f0e06ba671fd6d0fb81ae710672e345c91ef52a647ca739512f80a895437673c2c9e9f0402a32b8a6190f78a6c0962236e60ac78d8c40f41147f5d10827d36d5d18c3d72ed61fc79ec64bb72df007f95a6fafa60eeb2a9fca34fe74851471622812e9d340444e080027df0695c5a641ae9e84e56ac69552c32a2db6d11b285e360c04409ad8adb698d9e7d202aab87435d0051d9d28b6c9b9e83982e05652995da344f0fcde5b21b5378c05b2d17e758dea0cedb6c0721c721d1db029ae73fea5b2321046263eec93d98fd381187a034be363f3bcdf4466c08670581d45a9bb7601b09ad7259e68141a2fa5f2891bb7e3218cc93ae5c470864d0d680de24579fe6abf79c0c9c8b45f7724a245a67c0ffcf67f5a098b0f6cd6751b2a0906caff9fb56f6e2adde56843f52a9d872c4951d42080d18852f13239f8467ba5afe84efbbe858b8a8aeb86839872cf7dec59d285d8521cfd04eca17981f8a58d034640c2c3670dced6143449f01c6c3a805515bcda141ea805973a8feeb373558a8c82773116788bdfb614a5fc6120c0415b4a790776bc9a07a49993b96e1e1fb23bff213ed08bda008409c04e38c9a1f6c97279f875c13ff09466559db213d35dcbb3e2ae74e63578b90b6dae11bedb80b81db14fec23cd2d00037197f1ad48c84c0d6a345a29ec526f0eaaae51c53f690236d45882c731b4c1909400f0148e9c10eb8cdaed5f2969afeee5219a6eae26c43aa40b25cd17ce7993f44a6ce360f0c9bdae433ae809a8d128625221703f25af9c6a3aab383305f8a0baa000537c7c2148b3e7e5d48331cfdd74a8b82a5efe9d86bc3018f9031eaa53bf106241c8e7fae5b07b67719d1392773ae6f59f98589c515bc85d4e119d01824dc146623feb53cd10cee0664acc8de0dede376b51e643989d0d0f86b434844859272740d926e074904f944265109e28c469ef00aef2954d066523c53b78aabb74a408d254f04ffd69abb9930b5291446f2e304fc3cfa49b7903b8725e9f5dcec76f4aa503abba2d24517343ea48fbdf1ed070b9976564c1a4ad157f734570d7d7316e0d5b5e4c6c52ca0d971e92db44af4eb61e97caa189269fffed0f3e9c96669cc0d0eeb949681a09f89bdc40621e52c5d14c3f02cc1ae40dc37deaf07119bfdee5aad394ffd5bd8cb8cfca8400f4e0dfc6b127426544f20cbe5fed9d1d965d4ded9ae4f1200243531b34751d989c884bba746f23daa4fd277da6835a148ec040a8419945384120e8dc834c5ccf0ed97a2143f8312a8f02cbeb3884ad9a52b245c9ccd7de651668cf406eb364a449c80b59aa65a31aaa9c95db57749eaad29b2c5c1c8e3d1b70e7139c55ce93612c67f0a3cb38e4f5fb18d50ecdc507ba6cf157db92852dc2c1693470827f6e7b8e49cd9b4c39a7d7db28e8c582fd29574a8fef05d0be9a71a4d7c40606a22d232ef1df89d1bd4144f7b9d61b9cff0a6bd01da7b62fe7972c50940fb83ee5b0a807e1d2f33df4b3017063a59906df5fe8f9ef09a414777cc68d0428e6c62d0b9c04b1075c6be798097e9d5814659689352c3cdae64b7d0add2c98ed330d52a5bf79384726fa5a887ec26053c0f9beb483c7655aeb83b8a11e462bb5964e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h5a68bade2cf2be7837cc72051f85b3c24f7e891ea6bd9c8fc300327e97e52e40fa571159b781c1baade4042bee115a121e1bc3a905caa9765fe9de6405d36959db482bdf8f42b5ad470896610124328b3f0e051489953c95441fc72ba82346680dbcfd6c6a6ceaf4e90ed3638619b9ba694e6a55b2469b9f45e63c8db47eabf277f7b54b70d83e9039402230fb1795610add61ab1381d70a58b2a59216014cc49679fe3b45d5eace7c47d14e94ff8d386507e47a3e9eeb36d6efd012a11c2a03cd44a662e302c1cb4d3fa66188a249c24a874e68bb0e044cf7295bfbf26b1df835c7316ca4f5cfe63d13aed09c77dd5d9e66febd3194e30b2fe30d712e63bf6d9b451ff596617669d5ece49eb7589dd39e7e45dd07f38e784d1b94d9b0d0a91bde6a6633dabb3ad027e7085bf005e3bbcb97ed5dd304f812fd0da0a929c04ebad4b312878c2f4ea510cc3319edff6059674463b55740f045b705ceb6fa1e28534a02815748b1d315d9bbc45cadba4dc654be0cbc7c89030e032b5338e3e2a3ab0e573986de6fb4faece2d16d2399bbe13944cbbf447d78b3afccb3f339d16a7325e7324a402152d5bb3f995747391c66e21b002ff792c63e709dc0a2f9eda59b20e2d47d05a2e2d17845a3e3b554e116e7298a44503bf7a9db982caf76da7dc65d37fc9c4a4651b13260a876a8dfc1470e43b952c8cbe267de5ac6220fdd108b44fec2d4bf09d91aa45b2bb75cceaf0496f0489dea41311698388411463c6572fc7cac7e356ee70ec60da5203fd4bdc4af6f56b1cd92bd1195bcffc6a20d7dd63cbf31d4b721243373dfbc6218400c79b602f77357ed21a6bfc0e05f38c7600a13a2a5a2e4dde6191da4948cc29da32371c74481e96e9fe49fcb9762810968ce7a64239c5bcd2762303b28116d87043f33500d9c29dee668c4aa5100ac4e318f0c26ffb34e85a8fdb71d66ac0d0e0c1bc9b0fc1b0569f42ef31d212ac2276199999ff2ab52ebcc17d8b55d05afa53e58bc39c351c1fe01ac97430a2022c9edd9f76b6c12b0e6bf9759ff5a5234460a9e07472302961e6928fd3e36b008b3aac8a8934bd6669327f06f1f6ca7ea6bf0bd247db07e13560c70c377a8fb86c8e7906cb7251b6586b6de046057cdd578c48e069716cef7affe1eec2c013dc10f646dcd783bc0326f7e86ccb65305165fae39022a402d82081c952763afd1e4130d64fff26642f74e0317541300b1e79ca00075626c8087fc43034844e7a1ea73944c8a6999acb08fc2e47fd9004a5351cef729c78d012269665614ae3c53ee04d61c93867bc9ba62ec7b3832523833230548c0af59a842d69b190fdcfba44b05a2c9336020ebace4dcaa5178dc0b040b9133ee27f511c9f70a2264ea3f69a8260515c25ec07f8a3d58991e9d6bbe95f06771fdcc7b7314b017a6b09d49a1d58bf7d4342321adcf4ac458ffb753cd0f5329060e9251142cfd418d138a21e191a7e35a38c2a5de9b1623a077ddb1d8f52c9b5c3d44659a6f489bffa59d745ddbbe1ea616e9169124270be1926c9eb9f8f587c87d22a1df8a92ca723140b22d45be0566d735e3620d2b5a5a06606254de4416e943ee41cd7b739abff04dd6a14835d7ee971a8d9f84ca71cc8abf51a456c87b672afa61e91b87a2e47e0132aa5b026f68c2f4aae61f4b1ee4b428d6fac4e63df6bf95cef5aa330474100801d2c3a56cb4c275f1acc65d16052e350651630ce0720cf1fcbe4b5997e7a2927b1b168a70699e56557ac1f717176ab1680a1248448c9b059009b9882fe3a2d4956d50e535c028109c1302b619657ce2e20ce7db58cd3ffaf4ebde4096676f5a5b30653b4f37d9246b60801dba7bb8712a3823f9bf02f8a4d0aec31ebc01d7e9bbd442922911efaf95f597a1f67059265ca89abade9b3d60a62bde31e85827fffd7a11a0e72bfde31be58b02de68d28eaca7bd3ac360f206bddad09d3d73561fe96651a03b3a46b04ed4d080ca04408023fd8679dfa4927ad9635371eede38ef828949e350b97a28f416b8302b6d04effc74880356b0e22644488ff2c35559760a6ce16ca793a6ea707ddad5cf444db344fc7221e0e6364dddcf275299f4f926913185c8abdae25f31e6b1c5389d82918647415d150434ce37fb7fc16525c3d20af6e9139b4cc591d9cf23189019816402ccea9a88ef8d3dfc03a0430cb22edb1f2ea9ddced16f02d78737fa39226e19d7412d638a9ccd8a676c235e22feb6ef70977bfe6056091f3950aace1fb054d19cfc1afaf8c1729c51c1dec2e1cdd9e499033849a8f0e462e4fe25255cc7c7a6dd24d0098a5ceb4d44c96745995fa594ed55185367444ff08176dc93782275f6949fe375a5a364115c94f1b309d33ddd5ee3beaa897a4403d5eb3b1fb7a46ce4f174382ae119e548724045255b0b29fd42d5eb11546f6fffef9787adb43b76de5ba2860af40a99c36655470dd023145dd6c9b77501f66662355073cff0d01cef3ca8d45d0eac9f04dcdc28f5e03bff55abc58aea2a4751be9e14f24e24dec3e9b36d5e2d2177eb83e5275f5592d2fef5a09b1355c9bddb110bce322d974a2d0e8410a612ae3262ea1604d03214eec7fb69cd56fd7ae4f8951ef45d000bb22e772cbcb75b8f0bbd6e3608acab9eba14f7c9b73ba018c4fcc449941096956965130e23d0d905c22f019667079d5072eab38b9123d2f9d4005bb53eb36e801204c542c6079feba8d761af008c227d17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6a27bb4d46d9801d8e5a09baa30dfb840d2ac1e1ed468619b71b97a64c8ab22d02fefaa3902911fdfb5bb6b1fbd0381e01676856cf890efd6fe110d394180bce9259b3961a0a0acebc0fb99c0b51e1e1819a27914d99013684b57ec569a3408ac2c387efc9b92660f564a3a01cd4b6462281b5cda7c8dc5e91f23354de924f7aa33ad473348269dde853c6781670687925bc8473fc7107ac668a8876ee73ff49903554f3b6420d5a35c30dad9b4bb0fe442b1ac25dd53da98d1cbc0ce575c9ded62f3838064010e22ea6cee8d62e6fb676e992bb554f554e36d607d2f2d8483b5090de33d2639257ed6441c6c2fd3cb3d45f7e46be9fff722d2a4bf3adcec97bfe5d3d8906c85fbe4b6c3eeedeff84c82ee743794281be29f9044b7a67aab9d99c9250fc19773e94e35fa4714d37b55bc5bd820f7960128780765837b1a5a2b0487822ff8875c9dd3e01c52664c6d4c3c6c136eba0da7b4fd4b54c5fad43085b710a0a3018620981ccf976245d17c76ccd3c4784cd8ccebd4a7654649711445cfe6c2877e8eb44fbfb75e8f8d6b668b6647a70614c2877497104b3d8f8c83fd3fa40f75ffcf4c78f3573059bd3afd9e9fd405aa0608e23112134a8d747cf00fa24ec13a05fefd977fd5ac7bff8c84378b11f1d67a30fee2e680508eeaee0dbfcf4a4a69594f01ac037d9223b2e985612b197cf4b4aec31ee0dfb4421e53fd7467d1860019f41a90d24d33c85230cb8fa2cfd4875bd330314db0b145c8ccef0f60ba28d3d60aed33d972f80df92fd3a34108ef30f6e1cbb7d43a58f33b50555df9863a68c8ea7053396ed1f6654242ea06f15beca4a04106f5bd0c5311d1754d124b896b528f5aa8a1bfe66015b2dba5d2146c2a09a2121c6e2b4e3af9a55dbaa17bf3bf1504d6181d9d4566d8eb5c96b89caba3d09a9858f8b029104712df055fd497f5d2b29e07b3f1e43ff3f2950573ff3de27fab93bb0228108d2ebedb99547a5758804fef00d6a78945333f06210d2468094136aa64ebb8bdca66b228c636c36fe3566d9b3be08a077d608643e034ace87b578940f0c14c24bb1e1edd3cc2b33f60f8207bba2d8ef9845b1e7f26a35fdad9bcfe5d5742cc879745cbc9dfbc99e445a47680ed7674a23dd367e1ddf75c8ac6f8e959427748fa7a5633b2d78f48e48816ff182a63fd13c2c1eaf96366fccb9e9b2c51584e96af6c8026bceb241e3c75e4c845d39b5796f6145eaa8e1c59bf67018e35b6ac8f14af2f0972a39f2a7e0be73be0050e19aef33672e2632341b36c07fb7779561db46e6950eff8847d758afb494ad971829855ed31b51a8401781bada392e54690d34692f57a7079fbbe8b5434ab84f5cd7d4c0e8592b980aef40fb64c2666ac93ac0ade034e9923619b87606b7525a50ceeb157dfe3fb5cede6f24b8884fbc3254a0b59f7fa3fbe3c69859b324a4c3058b3a1174251f0451a007ad3dc23f746f8f7a014c1915fe1b42161b1fac6a63f0078ccc1245e85cc66bd0637f9f33e1c11302a55062c3fcef5d82eba74a243cd0411a5cca9a9d9746f3c068270104ae553a600e8277c032364c7624d4f1d264f0c7d6577408a3131296a9ebd1577a7e758980c69974c49d77d1e5a051bfba21bbbc5c3c9d6ae253bcf83194ff641126b6eccc92fc7de2c0767b8d12638b1a1dbb08270e26d85115fd09b2b18b65778bec9feb4fb3b1fd48dacee28f9becb097d0d0262a92c8f02d7712ed015087a2c4636b8a61a9a8ecc42b1a9305f742bdf4f60023f034665345f22dd08162182346af8a024173aa5bfbfcd7627caaf9446a462973906679581bf6b695b6719348d019847984edfee257d1e31b7517f2a7a7f206102495a3f201ce89a5473e88011fd5727fb45c39ce1d8a88a0bfac09ec016f97eb73bfb93fac3bc8dc027ec6758396b6a9662cc984f2b601e3582ab5a3df5b73cdaafcee3299d8fe0606ee981ea722caceae104a98beb59292e897e8e29ee468a98634f12c59a49ad78f3868b8fd4355cbfc77d55e19dfc0caff691c704b1da3e4af94adeb90eec58d36d015970e7749b271f767defb26ab952624655c1e54e60cbd0812fb5ea6711143fd785cfd6c25ee26951df8aa3b057cd5137703ab8b1c139aada196a26d49a71655dd1541e4587b719a0587ddb66c480acfd50ba62c6ee459572192928cb679d48de320d96838d868722bc4ea5e671dce1fdbe5e0a6fd1bbf2174e5b292e2ed2cec08692c74907552885f72640d0c4ab3526c98b4c1080086a2544918ea300e93b0d0166cb2278f1fb023042f16fdd0c47c56018f4a0c1f799e1911eab0ff5c0a3e1db4cf6c7f34d2f81dc340b12b26f4177be2fb1ff376bdb1b7b7391f9f60822aad263acbbfbb77193bbc54e172a390ac3e6481339ce304ef832df6f15d4d9de8163dcf967e0e91e215cbb169e86d5a941b055c69c5f6229248e793fc1211915a34e132641a226c66ca4ad2fe98d7a2afe0b5af3d3cf276b4a505e63d367e08c7769f9388e42a7e13079d13abfbd57e7c661ff992b877389589f65dfa1d7ce1bbec14bf495630a946f9ba36c22165e68dcc1156cde1c0b4bad2d380dd00023af40f0cc42458472176949126eadf96e80f33ec6294477c4dba0af61a7d6866b679aeb561fd965149e539e1ee9abc0c12efdc7496baa7cb3705aa23d4cce88bea3fe3b274efd3b378567fa41ae4b304781aadb90eb8fcdb176987e32cb79cf5fc82237233;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h86a1461e55e1f0e0bd578c99b2e1cafd7aa4f49e1424ec73d4adb9118e6c8b3cc77083518a18ff91cd7195d6a33b183acc3603a02ef170d38e8accd02445a56f42b9c28f529eded78e62336e2285567ab3fd9a545da6b5a770463d7f9241f94a23becf8d09bb64465ce1ae0aff70eb77e2522f91802ce8bbd8cc8fd5acbb5902d07efa944e534a82d1027a29d8e6df20f25c124df9936338729087cb4e3118b9554b4fab1530f48627706321d24e06c9de80f7dbe35db2ef87b70a5495c017b352b286ce6ae5cde7c31bf651b0ef668fa92d98576d3d01fa3556a2d7636537ca8f9c0f0e27eb044fc5c6a88147af315effdf6b32c740425d7a9e50a6a0b0b516eb4b0f90c2c4bfe6d3071f9ea0874d239d96c3d48342651d51245497dd66933fae4f699e40923fb48bd1d9cda64934bd6d3ca95e47219ed8f2292e74eb2b5849ea4ceda44e6974c7e9e9e17080231dee3543490f05a63ec8ec481bd15fbe0a84da5ad8c6a2608ceaeb615b96b1d4ec619efaa75c9ccce220feb4812b811940f5932d0574c618cc35e91739c0bcc437a159a6b3c9438ad66968806022f1528761cf1248d603b0b685d9bca71969c584cfccd1351b7be40be33a56e942dd38206d839d34193f2b7631c5148619cbebe8b6e97691ede436a0b3ae18653478e59ecdd158e2ef9fc5e882fd94741889662eef76db48b0b4dd6d5358ac28d5d83422d5bc588383e0dfbb7909b4e546093b06b325a1ef87abadf49c228f9be71e7c973680413995490a461499d31511e425f7db2f555ab94322dc21c363f91d4f12a0c63884d889717e4cb45003ec8402e0cae5a21486402ec2adf29655e5cdcdf9f4f1992a0a037f59232307a0079bf967448bb991c9f39352e1ed5acaa64b2c6e72b505c005b8637e63d6b6f046c5caef7871d66544124b82dc8e2399ae3a1275cd7fc2c0cc83a4c2328c7c0958a98485e73329e5a2dcc0eb02030a87decb590c21d6d621dfb98ac1017f7de1758e9f0e9d17e87a28ba9259e4a9ae9009a83e5699ddc4a25493226390e234a31c37ba8f594114d89f95833a9ac38a56a9f5bcd0a7a8110675e06dc313749e615b02f41796d6b4570d5ef92d0920d9a40079f2417dd7efccef2ceffc80cf51324dc7810ce335bf326eac2388e73f32a7da2ffd49d1ceef32081583c50b2223131d193e443a5f32c9fac306d8621de866dd0efb03cd53ef1c91989eda25b1b6a58dae554e2e9b071a39bae2eba936a8aaeb6327abb43ea82cb83452daf666a56728d10268a0cfebd62a2f9f6d139dbafd477fc852eab50fe953348821155f5d81260889d475b2a92095dbc1201eec0a94b28ce95a6cf5af1dbd1627e40b60f5fc8882183c0a6a3136ceef55700855974c88c33bc0c163b9f75e9449f1cb5ace93a868dd39bfeadef98fdf84807957b8613e5000d3bf9fbcf17d3ed143701d37cd5919699355286e466ed6a78c98df9fdaf1282ae64d07658a8331ef943c33fd3979059b0e2303402c0091dc470bcae30ad1a7e812813d6275e6ef0ec3c02b75916c325c1dbbf9c7ab33b01ab9520f2d935b5d433c7c998bf08dd46a8d9221edccac7ba3403fd10612a9607e5e4cd8a12d167e6038a5b9c234644f1234b76652f1f9eced9ecd32abfc1e27c2e6f26858a7be425847cf6e05cf2ab633b8b0f36e919dd04577d448cb04857c35051b945f93874578292cdf9ecb8c3169cd9f0d6eac963c90db845b45aa807230185bd3081827ede77bdb8a2409cc8aa4cc515ea378bbbbf7e6186230cf7e97df9e9d0acd7265bdb10440c00c16bb636368f85db8d3e66b9b10f756779159c74d268466a090db830b602267f0e8425c2fdb3b289ab0aa397829f675ae92ccc330ddf4b2fc9848df78a97c6c695b64619813a062097f3873161262cb978da823478090af77ece7525cef9602af88325aed102be69c6cb9b4ea2b9467f9a260d75e87bda5cdf24ac5a42a24ae0e228fa7f01c1fc1df9b490b00866158c02be580633e36c2950ac6998b97bdff643685b096ae37df8ec4a1eacac0baab88cbdc5aa5f09c3f2ed6febfb4a9e1ac447ed788d966953c6e6784455bd5b04606ad23a56e9b0f91b7d29ce1302b70a1ff3cc3119b82416a904ba2fda3fded9c2afa25a5d9021d9ad07a4c08df0822c96d87d4e7ad9483482907c8c0bf6cc255cd5ed4e1954f3bcc0af96ce5a93014b799f3c372cf6e6533d533a835118d4a078d8abfa13fbb9183a42b55de94fde4b83d21ff438061eca6b60e858804f92267d95689c1f378905908a282d230893d4a526fb9443a28a5de099006ad6bd474e318a7c970ceeb97280515426c247de371c7c9d9ec1c383f952995a66d7bf34cd235c66098075eb71679f9f3104d12e13d8ed9cb8ad720cbe5ef3bf2c0552a7092f107d17915ab546352984f713ed21bac1035d2495ea942c0baa0a29dfe34df38cc6645bae5559cb3da56b843c622f3a5a51bed64022954dacf2a72464b468648c788dc1e0784cca8fd27ed73e152a275420916f496bdb47b26686cb893307cfd43d813698b6f837035f793fcad62344861884828ac13ddd5228ebc5a4827ad81f952c240efdeb21483b48a4eba7718a1397b8ca2be78d9a9725028c8af8a0139ed0d32a86cf81664bcb68d2d16b9082e164c40486921afab14ef4f06256ada7244dab5b0be569378ddcd28fae98366749e4e633d100c6cf898e3b8eaf38a0b42a8c44fbe0724196a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb1e8fd9aa2c1544e94dc968d2767e9e2ff107eb6867b71269f1343acfb66532669f2a7f74862c3d4c907e7c4e7092fd0dff8f1bc8c0e5aa052e37f7a184d9f1dbf0bef9f43f606f6a67abc60dac74fb4acb953d9d5a427a09ac5761e75a4249d9d29c8f16d17fddddfb863ba5e24884c0b030871f709d3b6353bc2e2174f730e4095fa7eba99985eab2746ddff66bd28e9376d2e1841c0d2fdd2c379c1559690713152f9c3fcc63a8b43f83dcf464d1ee5049a828e6eef6006919f51fa793eee4dacfe56f836bb82a1546cdd7313f509537d7ec86bc9178ccc55952d7b620ebbb1d3725024d63a3df21f75ef6ceeaeb95f166ccc3a4b24ba5d094ca7466f40aa0f64b4e93d098736f3598a9b5a8a18b67a75b3d33d337f5db059c629112f4475b149c657f6f3499dae184fce8c24ce68e600859a7ed73696215b7295098c9aff45fe9d3bc8833cc5adfde1d2b43774b9234d26ae3e11eb558d779d137e4af4cabd755d4248131ba33e9d55e442832f1670526090b6aa3e16acc03418aa205263762a8be6dfe5f34a4464b50f3b0e9323805060692a785686036da893a8feda7a99001b136c984a9d93716f75c487160a79e0c6f755653e44a7ab41dd42c6593a07f22e3c0d5bf63f8b6bc5747664ae78bbdcd61e9782500ae5cd347fd2f5f5725623663f08fb8f759d1694c77d824871a53d2b293bd9b00107b554890b69083bbcbc6ae7b6978b96c27377058a3bd2b4e337fa6f54f02056a88db6396742aeeb552f41813ac4f9c3fc12d45667c475a989d5372b2184b6ec757858b74538cc955ecb1b2b370e37d7b4200a6a2c9d8354e215a9fa78fc83526b701bff7b9a360aa21fb70d6368e3dd35078c5a7b8948abe574a8ea98eaa2be2ab1bffda41d59a64c5f1ef4b0cf0c2b26144ac84d67b1826d0d38fd647eebd1708d345667206359291febf1d6d25b35c383ad324a022810530d7bb909337a5229f11bed04fc36c5ee0ec7b827759444a3a16d42be39d50856fb6efe670809d485f00208b44e232bbffea0666be193330f0dec04702b7b53a6d9019caca7c3721da4cf09cbea1791ddd6ac8f2c7caf0a8d3ef336ff6f89053533e0d170807a1a52751677c7bf25cc05a19638d22c072f05b03320a1bd14595282efd8eb0c64e64fb06619be3da21bb86b7aa6fcd2d95c5b01b283e03ba692c256b3645c32a5976140c997838f6b733bd1c98e05efd10349d3bcfb7e7fcd7649fce42103698bcd2771c500a4a2347a0edc691ee1fa661923d5253ccb0899f0052677bab418004bf8aa01ff9848edb7bc168d541b64c06784de325135ca56831ba0b2a9210d45063fdc5270ed60b7bdc696b2f2c7c420274c1d7d5c9d449e39cdb7ddee2dcfa8c6752613a3e1a7a4c8c4e93a17a2d274feaa9c517a8f06ea2fc1ff5b09155fa289bb967bb1f4d365a26f5e9affdfc1282f9fa0d4739737b28e2b19119802c194ebd825a36f447bbf99f4f575626cf760bb04ba77697e5aea9ab2051f43550761781cc9f20ad77cfaf2430121cd031e05da26d6c702679af23a231824fb42e36af600726f6a4a4a9d3b37b486b9bc7864350f10e2ec0f11b86fc6e155955bead5870598815bfffb112021ba99233badbfba3eb8dd6675bc703aebab6c5daccd61dcc4e0b68a0d96089f508c0db1ac3fc7a70d104e9d18b5ac81b33db5f43a6934d640c68123ac1a61c1b5604f6fba4ed165eaceba3683254d115bec4e5cffa940d07747b28e1fba1a2508afb52fcdf82bb4f014e9829b5c1d0c42e19d8697c9e4bd61e5944397fa33cb95a453dc56488a75157fec661a0b7b825751414d598ef05d8d618f0000df60392afbf35e821abc4a686c789a0fa0ad94b04b663d3e4ac48b155b3cdd53c32ea5487471a7371cacbee5a04cc8be4d6174869f1f57de9ed99a7d908a013aca1a8cd2db9258143b1fb54bb777369e0ef13ddfe423fc002d9a43d48d04701aabe216ed4c8910dfec4c1d005edda9862dd17600acfa014fe4434036d824a3cb65882774ff61050c983255646459a892a771aef2ef73b23397e3a35c3cd1db5ac375874265f53470d4a97a538b27c27325d3386ccb6fa1232f1e42c1c83e96f4d093572583f09dbab2f78c0a4572c8a534fc7ee7751a4e68dbc2954875966d40228c55eaee4871157d01c0ac1a8aee5349f1b59c9d49361d62f882781ffb7c636efb7fc2ace23e3762acdffeb8130ae44ffb825a95d8fd0606e3dfcaec2989b150d2ef7e21ae8d8154a399ec14a31a15f112b9ca0ea2553a0ebad6da03d0da644c83bb084317b5192edc48afbe02fc84f205a3a9d19a97c59ef181b98c9550988c1d990468440fd6802ed1f615854557a2c7dfe5f1855140d2a15920eb077e9dddab1ddbf61a7e5aef54dacc68ea284312c1169061cbe0604af2e961468f10b691eeec20d004c9f56ee46be52d39cfe18fed42f4809ceb655be4568ac3559347527a5dbe93924958a4d0c9b43b5ada82ce970e88ca227cacab7b920f6f76c9b75641fd409a83ee2f5a2523bc74cf57e0e776bf7c2f2a8936561a0981a31d68c150e9a4d3b22f4ac853a2fb17590f130db8d0751f96ee1a2e3e510f78bdfdc07d7e5451559f87e7d7ae9cb139b77abeabbc7835156fbe71b5eae653fffc124d552464fb1527e3dd5888c32c194a0f1619fd46b015aa36c33842b873d6872c244e218aa3d0bc8b1f37491458d865d380c85c9ca4ed37c49658ff11f7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h91aaabbabc62c8b0523783980e933547b7966f8c17c7d79664248ae645defdbeae7aeb48eb3af7f0c1b80a82f2632050e2418214337c980ba5fe64256b1dfd419c5a9fa087adb736ec42b187c5ce0b0591bdb191c4850ea1102e45ce735b41f83d1cef1e688e485f7c6c94437657eddbabed27b82933d8a86711353a23f27bebf23735b6cbd0f271ef2099f03953c5bf01deada5f67f7ca0e08341bf8a6448438bc9123b1b0b996724607deb61adf6802245433eb02ef1195c11ba95244b198591377c09c88673a18925cb9221ccbe7124d99dfb0f3dfc1fff85f5a9e7f0ef460da54f3b427eaa71186340430d2c6f528731067b4f06306c30b4c2dc6ce183150e6923cfee8c2ad6ddb3e00f423201aabc76e8bd16fd4fb047a5900909e329b4b1355a4ff977ceb04b846d0c8468c2e8266dca21838c8c52a3c5865925df4de9a30781129c4b2fb439720c412c9040913f3663f2fe6bcc220ce3025bed88a7d6bb3950330902b0d62f88908053ae9a1ac8b865a4ff23477498519721e4b1da79ea68038ec210351de98d3a2dc8055dc3f699e89c553853eb6208d2f490c53f95462b78324a8b10d941733f0d7a87d14de7db774f5e74e157028b3d73ccbb0f164964d7b42b38e9bb0cb4d3de66c2d6a171750987b7d063371f0ea5b430d78d3c29b26770d320e29cec58fc585687284119751448765745c6babc50fed7146afa218aa6c2fd30c59b9a9f55d0b502c8479b23a21bee6cce48db1c7f6f19e48718a371b842532ccec012dc2c7cfb738864b0189a5483cd0bba5fd335fd219552c43e711fdc8efcda1691e930d7d6f6076618a8dfdf263da3503fa6f1e8970c17d37df14b3094b489739f6eb2979b4b6a15e618c9b98d377f5e13722e5e861f472e2da9523a2eb799e0d153744b9f54f9a9b79c4e839b5be93c70af9b19f795d3db5bf9596c362b90e3bf14bde3666d85f0ee42d4c6e905e3686dd50dcd580a3a43273b33e276703aef276ac9401089b477c703be1be4b3b716c24a5b65fb2e4ed90fa3445eb177bb1f524d12eae0606806dbf590dc5bbd2d0f117fd956555b0f125914d4b2bd906724f60e8cc09b4bf37ad5a6ae28142bb7d76d4dc0c9f9f9d98daacb8ec548b0f29d8b4e8bcb9b8976fbabd62adcfcf374c25716156ecccbceee9c52807a92dcf23e3ca3b9c6c3aaab378e1ecd00f2299a07e4113a4a611bd94b454c5a98673e56607f0cf0b3c0663247d8061498d846bb254f792281b4807b696d2a0b25bef548088e32cb584d4ad32e38eb1be261577b203a671a5671a65466a299718e5d3f2b5d378b0e4f41b952b484a5215439e87fa7ea5bdea703a9da588ea655c266163c8ec663fb68388f19d021e557aeaaa2d13b1f9d73bcbad56b190a615e5a9fd51d912e6de6a533d9329e52fa0787a9f0248b6cbffb85d98912370fcd99f09948a3d667cb86a433ea4dd37d0be8c73737159c41e4e2daa599bac054ae38d22ec06bee286e07bc21206a5c2dbf1e46a84f41fc73f22ed46caabd2581eff0e2507b207c2de210f32f4e501b1534d0e8d667af2892ca8015aff723a58a801d9d51f2774d73d5a03a3607a5e70d7dcefb78c7d95f70469ee7cda8721aee1227b4d7fe42fb3271e329a49d96da4634a563586ac95fe0346ff95d1e2412b57861038248c6c8e2e2b0be3cadfe773a39401e9ce36f7d26e20004d05d3f5c3459fc2a93ab662804be84796d0cd8e4ec9f12f49550f1cef3a85322e32aef1334378bb73fc308b46c8008f4616d5bb24ca362041b405b1667d35b55c9df4244c7342e97ad34059b1d86c8a6c948bb675fef5cbd6ebc9e9b2f5615af47e67bea3bb59faa899d8712ad7e6fc9740a959844146e15b63381300507ca19374d61a29989997b23e20adc567d3afe6194e417f48be0f2c05a5d02ce82e1c6735de13659aafec63b50d309a5cef4f8902294c954a719520ad4f8f64c7340d4dc21287b6e43bd2effc7d2937aea97062a28e08c0b3ff112f294907819090d8acfce8b0824f4bffbc2db1acb2de65187577fa9cecca15ba41168460a6831ac5a2f8b86ee246f8ef5fe3d77bde43a6c3bf513e8e70e1d62326959366f93a3566ff0d97e95a46d9f3a44c8572452915112be029763d0c1e1cff3ad258a919a2b4b9738736a4622f12cd15e318c392a119e73912dfd35224151c37ad7240c15212f0b74c1e4966466551bb7589f14fc0aebcd046008a55c630cb7652bb400d95eb1d5c7ffb41010fb79df16565b11a2a345cac5921fa669e7457839f597ba41d7e81214004184363e5063d6b99fe04e6e5b0a4c733f71189d374dc3589cea68414d5ffeca9bad8f6e1c85e13e5de57247d6817cb311e40e0e2567974cefa623635773dfde2891374215cf0a345dbf10b514f29dc58d0f9d1ae3eb21144958dcf89d7c27bc58cc1322a4bb78c8ce7ef430b7b0e661a0f2b0bef1ff8c6f2072f714f636f5c878458abf8217943f8b9d54ec4f669a3b8c8034fe98707b2578c76dd6bb79bd9c2ad71749a4d39da13b2cf268c31a8ba4506272ce1957a3046dc94fec2558811175f2f82ca1e3ebaf16b00ab856c72d063c532403bc34cedf0eeea2178316ab6e17f8dfc4ee391b014c502c7401046f0387f462e9ca0745474d63e6dc1a07a45e7e0d151c471c1c782d567b2b5c6ffe4ed82f91634637671d5abe149a9ec4bab15f6d10cb97d8cb8dac11bf38e86d8eed6a3e08bb45c5ac916f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h5b9e6ba9275f17ba49cd8d62106839fc867efa4eb1202e4e79e406256a43f2f54dd4b433973f7f453057a753d28ca86092d557c6a95c86f4ba82f44e04aa67e5d77ca1b4fba5c556d61526b30b01ae7a8e6febe7827818af00a5d5e82da23238286297aa6f951708f4bdd5bedd805261cff5a1df865a2139370e8f337b728c04dc32084cbd4629030e803b0e680093c9544ed282733547b1ec7687b64b535aad7f02b2c41715637310cc63779c372ec7ee7f9837c98d95383fd31da8bd1cab3828894855295dd5dc612c62a0fd6874f28cf55db8ce98fddce9b8a9894409d86104408cdad2e3930c7993fb706f8206c8a383860974d594785c858ed8a43ebebc8e6302a3b54dee08e08aa8d05b5348f470ee2f6318d7f329b2f10b1cc1b787d98e950b7b3fa0c7004f896c31c30e0f4f9b139797ce6f65fb2540803b54f5c802d085b59225aeddb99a87cd303c730eed5a2bb5e577aaace435d5772b903ae3ad9c93ea860d873b7eb53df70020f79fdb77b603e5eb7b60bd63e0baeef48f7b65d48bd8bb42093e2d02d74b4ecbba8d401cf3917f6d1090d0b70a2c4648ea853ccbe3e4ae4d32ba64d4984c578ca73c3dd601fbf9e50a18668afa8ea39ce25257b7978182e6408105b48606b3af7f56f7199c0388a5e713e22f8840cba7ed3b092f3be64cb1a74c0eb39a5eec8bcd8bd2e1d2a50432a61af77521e21e07edacdbedb324513f1104175d89348399f29b113f4c168980c6e16bca736c16b9c816d5b986160512292c9e19d07c64b35dd30875fcdd264ee29e16fd4411cf8e96f6121cf56505498a9de5fdae3e4a570d350c8a1ed197e3008fbdf1ef3bc02876e0e0575a3a893a8982d56b34fd71f7c1e55568c4aacac15d3fe91e319cf2ab7b082f0a75c83f4ab1f420c7fb308aa1f2c0881cba4b142ec4aa4106ee03bfbcfa03803a9aac4ca0eadba731be1b60c34289ae234bd2832f4e98b61c5300180b9870efb4422a5c855e0d1bce0b0e7daca1533dfab61958ed3f21562b3ffd19cbfd4695a19e214c37596d711313441ac4cf63863ace259728fb756e58ce0957bb1f9838b46e0d419d4394643fb81903e913da524dc8f77a47246866dfdc9eb0df04cfe9e6cdd69b385500146edd78db1276a5c83cc179b070f6fa2d200c3693a119190b7a82a8b87198debd4ebcbebcc11cb5b0ebe2ebac6eaacead439d8cf3b3121545d01a4da65d5d385541ccf31944a8c0c52851536867b34af01b68c1d423511b40b734b9ee4c77bbfa16830b390c3074a756c3513059862df8e1c145874090b68205f580f0669a366df10fc12e34f05f31b6a3bd72b1446f814e35366d6d5520d4849860886e25f4488a3357cf908ba4c77553cf10477d7c509c2061fa4f740a1f2efcaa597fca223e294437d5de6c149659ed7987787c36dc013eb47be190441b8a7dd43869cfd3b96d1f03dc32756779eb32b341b8388106d0930c2e1020f09dd8d11c4843a6e10a1f254ce476d4c95f1138e07b43bab09298a1db817bad1b887d8d4d9ad07bf7388615e096bb193f948139f43cb360d886741cc4443c944e4a6c14615cf98bcff12afd5c9844ccc0b3c1365a5769ef525104c89a64fc208f228f8956fb1cf78f334580a49746857c595b70517fad322975ed167c9c161265b81b95f7a5a1dfecda46c63bb9addc2ecf062cc29479c2315bca97ad8168b135a72f418132bd2d2cdb3cc2574edce24287d7d2fc24ac654d86900ed0d68c7b9525ab032cb4f2abc9945b75e17215c737032f0123a406a5e19c91029cb90fe3ceed51fd9e4d01bdd300daf89329a8376018d9e6f6b2e6e0b8e91bd785fbdba031e7541f6f9985b3d985bf9b22b3b1ec2c0106ee7c00b7ec26e14a1aaf0efff2ad72250d2e683fb492ddd32ef820de6ef57bd5b6c80612d1a71295caa65026bef89b586f230433ee2ccefc80e7c514f94d498ce40bb666ef5bde986d0a72168566ce52a65588f5db25cb2a831dab6acf268b92b1172f85ab3cc91a82565813761eee496d81e8b80fa29596a145330107aef367ddae4da6f1d8d4ccdcbb5794d17239cf5bdffe7444c67925be9decb07d08389ac8bf933429b9d139ef31e6348a90f079a4fc8a06fe65b02563a7585895e4857eb6bb8835efd603c1185fd6df3f214d01261c056084c363aad76b6add35529c948adf203384603ed4a362099f45dc6ee4c85b7ef2fcf040ae00780507d203b96efe78626bfef13f722a7f44f9001f98000e9c89cfa59cab8561cccb61a96430ee3c48977cb5154722005bcad4a58ed217ce720fd6dbb04487f51b5f1a969ad0c31990baedd0bb7ccf24fadba8cef1b33d60bb42798af2a5b4aed1e84c6dc63dc472c09c46eb5d76733fdbb4ce42b5b50c4f3a2ae0960eb2be9b438e1baeb40812d5e250dc918dbe20967b7b9720718e82a1ea1753595b7758635e6bb76827fb894fe807dd48dc904757abb62c81cb2e8c37ac37305d3e4233250a7ed90f3a22d4e8a4f89c033e21c15930a0e09ff2c7aa74e680775963542cb4fa85cc000322e64a38728537c186c4a5a79965b68e8ede1a827a1dbf0054afb6b1144753740a6f7062cbe35293c030a0cd9ce59b6c67c67936873735a05704c705346a080e56c3b512ac382dddaef26f19af336f899a59105dba1670ac945a374dc499632a93a6b6f6456d6158931c772779f4c910e4f7ed5dcceef59104cadeca435b71ffb2fcab2ee4ef01cb18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbdaa3e3586681b0ad5b3f2856fc545e13c6d0898c7681761f6a69f220dc37633078333e64bd9338024e2f111f988638d913e95f6d37d67c0905f6f9f0de7f70bfa05c00581576c57e04f956fdaa785e1e7d892bf50f0a82e0f26b743b3dc045794eb7df2b836863e6805867d006d26f12e8fd343ebc3aaa3a72c8a92679d107fb91d872b179604e02758a44b6ef2326ac9a943721b4d32fe96167c73b576e4b0bd55b6670bd7cbbe42a488a66854f37e9b3c4edd797aa006737c8ed64634608760a54456c8d3ee35562555e2a962edc98f6491727f5b6ea63a9803db917244fe30faa160e89692beaf40179131723a46b0812bc5477c7df3a8c9ec7c1173cc93c4db8ff56cbba346e4dde1ee617e4c64a3fa48cdb7354546f9d514f6d3b10d003358b1a0de9e6de4236cb9caaa752444e6bdb9855c64c1add3c878ed9a36f923e388ffe4e61490237984e0a163cb2fe1fe9da4423c4f7a1efa5b9b5c1b6484f881c0e1870fb9696c06579e325115e11d57dab97f931ebe2e67992c179d9ec8c3f1ce5bc0301fc26957df178c84cd6a7a55730df2293e4d73d7f6f47571c436a174f07d59b4bd9a60d7b7b6eea6b20b3704126f474c6ca66bbfd880ad5d09c83d2eb8c25709d455d752803004ca037bba62728adfb5d9ddaae827e4408490af571cf8bef96fc450cd68d3b67cb236e923da5ec6fda8a6132d5739930bc7c6f001321c18b30a15b7a2f1707a4dd842a4c593133b25b3ffdd8ce7f4381a9bf2e92e59cf51ee6f4d392611e76b6296d4e293ded8e5d23b9815078aab43685e35f3dd8d2fbf47ef866db40f0a0adeb4d48de45fe36cb43c5cafa48e2d3184b1e5e791a71f93df22a39f2a762a288d54d9855061c8ed741ffd78a9927edffb3351c0435a5902e21645168f9aefe0f34326966356101de8dca052a455bd89662e83ae075adbc9f5f37262be3f787a321a8f286443b5bc035aa382b79aaf2973c1d682018219f7f58ddd26714c883e2a23b2815d02c7a28b8c230f7d4e834f2d8c612582ac73d0e69111b08d0f22b7623f9298d65f4a078f6dee8ec3c11fb3d28e6130c18db158ce332dafe36797320cd88b1843050c3a3ac0169b36424d5579ed8a4fcd4864d5d06d9b7739ae84180964c72e753ab1e927db369f1f65d04823dfd6671177114f9091d75442ef40e58d189b7e39b561189469b2b49cdc4d0624e76121afe7a2a70176099c6b82dae5739435f4337d0645976eee24215341f8f80c176ea01aaf44f8838c1069276d4d5d539997bfba3af76e91d0d24609c4bdae1f255b1c2532650cbd4f69f724fd8109d3614c9b93987bb77141a548dcd1eb7a62ffa091c1c41785f074cc50e821318a6013ff8c15338def1b07c916c11f482830994b3c4b864b343357563804f8ded8e4a155c799bfe495ae6537749fc73ccda520b8312158d800f5954ebee2c38d572928ff0c488200c19573bd0e46164caba1f1ebf2e718d1f7dc313200da6be8a63b02f76eccef4732c5a55669534d53f8b5edfd3185678a6b295d542cbf2750a3b941a93191722cf2d7f82d8c99d25e32462c7bc738b91b1780fe1fc29f4c80ffca2dd6a634c316bdb9d8f19f551b2b334247868342106712ab8dc1ae72e14f092cc8e4a8e5c5c350df8a727c35a80438c5809edf5e280d4f9ab7bfc92f9ed8b7956dc20c2eb4a85cb0b9d2493d9478551641c19a17877961efb60e0cb05c70491b927bbf698cbe078136cc24d87b6b68339fc1a967a598d3a557c2d5f197a1d128231fda758a5af9378ad779eab336cbf6efdf12820ded10a4ac6264c31dc7f216228be18c91a68c5f37c9c12a04b58dd3a02dde191e0e13ec9483402177d8ec148c90c96d4a961f41da92b7e59240aa312cab505db0848dd0160e5dcab1b0ab78ad6274c00a2c89946a20b3a01356805f84e136537406016b68b9bb78013b41543a3ba39146405aafc95257423e4f7b3fa911946dfbf4184439bf14340eef5b13608f6674cf19a3f0ce1a48f8727200d225a3c411e6e1b169801f3f5d3de44f93a5b8f255478a49ecd541dc484547e4d2a6ea6e0794c4b48f76f9ed58406499c8063698043c86f724d79f7d5d3fd09be1f508412acf68a89c13385068b3a2ad5028ed408752b044aa9e22362e470a03eb77e306e6027cd922cdd9d7e042e07b37c6802fec921e0541131f08f0a42ffae5d98344accf30704a0a0d3cd2abd46ba05274a990b71397223ef7899c54b515922be5a6b281049b44fe6c26a787b1b0f47febe4aae9d14508f14dc0114fc8d2dbcef79da8e494cd710b4a0d5c3bb2d8ac7d3e0357012ce5c129be6f1a028cdca4f183bd9240d9c9e3aa72467c99e4ebc95b06beeb339b45975121854b6f02f876171547cd00e587268b36c84bb22cbc68a5e076ea08ceafbc826246ef764dd4f0e6a1516c07670cd04e93784a5e58139b6a46d47fe65f47a4bab90596d318a89423d44b413ce2a28b85bed2231033c1d15bf149e42fd50e3e346f02f147c4522acb41d9c40ccb81d9e1ce565b1da683ef19a6a9945c07289d22e7ef21e1dbf03d9fdfdae844c0318c94ee28159aa0b08905b54073195d747f75f448c5918b9d08ebdd08543d388f4216ac430752f30f4f7346806808f55f9cf12b0d3d8135660cce6c32d2cea3db5c0d297cc6d951d3799afb3e1107b754ef4e9d353e93fe758d86f4f47be79c4e3230fd41359f29cdc22d259f7cf4940056ca8c0c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h347ede84cad36eae7a9e14614f215f320c4e12f1572786b4f78d29cf6ecdf9ead783f85164ffa6d9a184fb3497250bcabca178180a481610f932f376a48047674b57abe879f816cfcd4ed0cd94babddb205457158d348861375278a4afa5f03db8e6c0afbb25a98a5708123abbe1e424b2dff94564306626e26c42f057dd7d1c8039874ac5f93584fd86ad4dd31d3c8d25e011093b408b0884ef7be92402c29012481115a998ae15ffc892fee41ffaff6511a001ba42836057cb730c314492368d2399c92b1edbb5842624c52053271671ed475d62224ab8b08418efd1c204f9ff7360596d444a89137c027977b58e300004f3f68aa3b9b2f995663f40d85e99e0151f9f4fadbf77197609bfa51680771f238baf7f6cd1ecdd3f757c694f83dcae10ba8d5165156f65f5ea8d27c0d3be13bb5b4b1cfc6463adbd82b59b9fac9e9eb853964a15010c5ed31cd9e694d5591c3ed049c73670a3f84a44e10410ef80a289bfd783a05ce524094bc9f2dfe9971dbfc09bb09afc0351b075a9d57c6f50f5c2785f2ea22629a90feb3a7ee98abe763fb145735012abe4f6c1f2fba3791866d56444c968c4a4fe05ff92ef66858f5fcb827a162e243e0471f0a01db5250de0ac6dcafc3125bf57c2159f88e50aaff8112f2966250c88be2ab3bfc1c81b91b931cb05aeacfae691abec84ad4814e36dd9d2dcdb29cb62b73f0e86f489dfb487d068e6c149507b9e7352692c756242231379af63de4b64aa16f3088724e81a3ec5b8dd0b3fe58a3f467d83845cf4f0a04bee1852cad764b8ce65333d9ea7108dbcf24e1b15622ff62c44ad5f8b0c2cd70bfac5e4c89a16e37310c39525ab78def6931432c559cfd8cdf88c463d7ce5a7ff054c93720d87954e041b5d5b1b456cfe1e5c716f26aea0cacb2d1408b71d8a7ef90cf6c9261f6558c8f4c30e9e75135ab70257ee9bbf460e5025e2f81b8d132b996771435b47ece68480523b60b997f904ea075c0d5ad07a17e5f94638efc33981e549cc6aa25be99ac09296f8e0a964477e0f7c3e14cd1391d2b30c2b815a2a8706b28c823ad627f820c7e1cbf241db11ded323bd04ceafbf36ae6f0135b94031aa82de6d7ae6f693b445dfdad9a248355203b8bafa83f3c864a0e49d3d46c0135dca7f67ae1a8386aebd2d1ceb8d41c779110979c7b92d1d73bf5c6d91eb025b48163f1b6a1ce5f15525be441cf46e329782ea64407e0e0b9e6dc85b0c8d0de1b9dcffe2754eb626c86dedabdb415894ad4bad03984e7e0d4312b3e4f044cf145aa33c240d5dada4cbd78c817a4f5600512ea70aad52eb10cbae20fc76f42e49ceb811699630d4b35775c3a6e6e5bda43d40e2a08c79ef3881ade19e0060e66e80201545919e20bb87c65e80dd60955922dcde66f56152200bf35090313add90b22a502b01b23558cd6d4b06df9ddeded24d88874d7e55ec6dbe29c2e671922f2f5513c49e362e562b9361d35ead7b94003406a43fadd3719795bf72d822a09a918d110d857adf009ec20181113dc409fb8cae3f9af00805a8d74bdb67fc9e3471a4f08b6cd97e1e44c1d5563d704168fca58699252beec79ed0c9bee69cf2ef70a98a34391e6a3b3763948aee4656b3d6a0dbaa19bdec524386a8e0dda9af05184c9bb8599a6b90432f2b34a86421f75647920ebcdb05be3c89850f42124b907f60ed64ec754a5ed32e3abfcd7dbb174a7ace423209efecb08b74d498cc11b839dbb8db681ef34e5f2a5ac53ba528c620dbd8b2115237d0d20c85d4f4a081b9a1a4dee83fc8b887ab6b28c9ce889950d3341d66ede8460e7d0856b453e5a49eba291e02a52a84c60d40fde71d77d68b06c0ed3753113f9628630a0bc93773b244fb671b8b0870fac73c078351cfed752c773d6984b0a5e944d34fcdd13c21a18dd062f74d425942fe849d38beb83cac38464e4d3802fbcae8dd7f7af4f41a01663a94903189a536fbd538edd40876271c1b7897c91138669f6f7a0a94ce50903bb7f1ba17dd3f4b4749e4f956fc1c9f14a7f03b246b35fef280980e536c40bae12f904bca66cc77a450962ab1e470ea73b7fc4b5cb70c74db8e6bc12ebec509e5ff3c89365c2b02dbebc139710636951d4c61997d9f7db32eed0c14e85020c590ad16d52b1288afcc27a0254227cdb2ae5c43b338bd43ec15a45ee51f2a08708cccb1ed9b3fd33b802c20dd23b9fef3218086861b37c9948892330918d195f89155776f545fff7ea166cccf2c627a11fd2d0c47c1ce9025fd0447ac1853ea58fe1a2e86aa2f3c26519808f024aa40ee8521633b910beef2e372ab06cde6695036eb2fdbce36af759d11edea6a343b98d8d29132c277e173a0bf4cea18255ae5e8f31f810ba0e6e5ab8bc1dfa5d22cfd2ff6d4dadb0ba22b42f498315650a27259184ddb01cffd0d1488b0fb0d5f75dd3181213e0453b249e7a8c6f276d48d6156dba23279b77da4c6ef6148953ae8e5cd1555a1c34cb219a92360a967960f67bdb0bd5d1ebab093c4b2d64807b244d626f4102b6f5059cb1979239857eea788fc59d8b12a5e1f1d165bc29815c46498eff82daf584e930cd78d27f36c6ba27af49f6ccfe7dc8fe6d1f6b3a3dc4e4d5a6c0d51ff9521abf3abf816369a5df3a82b68ab35990f104fd047d34b85db6bae0feaf742fb8a332beb1687c7035c1e223e670ea02039fb44bd989317b818c5244bb30305a902c9cca6c9f4e3f01c7af16e559806be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hfcd774511b4c0dfb7c7f25668fc4532984c4fd0deb7c88c02c8a2e8261f17362c648382977e4d9ee52f73403b2ad2870467d736369a86b9edb668292c05fcf4b6c90026acec80bd879815448448b28d75fb54dff61f0035910853e8ae5e9cad10ce17ae5bc0a9b9c89a50ecc7861cc51d45910acfb15c80ac3f0041f1ede8035a0daeb80aee9afc28d8fe8ab9a9c6c89f7e2944e1601d472ffbf167673bf1023ef3eb190a24e69690bac5ba9d7ff319cc627cba9c2ac95cd13a4f6709db664229f3dd673105054bcceac8e7f72c40f0f63872eb4f8bd2f008042b5ba7240d01e3704a622ba9119a94a82670502f7c3f7bad11e7d7307807ec27405779d83ef11792a0a20d2c792f6ad21452e804d36e21aba1c6657ee00a2aee2013c8c78e46ad3106a8889995350d52a91cbe7fe5094bb74d2c49936008062778e4127cbf7a2ce8516e6d6f19cf9042d47271326c318f7bd12e7c58b5040419bc1ff9fd333f94759a9644d470544e8e7e63ffa8498a65ab8800eeecf69574b36a77e2de52cae9d19e9bb724b2f02130ecacd34ae8a20829020ae5f82df382a4772b03e010794155ca8ee8b4a131b6a934d07a6ee954953168fff28c3f8ffe2e458803205c7cca80937d5aae0d6bc0ad05285c8f2987beaa5ccc4e1693b90d7a5723448fa07af8bf1195014aaec1e87d6dfa8eafb50e98b02aacd8d0f8aea4b77e8eaec0ff4c4692af59a31b29777785264eb4717db573fdbb55ddbec31ca68964c273e2514a6c10fbd549ea1f44c846becb146cc1458a86404638665c4879decbf89a37e650e5e233db7127cc7bd77fb177c3e01e878120be1822e9b287a5925eff2630e28e4736bfcc5306beeb4c0eeb13a9e1ad29998c4e957dac866b6b40967adb25db41b021efd8158899125640e7be5839668fdefb0ca3f97a9bc74344d97fc593bc9152479ddde143e85b7ea11d6a5d7d83095b860970240e9e82f4cb1834d82ec33e0d148a8a745bd0aa842934be18eebde11b720e9cb3c004dbc5c3b12436448e37e5de8229f767550d9da1a540b2b298c5cfcaf7ef63d41855c7f32c28a0124b252f21177c02f5f2379e4afe18e111f724ca8909f239dd8b3de02a8b0910ca6c8993b815127e39d43f9782f66f26906acb60d430f3c0927424fa84556747fe2263e61e497d06c228da237c2444c9421b855132385dfa5a65df7ab8afe338747b6cd3cfedf599a4a1929f7975c78bf80b396659c0e49a07298a11834bc8e41d431d66813f7e8c866696171e11133a0316f14f4bf9c539077a0c1a57d7146e82f420a42fc1f0d57041cbacbf35ff90571bb6e4a755bd576bac13c49dfab77e00a4626e0be895434e9b0e8bd180731571aa74295d00450ab3b1af1256ffff0df3394d2e19a518afa2cf284444ef233c4fe6d8ea12808c79999e1d797850997ffca98896de2f6b4a2ba37406f368e65c1394b376ad81dc9f4f3efa5d098236e8c8da43927d6c1b63ce08cd2c619056d45b4ba936e07317b514e2870240076fea85aa41e38b31d0d17b2b0f97fb860fd2fc2ee9ead8b3cd1ac7e794561e4f8bdda1d0caf7f26537b9139873f95f55d601f0781e7fb916c339830cdff575af87881bd7ed78b3ae9f94ef55fd61f98b78dcf77398ddad5185464043c61dc3e03442b18b8e8c7789bb56da9a7e46a82016074077face03b1ac510220781ebcb3a8908e3ff0fb3cd04d87feed90af129948068a745a6448e66cd337a500f9f55c843827e7e17b898dcdd12fea12f82081759cb26528afbbe70701c2e73ac50e24e37dade16460bf5b607407794564f0e0db02ee9ef9f89984c53aa9e59266fb6a0e98fe14ba1d616d9205b937804139fe1fff89a875598326177353e6f61c1533b205bfd89e9e920838bd5ba6852ad877124d32f35f083abfb643d66157ed5ad3c432d51c30b6f59a009fa657adfa0002756ac913890a6ed046637d48e75323c2ba26d0647aa3e546f58bdfeed0b8d58b51407c4e81d3d1ddc620b07bd8971de61a3c0a85f0134d674302b9e25f647c12d3858277018b4a051a99d9a84d79ae0f511fe2b7ca967628300b1c263b62eb149d6c25e06b47021f1becf0e41cf22195fd180c6762cde79c997bfe313f08c21f0df673609bc22698956604c12f5b8d9128aaaaf456bf91c970a883d9fc729360b39c77730f4e601b8fa3a39209519be7c088503d768aca7804d4326e90561f43744af0a1dc1263c3c9ead8389148523b893074f66cfdc3d0d9f7118d06e62e3b424f47a2fcf5fca7c787d3918dfd61153a9a686d49c4a99aa0262da7b81366ae40c832b0d271fa499ba7c6adc4379178c2978aab84924730cb58c8dd8258acf0d59ba0d03146ffda3961e4d5a67df09e71de3ab50fb3f3a56e7703d2a782c79ac2a449d6d79e33847570e2e664d730a1ffed0b4b497d86aedf46913db45e05aca2a881213d68422cf578930a10541616e17cecfc4a43f70e44dfdb599cc900f27037c1a79f8f9ae2b94e823b2d922092cebd65b3392a8e9a372268646343fdb66708e2e0ba3f5e10c3d105765a594dc8c6f7d159e0855767878f86681006f3b210492c957c8011b5256ce1b8b1b0d70c17cf27763c1fdea6d80cd3c38dadabee6221b652080d8e0ea398001b073192a05d347b325be6219cc47df6d6e225c05ad1bd443011848d0114117167f29ae689fe00bc043d4a94b50b759852c5c9fd7f929aa9431d7df727f17551c5c7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h619b368a73a695cca7f8bc100aa42bd72dd6f7daf8598d9da8914d25d804e30c41aa55995ea451d7236ea21da02be70d83adf2a5395e438eac495f195dc43561ffd729b8edaf54f0fc5799e7f813fe045949280746be8d8498639913e743306432b352b264066e2d9868ea05103a19ca60576a9a3b4d3a83ec39de2d8a996dedf23697085c564ee5230211826f0316ac7a3f559de120513f69a2361316d97b7c4e54e3d049fa92a32396d798e1cee1c76f2e9b46599858dfcd133844771c09b8b9b45d35b81dbb02bbe5337936f5a421d45347f75e3096459fafbfeebcfe872c4493c52636712de23bcf8c8543a48f6fd09c982c30b20f164a7e3676f3ab4a02997cf451f1e97c4f73be7bc8f4c9fcdf842f4d874ec1dabbc609e7c25a2d266fae2d91f3a296568964a820eab5e7947b8a8ec889422011a6b8272e5731ba64b075d82175baccdb2dd026944e0a17469ea5782fbce8fa18989b1108e02bc6120914c88f1770402fad7123d4b1d6c6a734362927d106d04c88633a37f14d86172e32bb4abb6de7da662337a0460ae0011e58c10ecb413055b0a38534fb1225a450bdeabe56c1608a3de0a94157219044624e9d78bea0b74e82fd46cffc7bf010ebb89bd2cdf88d20596dd15a9e8e2bd44a41f57a715e7b333c174c8a5d2571f89fe2a57a7b5bb4ec8d53d549aafd249b2673cfdee0b39c1be7e6a3fa9b8711e17a9f3f8f38c2e621f5229fff1d0db386615da37dcd298772a7eb41b57d4a56ffe603d8b15740199be48648ab0711b0758f7994398c440942d26c3d12f657e360d8d89c46f525f928989e133410ae94d34e4f32c4598896c2ff927a135a360f687442732da867d80bbb34e74f0a8797bf01159d6499666b38324b478c17bda4d28d5d9cc292c8416cd673deb92ff1b048a724129ff78fbe450aedfc7e3d53dd47594c3cb52b6aa898f798495ac42ea7fe2ed2ece33dde576ecb126d6af4176484143aa9beb9e5881c9497f40879eec70d4653bee902e890eafc35b9ecbff833509e4442b34875d7c7150bdded5a893326d0d823376a22b3495b47fd95569b5d14a7a47c93646e0c047c26ad19297c5c931d4ba0b522180279d1ca6ab520e1a22767949479726e82a26be62414751cf16df5b7fcbc63b7dcd0e198e0df8b4acf5ffecd06f94c79247c516c32ffa361638125abe495ba1ae22300359103a142f5d7c9ea7e8ad61cfd795079f3f9b99b7dca4ed8d81e7e0b7f6c948858a7ebb69bd0f48efdec3d1aa9cc947394da8fa5e3a4dfaa68e604d5170ebefb3598cfe8a2cd3aeb89eb2f10aec69a7505bae4e66cc4b70875b83ba5f6f33324b09c9e70107cca21397430551a04191905c0cb0f8fc061a8539d582b988cd47264169f7f501fb2955c4537fc8bf9f745e120c3b1d8982294a4250f111115e1f8f8d6bff7d3635206c69cae3d543ec198eaf21c780a6fe73a42ee754920d55a3cb778305a694585b0e4494df9553717e9f339db6fffb8806dd092c3bd542cca1c6968bb9a493197782289a6f200112fc30340894ffef65c6b34786a1d512ad20da3997682b1a7e1d4bb70e1615a6a394a871236fa1fcb6e12b24c4cb19c9e4aed74ea57103a460fb94e4f3d38c18b4d517e6b6fd550cc3041e77d0a74800f72578792b75c0de4b95f8b7f6a28b78e563cb887e039ddbb9b3bc8c6427579b809d3c8361e9f7dbdf76281d308237e76a9bc2b1c13dec9af4b5b07b0424150459d2427cbe0f1f7788849d9b08733d6aa199ad3b314864a2441ffed7dfa0b1ee91231c279796adbbd5380769a4f8c15513fe11ba0498b24daccab3393aed1d29e741736d7f2d4e9d965b9ab215f7bc89e68432c534993d644ed86dde4f27d724fda281beb0b44ebf6f8826826a34fbec59ebf84b5f9acfd9a2256f84c031cd9aa05fceaeae2ce40489ab4a3a6122656d8e9e960e4e69e40b7ed741a91112e49a150a9b64ffef9f68211a6e626fc23e7906e653b5efd3ea926f5f7ce15ca12f371b3da369bff3b56cd8de16da3059b26eb1b0cd9a9414586945999e24719c6d2e0689f3fa8525bb5f61d227db3ab89ce6ae84f7826a363e962f1b5ce7424e779664da6f61bc53e87649f1b4f1a797f83e23ab7ffcb54b009196db17775ac02c4f73ebaaa21667ad5f07bf36157c0df1f56ade74194a354cd787aa2c689b07d2dc773850aed9fc7e726af360f2ae2c3c5c94e06d414093617c23d745c353bf68fa5904398de2facdd6b8f18546563591f3f2a7d66449967b1cc4241630366e1945acc640bfa5d95092f692d76e816e594013a2c67bcfa07e4455c49143ac0a484f575526ecb5587e83ac21a4c3ee460125566e0345f587b730efcc067a096d3d692fba1e7840a80e20dc61e4440d797447ad13e3b9a8a6dd99e490e5f0c8baa649b07ad25789456ea086107230d4469a3fa066c9f52ccdced751933d00806adea48b73b81a60e5db56b80a0182c7e7e01bedac31b144e5bfa52d8b320fbd41da06e455103206ecfe04e2b57c92154f887257f2a85a8a604824629a3f0910aa8d197736cebd49cc19d17b065563f36bdc27daf19e8ed706e3966664b335357fb0124d85c93d9d9192227355ae8f4f2356693c9b4fe43bfbcb0595f9061ab43f7404771cd1711f6d27632372d5264dcd8a85a3bcca5f4af0ee1463e4d877b5078f7723ce4f365bc4ac08eab4453b37ca6e4c5cbe8ea9788c8a9f6cebb4412a3eb994055;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h97d37fd33e859de686b84e73ff07fd50a36e90e9e37b1d070141e33f4617ecc3f8ce547c2ad59839bef738e95d8e7c211dda9cc93581793f5c5cdd1c6050e9e40ee14b045813f78872f63d9cdb61d67d9316c37259aa3a5fdc64cbfc315e1ded862831bc413145396c8d96fcd519ba2472a65f8590542883344ed9da255b43450eaefc7b6461b7f661e37c0cd047fb9e6fff06f30269aaa7f712967e13078fa2e5ae3cf1ace39470ef2e5e52a74796fd1cb4f47abfc6da51d3a5e43967295e46d04352185f654e551e9506f4acca4c65de6133ac98219760d7f667d99b8af8c178c92e91938e1758a95642a66cf65dc365cf24e647cdebd601276f58c95a32419b5b62103ac11f035195d1a9e92abf7cff5acdd9db151bf6a681fa4aa03c6dd6853334ba8c94bd2e913a968e6786b8e3ddd526bf94de79abe3359be8a475c1d129e12f38ea2f96c8f9b1f1dccd55ffbe582f0e7fde6277c74aa9abbdc927aa0b8e1bee9254383cbdf7844416bd42a0aa40e9156a076c1c58d5769a0ea26d52034987475701755b9da11f59b2cb384e49658750041c319c23e318fa0b95daa969c80f43c4dc7d7041ba7de8448cde230c5fe2dfff0b68d6c292301872217bbbfd3bad1d9ae9fa2f21fd590202010bafdabb9422ad2c480301af19a876d63719d858deccf4686339d0a30e7014f7776d210c5ecf3af8fdba9faf8ddccd266256e29ef03926bb85dfc485c0c5a951b8a9d64b0d075a0e66cf0c6c74d8bdde693016249d47d399fdd7663c49b59380606e0485cfe6f809f11f13456c012d066bd8d43090c9c6befc3ff7a29ad379c9e73fa96b775671d55f0056b42ccd3e1bd60d3aec02763e54d1c9de80ff85f972f8713d11cce935c587313962e25aed10950e16315881639b083a61393d8f96b41a9ac954fbe0fe836936205970cc02656c175a4fc3d5c0c5b091c60b49065c8879565a46209f163c5b4ad599713a86de82adb75b6ffada5afda466b8ec370ecc14e155e59ba8ec8624e8fa97b0e1de898cf85aeabcda82d72e9e2904d1fc9e70b1f260ede376a7d53f9b9413041b010009cf195e3ad9f137475010c1c3ca4286d15dc0c3aa068042ef1518e341b2d5e6eeb2cefc11b048a39e3defb87fdd40b24110b625cb29b342b61dda9252e30f698c39d47cab012b5752cab1dc20fac6c8f25d0b725866abd0756b805c043e6c645b0a7c43b72ae4f6dd47dec5fb891f1183c36b82714289eab2e40b723b8f264df26bddce91446f9e090e581b2fb28282ca835f7e6b2bfacf5fe384f1f3da67c5ce6eff4f513884b1d037860df47feea2cd8cce84dd1d5ee4920a890afdee4e8f4ffd6dc427c747fcd4615d4543ac06729bc6f3eac1b0b7fd1f06e4652d2c02eac46e3b7c235f8ced24686479bee0b9ca226ca85336a54028103fdd8a7e686cc221c363b069ca2ae7aa34215caad8d6860dcd426e022190b02a0a90610ae4ed9c1fbb645f1b059e15dc88f65b535fce852042f7d1fcae72cafcf7ea958120fdb864614308d3633c36c3f081b0f3902d893e40634d60515d8a083f53fd3c0b08a6d9843e3f2be6586a9f603d1b26e5a4c185d88c028bed84130bc06aa31fab46d497a781dc226ad0e43a3640bc06326634ea805b06de87c4b7aa58b0e905c2960d6b3a40db8926091676cb592889211d943b7724a55b36c7bd61902c3d9f5c5ef2d3bce083cdecdf4225483bd1aa2be1c4e977f6d6cf8860a0db022bca82791e79579bf65da26c6c4641410ec2f477de696c06d57dca41df16641f46a1cd0c99ca61d05e95a8209a0bef9bd6cff3102e12e2d8cce0de95560f3c901bcdc67d7d932e4114304a633763880966b5e59f3b326b7ab023e86b155b75a0c817cc95ed47e637a94c10fa506a5e3173a985bc943ec73f2f682e5fbd5114b4bfa51fac8fd507c238d294ecb550b03f5ea59a24287ff4478c7f07f9138e46f9c88f4dd31ed7be694044973d75f7bbfc66621f44f2cf24171b0cb49eb6fb8f37738362c018bb3fe81aa4355b296b8fbbeb3075539bb9b9fc77c5ada6a8d90b38534dfec100f78ccd75d46c02640b920c6354604a43eed332ea72b4dae92dd06d2a6a185e600cb900dcba101432f0ffb01aeab7fa102dc3d0e789f829e224502a9b72e23ce38b62c3a7e92cfb11ee980bc7d907abf9a784392b7de3861446bac14e02c22695d9a29ac552b5918270f00b86d5f820a2a6351a2248df52ec8593bd3e69bbb83cea8b036889a20b8e0c3bc7f0a0c6ad7c0a6be06edc4dc1c35f1b0850c79848aa1c5e7b1d5120c1d1366953c41f0bbd024288a149daf85ba7e8cabe31849e9d8a558f23cd26f2627cf972a1de57ae129e88a328771f4121c9c7604c04acd8b2ee375e1704275fefc82e75b151fc5b5c05c4e5c244474e6f8752fe682679faec4f61320f2c0de4c3488d5b975af24033bbf48084c84b53e58b93cc1855de7025a0a9c7fdd8136d0233aa84d59a772452e71d6ed06e568d23f6cd2f317fcc6b0428fcd65712afde3f192ec4d826e665494e45f6728dc8243d6c84a775454ad2683094f8369095a70fa5eafe1b550593d633f5bb6bc9b4adc37a7034422c8eb7a19f3c4152687c0d8dd04ed03ba4cea4afeb0b6fc51176b8708a5f69d6324fd76e104a567d0965546c51bde135d80a46ab0ddb1b80fc0235def7ac35f5a38074c69382df1a5fab26fc93c92a65488af09e92f5d67eaf69828ca6332ab7ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'ha846e1dcc5084f48883502c120635369f4c98f557915b1afe6b33c61bd527a93b1159961bacae60201f2e0603da9816dcbf329a3dbfcc1d2a0d6b7c6baeade394c990fbfbac17abc2350ac13079f8ce0f6ff6d17e5a2cfbbc3877c9c8782e8e1b5ee57de1f846efd0288f8ef8f748119c8634a53db88cdd3c0001dc867fcfeededbd1072df84c41dc1aee3e7639b00af6ba31d8194ca6d8abc39124195671287832a562b1f462ec74a26d9e041984440da2593dfd09748b51c1a24260a0864233b957bfbc9577b591c867a049ff6a8b83dd99e1f8867347e695c67a829ba7f20dc7b53ca6fd4b29eb5556d632551ed9a42c858b55dc653fc27d21787b49ade8e955c2ed5d84dd7d92f40af5bac77cf178eeb3e2cff5b177ecc77bba2df0c53120bfdc114045034505a28737fe14c7adfcbd1c1379c4760883ded85c6ef49821df40208c79dfbe46bf5e5ca0ce10f69c2a0b8d3d40e72b7ec9a14ff4fbe1bf5ce99ba2efcc40c23ebc82426d6719d5e270762e748f56829806b18a7c235b26d1f9d0c458f4e3dd2a1f78e6c8f46d3dd2751afd60ca943363c6e05af3ab4d23653721808df8ffe4faca86b515bedd705052455fc83f286f629814409cac91517786d6d47ff6a3b704001747c6ce53642341ab574fb97d930ad95d4a8c5f11d25562d7ffa4f6df9f02745aeac698da0510369c0faccf1be334debe8d574d727bf26e610cc41e217263ba8be69c2a56caac548c11fe600bf943447132b439dc26e71a42850d88bdfca7b6fb1e80c1be6733e42e0ca6baf679df68e5f69210b3012e204a1d912bdf7392300360f3f94ec44f385a144e05d5d21ddcd01a5a7df68e1a9fb1dde9c9d3bb567a96c516dce3ecbef663aed743daf9b417982825e724a93826cde9221e86dce1cff0961fcd8535962d759c99b9acfb3485c802492a3f2ccdb8a3cfbb87b17636a390d233f88d1b057b0f78d13750d76239f371f96d1827b7e8547b545320cde9607ed8d0344f410767c0c8ca8fb8365fef16022c58c50e634a30004d02736d5eded006b02186621a3a14607f3d83df2019b3f51ebb2bcc41d84f7264035e629c4c6ae5156dabb583f3b34eb1d8bb8e5a4573dc9faa45ba1dc8183c530855767dd68cd7b2e33379caf35a7ab1934c06745befbbcd7f8b46545ad00260fa2fabd8494a12c5c7e6bf94c0e3b9f0211bf0e4d1e11e0945cf82da777bf68d1dc4c7a6019222c0bad765f18509501d05b7cc4a4fa3874b2b8661c071a9e3b638dbef31912005b3517b1242528be924c81dfa918d111e7672ea3bbd49d77ad63d5dca393e9b27b358dd07eae72e2aaa806a50e0385c96695c60da3b3f68efc4fb09d4cdc0b1f93b15169a3a76b0aab0a0a1f66d014141c6d0f21267a52afaf01297f6ef9da5762692a18a5928dc811e3a6bc0613b7d13507b7a257f2184490dfb57e40fa1537b48143d932c06440d36af66687ce47e68d357916ad6e4e5bf1e6a479eb83a2eae38145db34c70545a63810b787309ee1363286061c96992cb3fdab7d9ad2d0096a7bb6ed1ca2463d496908ae8a706b1738f6fa731191ca2156facebc2b6f535f241c00355b5e9f2a5996d8eabf9710df0a0d3bc67ea70855e9f3022ee87c2016d0688735b145981ce6bf027fe4984f011e3d23b9dde37dd78b90ec0a604624c2366f37963d73c6835f4223fdb9884ee5779c3df4bc5a733b9e6268ded4929447145a0665dbd4ba766d0dbeb30b5154e10532d82a4e65458a806a37adc748b0dc98ab76158b5e300a4c7aefdae6c140ab3edbdcd84e38f959135c40d430a1b77c23feaaf9eabdc0c3c217d5d81b2b669c58b94f28875348822fab2cdc271f604b43b0dbc4d168cf723be3a2e6d2a1a3c4bc4f95d98972da58a6a7b07353fd99253f3311dc3ed6297e01e811594483687898992494d877b6f257a8bf1ca8955407f61012bd26c99a121d263f3b33d1ab44861d87cd0c6e387d52650b10f0391d40a7c52516e660cb5e421e3beba513e73a6fce114232d5218ce492099976b5129163cff7f372771abb60139d403fc58b4aabfe8d40f25fe20e6b0306e8c73390ac1b58f4424e6c637148dccf37c2d4bb3d6aeda8874094460fb66085f24e6fec9f63b8dc38102d917535a111144afa0f3850d145ae26a5d030079e18dacb9e1b0d3f4580df548bd5e75a8e3d8fb00edabacbd3882bc6fd91c2beabc084bd3d882aabdc756bc8bc3ce4c9e1af8c0791b2154bcd34664a621ffbe3d594d6fcae43f3d944f987b41d9e858c6890818c3bb24165bfb6f5783781b7ef3caae24d901b9e8d9a3c0266608c2c774a9a099d506f484c2ae091689823a28a1e3f314982acc14d8e7480640e221a0b2fd474ac28849789ea07ed87b439cdd78640476f547ab404651956898cb8ae2ae84e39ec8bf127c7c3b90831a1e84f9565cf7e468456e8a539880f9da99eb9a7f236f653892a94e324d587607be82a46d850275037bbbb4f01afd981a75c0d311fc5f76d1b815b9fbc520cb86775896a10cfa9c06950e5ec1f72164bfce709e11a2ef666f53fcb52d06e83d76b74189f43fa38a93d4bd9303039daeb65e4c2be611d007748f38871a24502911ff8e4a873ba425421842e4eb0c62aac6978def44d441c1fc9c669b9752e1f12f5787cfda11325b052429f76fae9a152ed9bc39935278bd8ecffb10053177c10dfed6e0af9960cc7843264f1168308e367f7dcc87cb1897381;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb98ff671c7265b84ba0376afae9cb9b262276397d26bed004290f547e2cb5d401316be8828f19895c8adf512933e893011c383d09887cb1550dbf179b78c561ce141e4020f708ad6eefdf9de1953b74ff212609dd25d698dad2e9c13604a242a5044ec53acb4f7e009725cd8489f5dd63a5f4606ee3f317e4892c0ff8d60137fec4094a6c2d78e4aab0195cdb93f1cd68e916bf686d771fe8ced0c316dd2f46a5f30553f41766c970e8b14eada2cbeec1cf5426ac20f8572e7156a3b1c215fdc49ff9c4414a665c06c43ded44d179f238eab54a2ff0b255f1565b3bf1b928c9f45e886dbb98ad704dcfc878ef1e3b29a92faa73c5236ee591c0624c10408300272ac4ebdf80184f8d9d08e8402849ed921955d6c88937245757caa7e5a4506eb9069d3f69b55564e1b6a01252211e4cf4809476f9b5cd1b05d6d73dcc06ce300754fb8cc236964faee3ce0d15154102e35843aec129b270b967f77ae773c5c65295e924e7ed3d6b7c9954a79f7925b67fef88c6d8be1a7eab2e93b3694b35e829fcf0a8dbc7e6107bc1f776cd710bd8220d6c6d8a24e54bc7dc629bbbd23ccbbd0155f13ee5e3d7c914fb2cb8279cb2bda908cf5e7ff84c114061de873cbee78beb0437d533e34794849ef7e8c7914fed77933d79596d410700cbd40c1ed3a729dfdaf42c29fa8eb0fb04fd3133c858028a78cd80ae26c3b2a18766ac3e264f7d83b2a789e18ca5d503d66c5948de2b55b6482e63515a2e40ce4a48dcf56ea6ffa9f1fd8fd52eceb86d0da3edd52e71a85feea991480e05ef02c38926b5288b32ae09363d0a124b6458f80c480926c7dd7aae6ca235649fdf2107b1260939e0e41068253b41c6064da22edcb9a002b9f3e31c674f303715085f1269b9ced8cbce278eb9eb621f5bbcdebf70ecf788159565f78eb1bbff52ad5d7c916f080db7d3ccfff886930dee07a3b761372b8adf3e2c542d3609f79a7b7e6c73b2315abccd7b4c7045a076f574df07bc2c9f52c2f1cae4f8add905c93b6786880678943a24a5a50969cfabbb27f8f590a077535bafb9bc51d515185b66c26e72ab624f46d43d8f0c818372dd854a4d7ad27fdde9a580e90488ef4135b398d0114332a0094591a29ca9b29c05ba244204655ebe66f6642b96198988460ade52e44aaaae51ebeef04acc4acd45a6601cdc687284a231b8d264f79a7b95a18520dbc15c902ebc6788aeb722ce7e141857ec502032987b68c5aab574e16c3ca50532f06f822843ef202ad85a1fb2407076548c8f5a246a7d543b7d74439472e0127ffde093535dd291c0769c7a200a61a4de3bdafa0f21058dd5956ef4cd2eb60d7c344ac91063e5159656a1a2d7ad45c1911b234e17b3cc2b2275614a7ff926924f8fa54f138ca6aad15ed971aebe8c9058212c4fdf891eb23745c363e5f856184926b47486fb10b65c7a2315a4792704f68dd3999a3283896af6e1fba7de52ffa23529c10ab32d4640786a0a64f49534a0c76a9451ab5c2c8b9bcfc1742840ed90110bb406cf18eb4d49b8a7f1246a6b6a4ade662036d18c8f64093ed416dd8e84d0a6ddf8b856cd841236b4caecc82e182fb06579e914317617d1e82c8af9fc34412fb549d2c9ac2d7a3bfc8752668193644d9e588ae02123c41b37d5252f75a747eea858be96bb70815b103b9e19288e3aab2aa278553829b06a20aa409e128d81b8fbcc8a9d685ca6c51c81be036f21a76454f111d9ee477677fe760c4663e0062ebf88df7494b8247ebbe9c8d55ab3914aaf2d165f9a5c69935e982496ab47d2455ce370c62ee34549e56b34047ae81c493d4c5dd890b08c9ddebb9970922a07f9c5b4b9266b7e3bdc436c11b01202bbd4c88fab06c864d79251dea3157b41764125ef849a2fdf4cd99aa72b2b8f534ec35e2899a689dff3bc764e38ac5d2926526d70179f795d6a08a19d83c75e9d09b8ed439649bfef8892512d9d602fd1d12f9fbf21bb1d5cdbceff9f8ed068b52433534cae7aee577d9399890665bd5d1abf61536a16cf67da4ec66caa48a8bd339c3dd1df4dd17ce76da75403c38238cac8b75379d29b2d932e460b0d46f84f31fa4308b2fcd270dd657f9debcc6ba017437314a6ba05656edb9f765423a6e4649f8d956cd43c2c19382aad5f51d0d558aac7246f9d5a026e0c13120868fd4abef85ee9a03287112d1c24f22b7d177f1f6fcdf327b34487379a479581303d3ce6e54d63189cc88cdc2c0b048843e997dc8520dbe6e63f5267041ab1e1dc3a18e10d9fe5b7f1c5ec95f830010eeb3fa539f3753507505a0a43b1c15a8a5b60e2accbca72a77adb42d8abc9e5f9461d1be931b0feed13d528a2f3d92e3c2b4a745a7ec4289d75b00172df4d9e1ca9c070751ff6ea2d6397c64aa32422426e5d2e5e40a62d6b2a22d893b0f0360532ff2ce1012eceeb29eee82e50fa9b48194d3f86801091db246dec9093996898b3fc1952f765e2068ed06c77674a41abb08fad557101c0c74b182783bbfe008ea2b0d5f790494242e318528695d50ec3e6fe3ea52b5a6cd43116421c3984a5307f67683a13dfc135ccb12aedb0f172a3bc805027319ab02833c2ef30a1205985e8429cf1d67a35fb3473c3de3ae7f61a2c7c5cfec96e6e5bdba9e925f73471ccee750579e456f78e57e74f35c2f8e6f96ed553860912fab6befe0e8993ce4bcce065d960befefcee54ab6f6989b8012a98f9766312c1c631bcba2feabba7071;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hddc4fc0f25d14d5e300049559f7d95bf5889d91d9ba014cb630ea70ad11a52ddc7e048a4a2558fab98ec80926524bda38f55e167ceb6e6b00f13837946d1cfa59d307bdf4652240ce94d3961579086590d2475973800b8afb59ac3b95cc601d2d3e8ec5d07435a090b9094691cb6a84aebf331f91e5679b92919a5fa08d6e81351691a1501afebf0246f7b6d229b3ddeade0bec09636548c9e1321f88e894c3339d11b8dd72d27ea43136c4aee9dda08e462d2b094fd4d16eaac11ae090f384fb75e1c6a9cbde411e94f6a156e67a9d8614fd5e1d945781b768e46b73dea4b6d01ecfdaca1fdda373f8f0a6b514c7fbcefb77a9eff228adf871dcd19dd129bd700f416362c96ee02ca68869667f03d30bacec9ae32cd99598f7a49f016e81ce45f6fe44097dd04d0f0d260fe22d1022ca2dd6e3870935554837a30b18334fb74670fc040d0e4059dd9d4f3348729dfe7d8f0bdacaa14231ebe1835d230cc2db0a190d4aec2252d75a4dd87067d43e86a68f8ce530a689054d846af8e6d2a18a0bf8585ac1260bce863963aa85c882ae935915df84aedf779407211755d18b747bd0f43a8fb998a0a9e29d8f27ba5ca1aef0085bddce4bd764e9ce9c3bbcd092acebb34b5406c9d0a076e36d3872f31f3c1386de82e6752ef3393533689454b7da8035b7557ed2208d5ee9c0df4df7052e3a3f99401fd20546f7253551886161a033d5602ad06b3795ab9333c58a260717355f0ece55c9e9c37ff785f72ec7e130a05508677a934d26186ea3c9150673960937c452f944809d7010b49523a01ac33d446262d0a624937642289f06e84d83a00f8aa2ce873ba25739c9739124fb4dac588e5ae9bb3c746a0ce5694845c816543190ffd6e464b40e21410831b545faa67c202ae9a7cefce5768aabeeaf39a8e57925df745692a9ef1fdf078446fe3b80d6a8d4f3320bc3923c4ac63e651238fb63924eaaee6544d721775c66b0b738da17b9aa51c8c5c4cf1bdabcb0aef7f7e77f3bb32f345cefe7a7cb7fa3cc4a610a16d1ef4bec8f1509e91f5d5a180065a52f87f076d006834b81c4320ddf603cbb0671dedb334e0cf35a9d4ab60065940188e56d31b0e401edf57691263730a57f99c05c1bbaed34bdb1609fdc557093ec804779fa868cbb54a1af9b76f8df488360d6ce790e9484cfb41e2414cc82439c963cf3d36cad0b2eeeca43ce155a0f9db67e706a253adff22c00f1d51fe870115aa439437950e5656f76b6e804a2f6b40a81d23b2045cb1b89c1ebcc9dc7ad63280f077b590b400ba1ea0d822300de49d243bcf348a08784208783ede6ec6a1eff7c3cdea14c07feba97c9230c7ae431278042ae91905717809da7c570e0fa01e43eefbb620bebccfdfc1fa32d0aea62f5dec239ce942b8fbacdebc730b728f3db8cf194fbaad89dc00dae743d96bf618eb08fd878365f92407c86d4534ca88a957ae6f5a0de7866dec445cd0273db34658592fb59d39c9ac3977d61341491ec9dcf80713b1dc56296f8c941837f7e1dded2cea5aa3d5194654342a7ccf6be8cc43025e30fcfef8842f93c2c38976d9b5c856587f1bda0afb535bd1ea617b21deefdc6a4b8a11ad93d27937d7ea2afd21abacb1843ac436df67c294c24dfd691e0868952580ee67a8a1ec33f47291b8e0fb71ed9dbe9760320b880650d70df838c4985dabb0033be8bc9f09bd28ffdf2b14aa937e8c2dd663fce4cf9b1fd6a417e8ddf33567de6bfb1190bfa6dffd0ea09af298db9536326ba54db3e867b1a4511d876bee06ce074d0214ff404e1c592272040b1930a650439b61330a42694eaa9eebda85cad78d4e485d6f418362f08fd85ce533ff2101e01c66468c1f3901b60736ae4cc368cef8fc36f2016cff758ad2902177bfc135fc04308f452acdb0c9852d24ab18b3d3f0fd6980936acc1c25cb1f907bd9a92a03e7736da25ad6c58daf35576e211e74d74b2f9e2a75affab167b3e155c968b7c13ecd3ca694745017960ef686a01fe6d0cfb5a2b3337890aa77d65395c88d2061d8119e9ae97317ca7c32d4fb20ec2e7d30cfc88486d1fe7efb81888909f63132b3e61a1c7459c8b531556f7aa0163a2af7268c3d20fd593bb48080f19c2f32a7cd88998175c54d178aa056adeb03afad8594c8f543bc9bf771bbb4239e04574fd55be734437ffe67fefae4573ba9ba73b23957a8f14cea00ffb42fa4b9bc7e719bbb41294edb9e729cab1bdf8cd8cfecf36178c53170c4ce1f53e2408a3c3dfbe84c4e863132f70a16ea957856ffe483c3a03a0ac5b1ada5017546362877f1f1b80dfc2369a841c3742d86b48a7ed1702b824843af0724574088537cde8321ad284006f8943b6ff8a1e3d5dd24dba759cb8a8841fcebd8e9c5ad949eb9587750e1f1d9a7ad5cbecfedcdb0c1208269dcffcdfe58c5e8c895cc8d3948e92866d11bf6530fb6b7f8b65fb5f8475ba2b0d06ce750d62aaede0f9b1fa5ef5d2395a6d157fabc33a7fb9a420bfeca69f50f0d9c9a754dfc1ba8f478d1d407d555d891288e7d85cb3fcbfa45f67571e0148d8940dcaf7a179e25a05883c1d4183a5de09b371c45940465d363bcb0e59aa5504c3653cfe192f6d5bc1179ecb35e7b6cf85fffb6ad4eb4ca5fe7edd0cf2ed37c9923a8c4bc3307b7c059f9c9055e3af155e341bc2475ce24f22811030438a54b42758ad71a3763d478e0c96fa0604e78b35bd8b77828c6c6c60724c354a353;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h65e1d4b1683787b2df38002c9bb16278b16b2816fc3c1e8c23afb8a8071b2b42599e2352fb252829b63175de92dc955792cbab4cffd9c03aefb0a4d298afd78794342d649e7a7775c6f9914758686677a73795da79a2cc2add8e1ea82693229f2e0b1ed6469db85a9c3dc32586a36c05bf7bb85ccb3b48f0dc648a08aed2b674e68f7408d280df745048b5d4733098704f7c5b7bec7b5de792b84c8fcc0f63aea00bcbe96a1d08020571d030daaabb947e074da1dcb848e284e6dd8d4de338e98d678703585917cde2d53a6d1ca4280a8f2ab1c072f592bd175b67e80bd273ad4ac0ac20c2dea3d16938490dbf049e2b937df664333bd24a086c922794d8d7d8c300e20170a92cc4b6b1f3519139e05929870b047e7612a15cab1a0348eaa979062acdd1d9ef361855bdb070adce32afedc33acc6ef424d5a79b7f658a4b220d669f58ee5df809b709c420c6fe017c03fe18f9e09268d4d61b15e15a9a85b3679363020ff771449e658f01b7a97a5a2d9fc7458084f3a29620aa63541d1ebe3cc9d32ceaf12eaa86a3cff5e7733a30531c183111d054bbde7bea63f16ac1aee6ab4736e9e6a5b81097120f18e295c2ec4ba5a998073866ec4af415c9c39b20db5783710976388449bf1f3768d6591c4d2526a7bf45e9463e86ffb12840992915e03915c67b3e230d7cf9a34826471b64db07f2b03dd1f82779cbba4447da092e987a12f62eb1d7c62a3e0d09c8a7753b75a6f1e1d453add9ead0ec29d295fe82edebaec60524ea59713f3bb6f03469f9648cb2e83c2b49029713c7eb83ec1ef8a5fed737025f3a237504bb0767b8763a7bdf8c32ed9cd1662d8410d2105c065258caf92d32ce33a5d907212c11d5b9f69dfe7096b0dcb4e73e6619be71a8efd989574d6a7ddbbaefe80dc8b56a04b7594815012e0b694bf2445c0d0a0a7abb8558c66a426b7073d3175f9467f46d197d5ad62ae921ac8d77280a063b4790589dfd561c976e3b40d39e132d577b7ac85fead61f6f705eec546355e46ea04ede86afb7687af4dd4a3904b743544f4c6e7136686e514effc46e4573a97aba789953cb73437e9b9e847a3bab61fcb59e14611147f8a3256eb9eac06b3d1a03495ccd88d54e01aaecd2889f59d2420bdc04d0559f7afd32e964ef46b701be7767ba79407a46b38ca71056e5ef664884338a9164b276764ae271fdb19173956e40be239484ce270725ae616406e2c701c86919bbe564240d67ede1fbe8f0fc4422786534420ca5a5ac9d79c6b0dd81c93da20c437a80b401c1aeb53c1813646d3540383f48a3eee89ac0288cce4ba6da02321c576a577f9f8d3c196e29e6cb96bbd9c54a1824436c56cb47d6154d982d71c91fc28d94380fe6b17f7a083a3f8a4b2b6aad8b81a810e0f2aea8aabf1d20e6ede056c732e1a64ed8af5a6c3d269ac819d454720cd6992f677ce194e1dc42770bb8d79d1b8b07527c6087b22074e99abaaf2e64cb96a3916a91ed98eeffedb5487f6a70eb1d6c4e18f4612763a00bcfaf40ec1fbcf29a5393f4efd74530c2f7b8b57e5cc46a09d1e38c531db8d334d9f0892cb89c7e1c81c1a1538b97a1412cd86304b4748d8f9499eae7969e0fc2c86c68874543969de62aaa610d35e406ba4b527a64392066268d82eecd579859c843b540a852c6d379bfabcfa4717d64abba8115b9911228653368bb90b38acf18c9e492fa3c583a011dcc3a8a5238edcc92b272bfdf6def11e21981f7cbd78c66e4b5ed1ce683e4f3925cceb4cf6c5f55ac6d731e4fdd3d7753b168b116b2977b401190171543b40c68ba0b014cb0260d09da1e2049ae38f115550bd9629383f6407f9d55d7c308ce85fbdda1ba2fcf6c2b836c2b8be58f9f62f996e5c6b4048f02aff63d6144c15ff3da9be79c1cedca09214aefb2ee6ff2fa23e13e4f6a3c0df93c72067d73f0af61e3947b35f9e4e38b7e75c92afbc0de0588bb8bef1a09edc881dee8e7b187a236f136a22d341f7929721ee9f0f35178861fa017c431d6b86403de76735c6200a7d780b5ff323369070bf76c3fe334153a8e1a0f4c8dc2731ec618dabc4e66ba4a91bfc169d91242290584c3cc26305f8eaa2fcd2ee7ad7757c422e6ff7003e2828583f551dec4dcf8133f2d32cfbe7865c00f079b645137b63ac5073282be46b17cad49fed77e076a5a0a96cc8d54325a31c6af2636fb4e7533fa9b09330f917f8b169a0df553dba1359e8ef31cd0d91c38a6b1429b58c66bc8ac78674be53ce941c1fe040cacf7c59b20611f8c26e9824232535a398a0d4c99aba12cb8b10dd592ecc7844252bf741e7759ebe8efb717256cac9c55fa8f6b880b55e3f66c07d720b419af5bdb4e5dc788318fae6f147f5cc7ae2b2085df7fa1a11ef04b6f8ac46fdb9b2a4fddd6403856c2534dc06365a23b71c9754f1b185a9710811d5850278db98c14b7e28858cd79459e35afaf0ba8299039efb2844c19de6b8ab431b129594d4b63fadd93152d9daa1d1c48f30d24762c4c0eed89453305fbcc9986a0b4eea8c4bbb6ef25bbcb6bcb8d9d91a8000331703b7cc3aa3929454041fc9d20f28260fcf07bfa1d207d59e90c9eac8574e16ffec6c55f3488d47235ffda99bfcef85146c00acfc3309b4bc7ed230279251ac18812b36612fde42fb26e3eaea9e5e82b9e2ed6713e99ef21586646918d7110dd12c3444614aea4d4d8685402d6ec1ac3c2810c914f1203755fe5434cd5215f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h827a9cf781625e36ef5ce5a329383f77fe8197d863b8c4b7d7b364fededd1f232dcfd0acad53c96fe0defbd8b5ce8bc24050337c45085a1cbbe96142430518e4f61e75b6328ae74cfd51556eddc5d35584c3eb35d5a85167d468122ce88cfa5d980acd6b09f728a84d158781f13e1d953df5a7fb28775e7b061eafaec2348ba2846e5cba891f081fb02380e860c7a972b88003266034ddec4c407148cd4afd14ee6f7be4e0093b1316a03b1d178494a5e78488a834d85d01112a74fa24974b680a62ab2774da19c71853b8ae3d9932b87fabccf76b8154472259c117f282eba3bafaa55e4403ee0be1b680ded004908d04ce148c6574b7c1314d4b22e0e088f26ac5768d0d4b201e74fcaf7c10c0f1f8e3238ff7f11466ee8bf0b4408c62d8835b866dad670ec76528237b35ecd0f69a0f43f19fea21bf5d1f83744e9c1880b6108bbad40462cf641c6ec12f66c3ebd6bba33a8dd5ae16476543eaf00e7df01d7d3336479d66753748fe2132e066c02b9f6692a765170c8a43adc2bb32b42949712306450c711928d619eb82e09336c39a0e34036bdfbbcdc6d796abe15bad67e5fe716b2cd830ad44e77bd67f856e37757db83e2a4be0cd3a640c07165b95b1b9c43492ef10174e18dae9dde18d9331d74953603a2b5e0acac9e5f7234e8c81056d67d062bedf60d687edcaf91ba9f27abd0d9c727187a2d2938428adee0458506e66f8419ea3521e646535893035dc4162b8a2ee91cb9f8503102b8e967b0b75adfa5e4538800815f1e7f97f1aef1fd5dd0040f0d47574e57b406f3402bdf5878bf5d1dc92e25aef1f71cee9385d44bd13e49516882e3facacc855afc25ab03c87877a82946952a7dfa4b1bf9bf77d05befae187e53e401017c9386708d522e1d4cb4ebe62fb4ab255bfc23146b403c205a358bb0c83e3f405f875f7a6f2bb9ca8c52a26010d87c1c2a56f96484f8411a195633daf6458fa645c67472210512597779485dde52aaecf17ad911fe15f5a423f62ac09c7959c5b5955368a4c488b1ee0914d0378c152068609735aed5ee12355d4103ebd41f3b3a30190bc01afd78d0d559096ca8bf11e122a258ebad6e82c2e20cdb03c1bb42e3f49e7f4646abb098bfbcf271784786c82d1ef757351e96d821fe52e84a3d1ef241c0d41daa9501930ceb05044767eeccd7f8d85b110c0aba68302ee54c98e4fb4746db089373507e067bb08af37c742afd60c55864f7be10cd898fa7cad3319006b6daf59b7971e2d644d32cae471024c6655120ef347598b79a16f3993849896ac411a68522a3575d0b94c72df3deecd673e8abb59da5cb1bf9b35a781673dfd940aa92ca96de4056765dac29e94321d4bcc03bc37152ab4afc3d47d703f6575fc0e136f7c7947d77dda823345fc04ca66cbf1d683a40940124ac987e4f7223efe8338bc548dd99b8489b07242436046f3545cbf062e73a1ca9e182fbef527d2f08464073114cfc75c1ed34fb0568c8319713c3d512d93d09bf8d0446140363f00341bda2289173a937fde9dda51bafd60fe4c72279c720ca3781be8899ac2987669707d2d4df5373b19031a52b42825e6a7a3725991418f557f238039589f3ae1a03c2a0040d03ff922fa894f9d94c92962b0cf8a6eccbd6fc5551cdc8477fe06a0024c7257f81b7617e8eac61c41475b529d98b4b917c1d5c085570c6ed993dfb55b697d6bd1dfc316ea50e53deb639a1c2558b538ea7f924ca6d97efcfa5464f96e9a1070043138dbc4a3d21ae7b8cdbd209e9004dc0dd0b185403a7717c85f5fac276924fcdad22c741ab5fa29cb94f0a87d399a58956c88c1cd3e24b8f5cedb9dd93cdd67671ec0e919c438e45dfd14d347022d90991f76e2ee192555a9620c7770f1e269aa06d84d2b93c35f8d4579d3e172bb255c8816ed18427df547cab131581f7f2eaf9c8cd8acedd961f4393b31c16be373e7013fcc224d962c83a42aef42f7f0e021955c69161342a36faf073d32ebf6ccc7b58bbc6ecfc6b6db3474dd58040fc87eb3eab53b3b25bfcbd8fc2746864626d73634a9418d0bcb362fd7e43070c538f4f3fe4540e3163906643ffbc46512c232ce16b52b8c2603d7d7ecf677751a3951d49320398a2a57b4713e6c0723e681227e55a592757261dc7daa375bd6cc99931394aca38a8d0a41c8f63e038b1276bdfc2c3d495bbedb0ef1c5fc759867b7817cfb3939c4f1c753fba4b12b961000d8a15a698948c6ac5f1db9a1fb4bd8af31ffffca1510b39827a93f126ed7040648ec35188a31ef3c9a42551151bb91868ac9be7cf213b4515a90a4d42240b1312951b407d1f852d7841887f7b7bbcacbab41f2562a0a8ca71668006ae567be61f2d2b6bdb4a1dd369cd4c1f8f5e23ea2e5d0d775b7596995727d37f2c329638e4961b11474bd0f4466b45da74a47df9d7a69e06eafe7f1bde600f2618160e5ad8fed80afb615538a9b79adf0b31874f3cb184691cff68897bcca9f1b8225e7da0286b939504f3145e21415bd9caba87609ee013a22b061c23b3adf02d80add4dc4904437cb64e580f37f107446e7410dda8ea4dbef72b2edd702f6fe03dec54bfcc8650e500b1c04e07033c238d37f0087db7349fa4a45ac85643098ecd5bd9688f37c88f7340e56a1305c20ac26d0b7490756fa7fc0dde26232a62c3186c82261db642692a5140e0f518c6ff0569457fa9da2d8e50e38a21a0b8a3944f61a33d15501fb66bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbe9f78f54e9855b3e6b4fe8b90483d40b4b8929e8f6e7183f81d0687e9b0fcd4643e474f76831bd134e8470052ff50672ac4883e74b1d4c4d8059a75aab4d4df84d40e5093360445683df36a17cf83855c0ac4f5153a77abed7199ddaaeb3b61830b8df7473b19b0250030dd21724c0f388896d04c07d101ea5793af93fca27ce3fcad9edc394eb4a88315210416f521ea2825a775ed4ff98a670a87f4195cffafedf41ef02b98446b958863917a50bb6073bc22f2cd464de0daf34f17d21db28f95f2d806a05bd7148465b7ae094d23e176005d1f0b8590a93cd67b02c5bfa738ad70706ac81129304950ff09dd46ecac16fa8dc3025e48950388c554d0b5530e75a10df74bab54d540a4d88886953ce5c5774e3120c0fdcbb07000934b22c16d58d588200d4b4742cc8d5f8655e955ab8a2d80d5ef50996600202df306e72b8135826b6f80ee5dc10ee571b89cc0d2d833e269eb68583eb546c01f990a3a88983b2fb09988d53e97ea2e16e6e05496a5bd5489adc3e74402b4675610a01e86138f8cfe312bed7d9a1c1561bbcc00bc3668145e796e500f08d19c775dc68882b1cfb1de72ff444c37605a5fd9e86047a82827487184aaf0aaadc6da239a5e58d50d1223cb86aa8cf0160895c4a5fc0299d069351d0b03c8d70f856194974bd0e15851580837b53daf8bf9b8352a9cbaee52b5a9d5b00b112bfec7dd54625b164d99a81abaafc1a527449cd99af419f45dd7de7707cba8689e869dbd80150579600a5bee3fd07419ab492651eb308a2f5c5302a96ef3a1a6848969a205e54d69c41b0c00e83d068d0e858331edbd1908930131b307177d7156f918487d64074d9c604ead83d6ea59ef4ba0f355ca04a3624ad214ff7afa83614efc0a84540537f3b539d86ebb29a6d6a00a2857ea34894ae83fd781990f01ae4e966a2b436f3871806a855f62e164d69379c8f19bcdb57207af6852b670159529b84a6b3c7e4aa76baa76b2491df0b9a150fa1a61f9d871d4cacd568699e7811bdcf7b5d0d6be9a4f82f8529b326b2a796c3188757eacb873aada781f2730396b70e44076b9c6c7bf4857d7fcb16c53f676192d6e19f64996586eca5cfd66c8ef00c60158a97396d3eb76ec5ba52b80dae0b0288f71f9551526d7d52769daa23a2bf41357dc8aa6a2ea207d27cefa4492ba06a61f00e929f226288cae48eeb989d40196c6ea2d20b6832973939723cb8c3a57d1e8561d1acef43eaa66e67ab53c9bceb534babef203692bae5d3406aa3ca3b605f31dbdc4656e2fcac2d0ddac595e68a703612b6599ca97d9b90b7fe53cbacd09804fb0a73f188110e5cb479d3b10932544ef3ffd45737e382e8e4065525acf5161cbd004948ddf05397f08b44396a2771ed27735e6bc0050dd3d68d46d7ab099859e09c0ce66a4455f94a1ed3737b7e5863c3fc7343814a9683cdaec4e5bf0f790d985f1ff334f7d9f0f290265c4367f1f7de6d1fcbfa4a7300d2de42c1c7e050fa8d7bae05d98273d00c6ad49f93bd63b2c80570949fe15a294b99fe0b28217e7a06f370c7775d180e8fbea2444ec3f40e41ec868682656f9aa754b3c0a504f14dc45a9407f1c895550ce629f48a6e4cf1f278c8537d246d4a591975deebbc25af9936adefa1e9eb31d881088e33045509249742df74ab89edd38aff59d5228fbb3cd3b77612864bbdca03134e4bc9857e263e7dbbfe4f47943c9323d7fc1dfd2ff880c01eb07b14cb7e2fa4593008f54a3e934e34655c67e868e59ef4b967dc9cf145f9be06ebfb205930519f93ac052896555c421a1033f89389525d3a4b79a6f15c6310ab43ec18d11354d65a1d1f1f3651cd5d8c795b4a88a57c03dc2d67aa2bc4007884f7ea265cc5a1eeae1d43439fde455e8060783ac8ae03de4cdca15b873dc6ef4c405eae3d024300bd80c5d6997789550cd4c53efadc35534ed1c7d5ba19db6b1cacf73e253fda50a986e8c5535e22ddba3866c826c36cf8de04f17704e34554719e2c91f2e4e2f79cd9b5e8aa3043b75b7130ec81928a18dc6387ef418d086279a43f0fc319ca609597e8552039b27665474a4ee03d15937be0d3f68a35fe574bbccaa8ecc274d1f65980552f97d9f2522e84d900615b4e8f7d82b191946b012f10e2d2bc5d0e307fa913988a630f21fe5fc04855c80892ab960e4ef018b702a4ad1c09b157ed2dc0e38e5b09c654d39abbf8fbb273026e334a405d0bf3bdaa725235b1f83d8ae052691dac74b2e023fd34b8aeecf417b163e3277f5edaadb3985e27d84378f7225393fd9c6fddd0a39e9e4c39e85f9e1283ac8b773b924994f3fac10f2a47afad30f1003a5bb14048a31ac3d13c1b679f221e2cdd8e8eb68827ff4a5072f9d454c2eaebdc110772a36e20330cfea73ca7521e4f21bb0ded89202f13493cbfb95fb3c211067fff377b2f20ab7a04c65149abae057433fd30df65d26027bd2a2437aa460dc8ecd86a8e479807175e14c2a69b078edd2a92abf61ac9116f2b2f9778ca82ddb8578013537f7236e1a1f281e53ad6a7ad49c56e53a2afb3e5b6dea840e2ee7ab08436b72826b14862a38164edab52010f46b84cdff1bedc794cf22a3e475430cf27b55a56547d7ddd8c11aadd6e18b0d91c1e46b3239ca75423d37f62f604fa3677d4dceebbb69fd8db6ac5efd83270890a8cf8b51ada797a2c2108e770043d8b7d88e5c124b448bfcbb649ef2835ef60325b3bcf96a13d0661b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf581b93452e630e71c6f9b6af6d3e6178603f3301f0077d5a343c927f609b9970eee68e169e7a11d2a6f07095bfbcb54cfe2189b9f5c1da661d469be32b0d173dd29f4c2a6f89a11f7961030f0bb660edc10122a4198f5ffbc6333c399e8d8fbc92601720b700e7067018d594dfe07b5eadfaa51db1b463eaae00e8a8c58b0e0e890b158c4f02ca02ea9113c6ac9990ca3b8ba00d11373980b7ac18503351717323d249e759c156a16b5f734a9cec2e2de85b960e30cc32afc3bb502d70a96ea7f2240eaaebf3307e7dfb2761e173e54c9b97af47b0b87e9fe1f48912b281d3547518218b9d1f86a845307483c8b3222332ed1e48ec0c7607fa0925d8a5b8e4b9ca07e82277a93aa54b46338871d13facf24893325b1a1b73fb04df11b770d174083476160fb2ae62ae37c33c28880ccc0143f6d8fa4dec6457484b845ba25a12e1708ff4b0626fc273e14bd3ff2ddb8d32386ae0f87208e2a243681efdb1f366b1ac47b161265114012d4b53c8337ea1dbee41c1e5e448d232ca56d0d8038258e3611029713392a9845ba4713895123b6e2ef4c3e96c7e5bc3f6698692dcd57173f73f999a2c10185b6a638438fd8b867de2e0668b20be92162a7543c962dae0278508f1b40a0239c712c21cce907c7d9f815a94c962f51e6a3aee31448dee2dd7e0670305e5c09a118767336df1c87d523911f32173d640fcb4c902e71ca084e8b31518292d9eed33090fc34f829b3e8989c84db92e14cf26ee271391c5ec1d036bc9d151431e07fe9d3e405963ffd764293f42983e476b870afbc4fa462f185f37322ddcd862a064836f390ece9f6d5ee9b25df22b9c4cf24762231f1d0cb41d032a057aa8ba4d76a71bb95f80ace9ecd8b3173b5a28732abbc0ac9b970942038ad7f383eb06195ee8bace76b119d15158a29d1cbd85f276b3027496306b85463ff59e351413607952d614dcda8e8e2a23a9f86408dfab5b8b2af27b56210c03b62492cbebd7cc186c941f346d5e1d798a784f87e53a32524b7acd1688eb827d6fa74a14c38736f4fa5b5c4446eb128f7df78af5646aae97003aca2be2ee1bc7cf3999d709735d23ddc1e3c72ee203b1f7559feaf2b8fc3da0e18c1ecfcc649f96bad7bed6adc55fc1b0fda2f0ca724792f92624f06452b09939a70d2f554f140c89f0ee3a87bc93fa4fbb923c7da5dbb4d04e8d3bd18202bc0733e9f2323c736a4576a330b3bc69727efdb87e7301230fec7cc964b7baf25fa38f8c8bae98143f28f5be869888d87b8d32b3b4076f4d5339a8cdb394ec5c4fcd411a0dc0736ca6bd66cb123e4614a54c5b373e9daa50d3582cde9d01d82c196e495f1e04e556860751b5fa4c80146edace1252622a3c716497eee69cef1b7dc8ecc6f4b22162a4d52f1df922ee8b67063014c7efa47c109b94ca553e340dd04fdc5d651dc7fb9f990b4efd99cb97e7d464dd20c098fd0b86f73c5bbcafe1080f3f2253db8e0e1100771fd8cee9b1640c31d04a9443d42ab9e7c22e20258df8e5ea66984fb33ed637fb085246440ae0c279095a192e27a041f83cbdd0b2a8abc44d3dbfaa809bcb6dc32bbc23e3ec485ff7752cf9ac8d9bf2173580d2d5410d52ee2746442b43315fec53a32feeac3fd6289506f941c9c6c8a682a8a7eb6eab104d1f03368f50bdd180602ecf95ee021828598c842f96e84d92610db3c6922d68dcaef7c983fd9955d483792f42f07e0bf552cd625ce980c4d08c049c463006f0504a3503f0a7ddc790eb363efd1af321449204c9221a379bdd2693c9e003a739f489db3c0ef6a1f992e109579edb6d3ef9519852d5eeb422cf354c08059d5a8ec4535de78adb0ae778a33fce5abb9036cd44a1a9fcafbe896ecded5ec4380a0f7e6bb581d31c9eaf0ba3a4ba347e4b4f9f2677a35f623d781c16f56a999928ee5208d3fba1236c5eb3cde59c10101b239202d56f9f371d4c857483a57fd1decef36aa2bc9481bb711388bfc541853710fb879ffacfddf853a68d7193962f28f3103e51f97678785ff6e617792f85a117a5b6686a0a8817358eeea76a35e6ec23b87c69c6c9d99cf5c8f154b92567b5173387b461a14141b5d2c2fccecc5fa8ee1155bfedb804eb68c6462932f6a3cb3ba369edbede3556eb6f8bdaf4e94e740ab8e5283c2c3fbf5282c0a3634a01cdbc54a34fc2c3b7f91e8e7317002dc8a6c13d42f659622fff9a181a53d3ef658b9b3c12f36c127eb2915438af834f993a6d5ffa722e0fa9760e43c1f7174f9578c3b4eac1caf798dac61a747e1c8100b51f0d6bdf0ad682e35367bd20e6d2e5a0ffaba92b1ec8caceca98f64e8bd5c0e0a2257ddd639a1bb8890e0318bcb786a1299f0ca222914d2b2439ac0a3459959992aabddcec3a51d91e9ecb9761cae87f9307c21cd75a9f12a1c22d464f6787859b077b1f5ed41705bfdbbd6d7b86179a92b4f052e42dcfa2364efec65c8cd30621d4b5381e9e4ee91c60d35083be29a8aa285c0b84b5df9584e7fbbf213e2d4eb00412a3f7902d1e6bc4eee65b156091720d962f7829e3414a3db5923ed1ed55843b4617a5bc3d3103f38af2ba4fc08a456e317e6321983782ea25958dd5536eb982ec79e076c049c39f8944526c629811761c0722ad069de5c5742196e8332a45838eeca797c8fc12defe7895cdb08e54b11f63589d3f086aa3dcc875c0400088b498a6e84b57d1ae06e00365fb71be4fdfd4fe52c3c5389deca11ddc2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he5547e769723a1f92b5fddae8d09a6d035997b3b9f16399b4c2ee305580cad7be633de9b5d1d62286b52032e937509b18ba1543b46c1242eef3125c64e9b037abc39c834b864ee33f7c1d339fab923243b5e44e7f0384180cb9c6a764640608155ef7fd3cc93d56953defe6a110a74dbbf6918e4083fe0109af906c00100d3f12e9d47b14ec343109d5e90712d24c4336bf1d39bef4740096593a945d0c58683d81aaa8934cbcbe46d8e4961f88548c6bad244234d2163d3b313c69d9b1b828f51c0462c87f15c2c72db746af9d564ff5cb307d95f20be9081e96feaf89c25e0313190c4aebd234c5756093a5691ae80523d25e6b354b994406a174511d3b31c6691ffb2471fe838f1fe93002fa85cff297fa1d094aa7263f95e0dd6f3a9de6001d46c9bb3a961237ae776d11a3089c186bbaf91594d66c1fd5c4f73b98f0d70eaee517f262c8ced634642ee47352e0f1d39fecc7502428b6694242cf872f585218cbe7d348918e6ea8e454c040b4522424bf49156fa2ca332a88aa8d3d931ee6af75b731e493006588ac90b3b80c9ed9c9de8cb28b84b0617bfb9f4f73d909a5eda348d2a4dc7ef22428629a2dde4e26d8730e1421917e02cd29d39208cd635795c9d273186a3b976ea8a0f2d9c17f145c0fdcaad3eb751803c66d294942434dc01cf801a96a9a415eb91f808618944645c22da4c0303c3c3a357ffb93b2520ac65a9089c0c1ba239587709daf6cbcba32e6e3e48d772b15dbfb2ab755757a51c15eba95e65a602fe68a248b9a7b5af7f35ca19a4e0ea72d630557189f716029af66e12058e79a23e0ff577e90a094d10d245aa8992e74718cdcb39228af3eeecab184049fac356a50f9445b75ecbf688660840d19144331679c15d623b279630ad00de4fd2eedc1330be1de7000c18de38252619cb54a874692f9a4846fc5122eb9628c9a64a881045af52c11e417abbb69ae448e3c6d95a6050f1c10241d1e53f101bbd8532dbe69a5479a6119e6aceab33d88509a026869655d347c7e212957c44c5cf74acc889a9e488aa3bc39db9779e7cfc65508c67eef37cd160884ba577d47265ebacbf6d3a6fcd4cbb1acc2bc017fece7962f2c63e918970d3141185bec44a7eafa0d8375c18ecb764f50b86e050b8a9f5fc543256ed8e57465f56c3cc94c8ec200fdd28ec3fdd01985c9830480cb5801e1b202659550c8ca5bb41042bd74f2af9bb099fe7e29d921b8de9b190ade1ac45ebd4bc808cb9d94eafdfac966d463ae5513b41fd4c5b9d46c51ed90501110f08eb69990bba96fc6bb3a39d505387c4776fc0db0804a36115a7bcefce6b71e8a4d0d66d18bcb6b666ad06e2d1e95dd549b33cbb23718f95d64680d4c38757eb1acfba20d8ef5ec58ebe8931e87fc67ae499baa121cee93dad2c58eed3cbdf10f28ed2567a9ca51c3f738f8920a790251d7675e2a0bf38721d64d71861fa8425847cd08766e5123bff69eb41934046a5e7ab4e7f501ec314ef7caa9e44ecaef0427e80a78b30ab73f9c504c5891423d4c91a750a284ad2096b61bdbd815a8084def6471408bf448aff282855a01e02af101aa0887e2855a1b39a4e3ce05e2c00e32f2e1f3b2fcab95ad2c3a9ab0095450f74208d836579be1dc04d638922a0ded0c4cd4e706fa557647f1344ec6250cbae32f1c2b650a90755380bc81c337d12b799733999923569bf0089e53213fc83b94c2dee63351a82840f3d1a3232ce24155ee4fe5009130f0492e3b5375c90e07565e3fd3a6f9540ecf6ca7a3442606232f96891f8eec1e2211eccb77109322e893beaa78ce7c28a64bf87f94a55dabf8963e45545c74a22938c1b5f236b398daefd265de3cf77f164380b55931f03fbaf7e4473d57cad25784ad79820ab18d0d943b2a241350fed2aad06141c74cf849cad4df80b7860ff758232ac7450080e3694d0f653a791404794113d5f529bccf035947d76ef09e817451d70d3a624db45081f763ca0db7bb51b5d43e1acafc7acc7b917e206e1e151e64587c87b4fd0c13e252dcbb697fd06633a4d1b9e47c693cbe54f961a73cdb3149c89f096b11836a232651279d899878402e4974ef06c0c2d137cfd0d7244870a1fe2ad7e2ea94610c1f6660890fb3d96341c1b99fab479ed4c68b4706521b4e076c085aa6c202421a3715c207926d4f23667d502ed12eed0330a44c8c9e220869a799273f9ec3bad5be3fb1410139bf102d046e634cccca5be7a0ac9a1a982e8b4ed9fe969dbb20c65db884637ca7f3960cc65cc90608cc4f2fd436df7337639822f5af71a28ac6223251631d60279e0ecc63135fb58f2e575ad8cee27646c29189046468c8599a793e45416352b13f4d887e4df382994d5af379b7dbebd721323b284df23928ec6e16bfdadd08a43a12f1e3059c51c09a100a313b5cce37ca0931a2a4b7b755837d2f6e2856d4b4cf739aea3a5b91cfeddb333df1d3218bbc4250e17b9d4e26844a4e4bb6665a67fb88d7a94f697396511eb9ef09c87c56d20c502b0e19f66c9d76ec1c5a42a9ab450cd19ff33d0b4b0ba12928af7cdf1f8ef371486dbf6d27c124095c709658e3ac18ef5ecaf61475cda38cb4efac864530896e82b80634f5a4484e73f749d76d060d968b2352c95d2e1bfe4ddc7786d2a562106bc89db6f378fd3336847c53f38145d1cc87421262ab4f363d95c016cfb450d2299e31863e008cc0e1d95b46150c248c3d82c342a3bd073;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hd4ddb96dbf627be9facc1ea33074ed20b1240c475b6781946bd802e112d2fb7e10648af1e6dbfa940c79402512c4348fd7956aeb27f884459c507e9a55f3acb5a7d42e982ea13257b8d47185dc4271bd795b2f861f1136b68e061efaa155210a93c659a8cc0d6aae3bd5ed3622c2939d1b4470e0163bf9dbb90addb7864862667032949389731861fcf465ce6dd43343209bd3c359809752a952331e85d8cbdd95f12ecbc217cef9d4c8b9d939df4f2a277694ccd8ce25f0432cb95d4ed26b5463510caeb8ffbbc733e746e11706efca9934a1c1c7b77ec5f16495b65e1200834151de78d9a361da4d49e97dae185c64d30544436d50c0b639c6dd88ea8631224903fc0f3b41dda851ffb3797c46859d7c70cc35466802d8cfbd1bd4cdcb504e64ee6bdf650307be34ff4bb463fada3b45e253b8522d8a9bf903afff75353d4ec03e3b39acc5d74ec163e0ab91a03a968abb585dfaac416dff45a5ca434368a7625ef0d01c9e412e538360da096680874bbc9e06f3974b7de30f722607a9c2cf9fc06e7cb06e4de5c989d6e302bdd78f8527ca9ef6de98ef42c770c0a6cc7806fe79e6de545e854d0fb2ff63f8a0243197440c786ca64d685ef92164447034baf8a0edda4f503fd5a5c18dec82f57b465856e725b5b72f0811ab8872d96daf81207256041e0f0c9db7943de414e7de03b93683d226538fd2fee9b2a8f11729d9afe6d57a1f77ba7a00ae1ac2f37599ba05b053a07338d1e28ac91fd2f0a4a08f534e7423fbf6aad3b6aa0fda1c9706d21b2c006e98b73f5dce62e73b74e550f97bdb908ba025201945f64f7997849f0858bf7162284bd547e0002f75ee019fd708b67170291db2e59d6f651f68a92133f341b82219bf9e3a21b83c549c1f2658be4e2e4f8ce27e54e5fc1287b06eef83f7cf379f6478a36ed37591a0bceec9900c3713da909aea515114d8e140d34685e63453bd2e2569d5fd4ed55694c62794fa1d6f41fd11e479b8dd2b81a4e2b34875945f6b0cf7eacb884756954ed3a1c430cfdfc000a67adfc8fe00cd85940e3ab3899575acd810055b145636b3a41ead330f60dd3710249c5648a04c81bdc1d8ff0d32e12821b18f6a636ee11e39110c92cf8da9f96ef87919ace0705a3bd713b3580ee1e8d4261187cfb7efc0622bce896db29611c53592a895f1a3247db4313cd91e103e377d014045ece4a06d7f7ca8ec704cdf398a64190ef2aa5069421419d1745a4b5fd23590d3475c0afe1498b4eebfd7b3f6a5b5c9a8f4d5b85b2d94c4475d8b483c561eba5aca8e1aba97eefbed46f1f5de58ac97f769f403dc8f28499c9a6125ae9e09db92e4cad3f76f82066af0653a70ceb7931383cc0e7665bb6671fabcf4bd89f92737705a3f5a589624f9b4ddef2dee461da886e70165027d9780001e918a9298a5af872169b9970a57cdbd78bf31b8a1e792d1c5dd8333e4be0ce89f775d50f327850b7e3fd9d7136b4f581aa5bf5047189ec5d4e9f492867b1f625c3d6c4009527d7a72f73ffc487dbbf432b2abc525482aed8bd2fd6aa4e60f84bdf2c99277319cfa0c2d8e86ae4e05761ce5731ebd5105d48fc05a978d879f7cebe5f47bed38ae2cfc34e92f3b1c73edf08c0dd686cb16e9387257a756013f0cba3b411771b1c7fa15a64015f6d034f9bd2eec73fb34b5a98000fcdfe0106141f3a99a1be63822371c410f3b538dced3ac9e67396ac4f898a8a4473802190a2a3197e9ae43cfcc3f75e5d2b4a7b43e7e85ca8a0c7777e712820f03672b6b949c9fac7e43409fc72844b744edc87e1613a520f1475b24b95ac230339a85757b580e6368955d00bfff53f8efd4effcbf857c2490a088029035bdc9a6720db64eeb73f541cfc114e11747f71a1e505ec12ddfdf8bee1c346c86643fbfa7a8d76c67073e9c96174a7cd71445d60dfb423e425a2529bef9477b65d31609b0a00466bafcbe45e27eda98cb34c0cde254bf7979a7e67499363fcdc13e5fe3129694eed75531feb104bb56cbd1a15007583b2eaf6031825a5927f2c1d2ae4d001d2aafe02ce48782343a3a52efd7d440ddce22bf9f5e9fd5712cd6a4907a1cedc85a44a25bdfa3df65c02b3048b0977ce5b5e793f16e7fa3f28c056d813f374c8baf936a50436433c98cdbc49c9152559f87cfc53f1f175d4a75e6c0085ec180a7300f88c6bdb74d997fa3c49ae1cedc3c1c0513945b6004919e6e9d8ca0d2719530b1779021db934cd34929ee451d30f80652362817ee4cd33bc406f60615b0b89393406fb4d38d7cd062afd3de170d609904f5c91befcad78a6571892c8d421c549f454293d7bc24538895c00badb09599a90fbd60758c1a3d33b7a2269d5e049303ce058c2c84e5859a558b75224eb99d8540b426b8b5b42e2d6cdc8ef7cfc8a6cc555f38ccd23900a73f94040dec7b045c7f37655d5324caa71c1f19c9f3111f7cc0b96b2cf7c813ddf89ba574fb20e8915c319c7e7ede7a57ad360c5f5d868a1298532351bbcae09abb59fc1dd532e452714f4bcc12dff64bfc01eaba424be947d139bb5f7be79ac3ac3743fe15dba2bc5604a3d70bf549282091da4e19afa5edd0506752a69bbadaac29c5e8eb483a315b6c38c09286702a0fa5b0583d21a2cf3491d62f240eb5e1f96eee4b41f10bb4551fb9595209b47988ba730e524fe96454a1f1fff47670cbe9d82f25d16207e36f739520a9f6c471913a8902fa624ade513fa6162cc8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h6b7d9e22acb1070924ca6d409c7f3bcededd0361e4a1644c2d55116600b29278bc4e363a0d1879cb484527a720e93ceba5f1951122240e4c55565a30d550ed4536ff1a69ea24aecbdf57cc696fe9d453fe99ed6151c0382d5c4b699b28c89f9e4ffe28a76c1808655d2e17da2de810cd2e7c66eff747ee3d7fd34c442de0601bb6ea35c15dd404e6dcaf03fcac620d47992e20ba209a4efd0cc6e06f576ab8b94fea9cb07617176dda1f5e0afd022ceb2d96e22130ee8c795823e9ef51c74439954cc4b993d69f2672b13f0723497e405f0f2538f7850b3c81dec8a5b106296fb59bf25fd1d342d414f98905e480f900925aab95191b5d5d6f9ea568e1339db232da8cd7d8eba53449abef36ba21231b4f22a654610edce17201b80339c4b1e8c5810a94ddeee8fbccb9186f8c570f5619117966ca79b5b9bdfe2e142372306f8f2fd45a40b97b69399f8c5c6fd381d3527c9cad63a031b8a31d6e281ef6c941bff36cd963e829a7875ee201527247f4b3347e420031ccc1ef2bc657736dc3e3981e644506abd6eef8066c6c0ebae8da5ccad4bcd59d13e8b70496ac45f3c767b02477e4f769f780a9d3ea55d5ab519c0d0ea9c89b1f9116e3b74a669bf8f9321172ff8cd2154a85a781c944db280309f9a677f155f703ef180af52767d5eb92fbde3c96f0f3c4faf4e35b65de0929a03a1fe3e05697e9e55ec672176439934f59c44d475221acad2207ae1b427a14082c63c5e3333d3ae55dbe65f520c93009de138e8ccfbe55b1196ccb946c9881c7e140934c21df95427d5697a9359aa7b89a56b6c19307d44a475ac0ae273d02e2529dc891ffcacdcb4e922190a670d6580a32e891370e26fa79d530fda8a7fefcad3d79cda700e4a614fc9850b3705bdb675ba9b268cd3aa523b41754337f67753c275df4b64886c58668c176cb512b0ffe78e247f376941e7a1c5f05f075dbac695256ecfec9c9da9fd181686a04f7dd0d69c374a4b9e0e2cab2291f716abc085251a97a461fdac39926194c978c43f50231efb41ef96d632e5bfa3f1d954bb3d9b377160a7b62b02ba6edea7847b8074e2688bc0b6270252c3c8fc23c462f3d76d95c1af771f93bac81638698db425276316e41f047b36f6b413af535a88f5cc3eefd0af1ebe7016eea571a4807ec19e1d50cfaa10d60a7c2f10698a04084d470349522c5a061f4ed796705710cb958e81ed688955de3b81d045c7619c619f2c23fdb483fbc0ffe2db4828450ad9254c725ae7f356f66f35696181d37ccd7e4b90764e98330b353c98254f3f3ac571ad251c8a8857707aa79a020002cd674462921072f2f7734995812dce643682987823d558fa27f38b2ab7b7d36b96db6f320c66cde005a1ad18f0545923d173462b9ff142bcb5c05720467709abf77c95ac4caaf3ce2b0acb74370e5ec5e7fd3bad4b6148c51e1478855c16860c24edfdc38634082a876b5c690e16b193e0438fd104ea2a0b3fe1661cb5074378d193a9d69563b9bc946e9d62054dbc3cbac3b4d8a0c09ef235ba1be656ee94b419fae03d7191f7035e02a3e085afe1e9146d88bad352c4b85ad8ba02aa2ab2f2f48b6e5b56e8cbfff2dbb457ad4872f736bad9c77ecc8a46ddc0a19108895dfc22903304572f9919532e1531216c44b3dc0aff165eb868da8b615c03d28d00d1207c239641230d3a7552016bfe44133ba34088fdd4f63a36ace4aba628fa9bbd4109f49bfa4630de44c5d58206909d5b4044633abc827d2c1824cfb937fb2e3d3c7f80c79b5a1c362f56d616e95a6b7553a119e52fb20cd7028f5d44c0dfd1d7a3c82ecc95ed117ab9e1c6413c783758d790213d37675b2d652d5828603a8e0434604ef180f5972604603cdf34b0915e43cb15eb11d95c9c631a297288cd8b87b0f30644159857fff9e61c04194ee4e8370fd7014293380e8198db1cf276bba6a5e9adf3b010bc24269886f2c2ff7bf07c09c760695f4608a76f26fb1857c1b7b748921e9c0d3a93bf2e2e29965a515f66fb2845232a726f6da6cce3a06c128b613a706c3b80cc3c43db6f4bb51fc8f100e7484fc28e75e2c63851a1a1afd1a43315c7116f4d9ccfb3b5334f87aad594311e30288b32ba53ef07181614decbaa17e289effcaad17dec6baedf89ff655d89e9a52358ae4d6ee17b500e063b56e7adebd6f317e00bba3ae0a9928ffa5ae90688bf804c3af44439f840dd5700e755dec836931b82deac0cb045606fa11686f69ffbe7251e94c70dc38592a903bd9de6ec7d89d6f993f0e3675dcf0c0ac596932507d4a91116e0c8b9cd75b28a72d9ea3096e7ffda0b827ca018c977385578f17ffc6ba721073abb53ca8389403bbcdc69778a9de85688156ca3f3932901a7bdb2aabe517ece7bab4f9c1c9be8ad122f5ab260a97a5cb310bfbe7425b2acba126a942552c31f76502ce55877a04af57dfcb6243e720be6832d9057490a7d53f07fdbf4952c78ff91f7a65830606338f4d5727e8486c3bd86d64bd86b9fc1d54a288d000f17d3744eeb5a977873d3e8ba522155a9c4571f105a2380d3c323b588fa38db62205c069c28dcd8f2510839ecd1a6616d4d0aa339af39b2b140dc925518755e8656268778087eb10cc6952bb554c392288f5da134d700ebf350a54b2aab365084ecc17dcd775298dd13dffd122ce3b8b5704b876eb87222298454ebd5955b16419bcfe614e8036fa783eb4a2e18dd64667011ad898582d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h72a809ff8a8b866bfb6dac4962e58853543b5c80f7f201af647c0ebb0bae1f09d5029e4a8f9b420b0f2ac22e5b8a2c7b41f4c92aabfec052fea773ce7527f4b700587f642e374fdde4d82ecf5647ef89c1632e4e6f7f53397fd9c35408cace3430c27dd9c3cb054d0cb641644295e4773698b928725aa52bf6c7e23434a84e513236e4dad7a6afefc84cf65ec67a0c031aaacde385071e0640f0eab7c2ddf60834426475a0fc31b28a815bea51a8d836ad6538bb9698c9feb1fdc3ee6478168ac57c4d28f3931445302766114e3d13835c7fa53e50ab5159057ae2cc4138e75afaca5432b3442fa4498825cde9af526f14270f6d81e4ebedcd297aaef3ff1caa64acc6041b349cabb35beace0dbbe81c32b38ec7c613db9242dbe25b95233c13ebfc2593a66b203c343846863616d7c6451b842457f3fe563649c915cb86a5d9b97c3e9a4713629605689a96129d9f318cd677f8eaf7bfef1e43c4092859a022ef26878a7e120045e9e1aa36ea3860977043445e69dc90ef89ab014e6b122a4c3b143c203d8eba2bf9be0bfb5aae0413866a8b292676ed4197357ca75f1c3793ed41145c7b9b110a96ffadd35ba4406a1c6ff7b12506b355cfbf83308afa2ef4366a46ed9ccb7ee2a18a11361d0897efaf8ae9c529e520a832936d96aea3535df859114066d57d609eb2ac24630e4a23cd12e08b5e59ab016fbedaf238869299b03a9923687ad5ab762b4984bc11d0b9c9687429bdc9aacbe09bf65a38e5ff4a94103d8f0b08e5dd037c81d1ed6e06f972f47031a1b6a5e860896e4743ef431b1dbba601b586561d5745dac381b2270dac3a6208aa15a10c05792365876b4557b701c7648fc75f388a9e849dc8d95f04dfb7d08395f255de701822338d62d4fc4bb735ea1ee1ee624cd12c5948466e712a19f2aca90c97b1aaa9fc273f87cdb6c188a1db2fbd0ba854ff3ba3a2dc28b94f6a50b0cab22a10945550f8429f0b69d11084e3f52fff1b7fdcf5edf00667c7757ff3ff3a47edf49a33cabb8a81af4707c03f9f64783a963fa0c2e4efeedec490ad986b12296e69088ad01ea5f1b998277a0ee59972ce89f1936a0dd7e9eeab4d240afed84308e98ba2a15c3e22a362c6ebc5636f29169f1e4b42af578dfe17fbc90c2bd2a99e8a513f30ce17e53687d424d64107e001d87ff2bd30ff32252055b912638e977398100a140418a1ba8fc6cde46344a00c7a028b892fb35eca5f6b3ce2152c909eb903855a1c0464cbf5f47746867a3d215da187bfd2fd94e61ee9921fe287bac56cb1234742ab953ac51dccc742c2d1418135f6cd62e536fbfd916c8139202b020d705041713578e324d2439825cf4b3a01804655ce4e40245e48fb4c2c37e5ac51dbed957968557f4404ad32dfca35881b4d28f99954c5110e4e7bc5d205dbb5674128c0ba7f8663a3340d362318efde747d733ec24ff04179c9610bec02f3d0f84b9a102e2b349c18160af2d503329ad97471e9679f07e237eb55edade0782e10cea191a4178f43c70f0b95a3e77ab7af9235126d366d548778fbc1020a909302c6f6a8c033746b0d2c85f7937d7022e8cc55589b25e886cedfe5a4d559af1733f1956f1e62e231ba9bb0bf12dc3d022a1cd14d7d664a1b97f82bf292c8d4a8d6ef95c0ee624198e918f3368b289fb1c468db62be3bb4793a0be8f2349aa46113256d479733ab39c74d181eff56404af08b0da2991fd1143f6d4b63d1fdeb4eb159bbe658d09fc2fbf4efc2677ecb1b351f72ec8928ebfb3ea4de70ed94d4508df9648a3da61e51b67a4f24cfeb6c20f2888b1a3a1522fa1798ca6f2ad5f0faa43b5416ebf408da876425cbc767110765d06bb1943150664a689c1b8099d5a2696050ea5b06808019fb8e8586554b8a9bc9dda76dd7823f9ac211dc952174a2782c0eb9996f275f2fbe864da4ddb56679c4437a54cb75a1bb6e64eb4e681ce71b255bf01b11585a220aeb9682eda592f81a4423fc432074785eb1a81d5a77b6d1fb3821692530913bcccf1a95a5eee02f53b0bb1b319abdc4867afed3a37dce33c7e6daeb38be3c941121473ab8f86e2af5a7363d78319c12521d13c0da9a539eb7ec7427ac7d99b6f249e8b95c7b5b15f5ab17cbea40004914a95dce3a260044d93d7267b2a146a97e225fea977f43123b5e315325f561894440b72f6c6e5e6c5a54e448414e262494bf4eafe15e78edf0171591c9297faaee9c6f00754fc4a47c91ed7a43130f712f671baccd33701c2589291bdfbd133a8aa9c5f0d13c40e2aa2cf6c8b9b79a4903e154739618ed31e1ac6b1375b015b42e80880762e686e0084cc506ab20189f8e6228cae2ccc1e29915cdec4fa3e5c51157c1f3fd243a3d74b0d103daabbc14dc6cd7988425d8525d2ca177b3bcc9ef971d4ba2d73ddb4c924ef60b612f08e8668c9deb6d18c060fcd83602429f9ea55083a8752d685d8638527c39625e5ce5e8d45d44f81f048c9850a129e6a670d57efbff954fb48b1031c1e2905737841c3cd00c675a4782be419110c81d82c700eace52dd94919bf23bbddfcc289345b71a9db0d5b54048c7ca84b382d70d1aa522337463c55fdf2ee80350cbbd302a9e83295c26024f98ca2c95ba0b692fca2108de249ba418764da04aa117be42347ffd05cfe7442aab51a2a74dacdc5b9733e4220e7d624d6671a234e9f0d82642c0590036b11a0eda1b8fdb90802d96f08872dad62c62b6c71f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h196c3099b54cd31720a919e0993a0d7fa3df03b37de3599a3ecf9366e8a133f410a27bd909e6a80af22265966fe0b58a06c8c6dec7cba51494e3f90492a3d6277cd7f136aa9eb68da8fd5046c4b99aefe8fa57228b8aa8913ecaed15b0167562df2627e03d564a865de590a75e6d01c143331317c402fc087c264c41874bc535f39c1f11a23311673cb120b5aa79f14c0a06efa09b1eb2769f2242f42f7f7e2cfea1ad10f4416b67e1039681a8b55693c90f086a4a6c80a18641ebc2f91d7efafc499027d2ec5b7ee406afd03cc328f2325e22a0bb9e611eba099bdb88b773737c1675654d17e332d38175b981a406f1c02a72728b9456bc0f87003485fb124a4dfbc63da7ff29fe36097605b0630597ae47f846a957315da651543543f8b16e89c132c34f2a9b9d358f73f4fc49b710e50f4b9d10c9544a0fc95d4582d9388f3843015b41e71dbca22fe6553126953b0b066eccbcbe514230aaf38953c4d4dc146305d1fc18eb17606b65fa58770ca94a842ac017caa05f45e7ae8e9b05210c36682d616caf195454228fbf172544178791ae432a8ea0cd74cdc394ab8614db9013270099d49b600cba995dd696caffbbc730ebbbfb73e3f925b707073c63317cae4ca610572ea045f87af099f40df44aa49b6332525ee91ba5eb5c3add179080c4ac630d02e64718977757a10515bef9f699beee60f78b4dd173ffab46bc6243bd223eb1f21c96830b5c5a8eb6bc6d3905cf3bce1778a4584a80fcbf779215d592f3c5ba49a3c6f4a59fe4fa01065a3abe7f02287a84f84c435c90a542db4ea9d1ee44b49fd46e7d8d30b9f13b4f0b7027048d62004500cd56b28a93f0de3502b2cb4bd113c769c59dbf81c20ce014ec51bf940c5f926b7cf8731cf6ae00c8549e580342867671f7c4d520850ab9511ad087dcb23be94a7749c530b925dd8a0dc4fa9cc0fca907229f448029f26d9d7aa9af07144c139e8212e8dc8a660b5906457918db77db71813d2b9d7ed13e2c1a8795ed2106b44c3d35fbae9a2044fa6b69315dd6248cc5569328c4fd20f2fd55acdcd52ab627a01a7c7375768607c829f6b5caa2b838092abde01bc64cd8922cf4af420a7329c124b340b9dcd5044faf18d230f473015e96105d6f2a59f3f7640efd1fad848ecd97eb9a212de49365f578280d980235cb91745216d15ff5c15e09511b118201992fc1314d8153549748a138e07512df62a99b55a7d63458c312cf59984dd37c4fbd47035edcdcb8185547b6897a71ad777d2dc0ecc60a1b429fe24b91365c8bb993c365ef8ad3b5823042a5941ba2cdbefafc0df904a0947724ab41ba5c4be6cc552aa57e4ebf5fb219802671d4725c40c28fe4e154445189058c68120e5542e1ea9192cc9e4dedad329e199a6fb72b5b08cd2a92653d439c2d662a51caa1055ffecf9fcaec598077a18aacab8f6537c80bdf3004cc5c5052131b56b720d805efb11f2e575354558c8e7d56eacd001a569f4c63ea9ae5a453c40f6f849f68a9eb2cf7af4ac57a1990d28a1832b569d3a0174fefb0c1bdb00585b4c8908aae0d5a680011493f7fa09391b12b8c62d7a6e2b32d79d9c40108f6d23103e069973fcba09e16bbc6994d0a755288ad1e2c6b92342ee6e25064d8b13fea4e556f08f67991e085936ca7e18fd81a188b80471bf76264d49c862958be797e2e4e966e4ae660538099e0128e356835f16e3ad01c42c62d72d4695127f8b5a8faa4b94a2c26006b5b99581bb42e8e284ce3ffe6aea8cf43f8a4776817128af2f24fe645fc0e78e41856ae320e8d23a7d775dc216ca3fd363fa9336c945d09f6fd6b35110251399c648b2c9b649b949a220881a73c62400b60fe591aa197ffd16347a2a4f308b7b93e3575d8cbc325fac4d3af6dd82125b9d6d378a8b38956d10c8e2432ff9d864444fdd43223493742ab194a7a8d6b2a15a9d8f775da408d8dbcbec3fcedc8fbbe36be35d3d51d80e51a53956582c5fc50867b69b8ebc59bdfae2095b33fb52399bf0bc84bdcbbb6fd5323f74150b5405599d85230d0e9d7867b030cf969de193863948c1a915b2af8996b987a8dc7132bcec0c654bffaa12d3f28381b4623c40bc38bbbb967b71aba9a25c86f508b68e04fb738d0c9b9faa774258ee1ad53274c6830fa92f53f35eda4a9bd2232e375986acae0d095af808551f6a726a999c1147fad68e82edc977aee629a59dab39bf2afe9bd84a9486e90f5d6eb8667a1798c05ba6d05503d956405762c37d30575ec53e9894b3c36a3d23f0a0eafd3b64352bfde1e75da8a9177dc56ff9c779f8e632a81b4e76059391cf66080d7af62d5210caa374646c7de80b90d6be55c2096300f4cc9fa3f4e18414ca721a9afa310323533b2a9d6c8e715a9397951ea80c21859c665af54617f11862c122b1c67de9d343a02cfbddd2390c53d57c7ff5712b07da092f200d50dc232b4ea49c825b4f544c7af78bdad76f3b209d1068ce8f78d96ecc77103c7719a4ececef5df5f5d9fa8ab8b9770c1ccf2c0efca37813cbb9ec26fdd284d586335099c55c021bb31b6d0baf238b992956476864d61ad2ee26b6711a0d81059aba49cee8dd9a41772bc1e726422e4f24c9bde76120491faf68050aa746f4aab6ae64b9f18e9abbc1b52d8e1ee3eb028548ee60cf52b962a8f06befb3baae20113add9ae0bbcedff955474dceccf4adcae553cc41ff08e731f812c411062d4536ef1d5ead4589237;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h368037dc2a2e4babb7b68fc4294765d76c6c7ec4d74b7e06e3fddaf3e75ec49c052a0775e32810dbad0914b69130ef4a6afedad1af4869a5178a9b81d99aad5967f7f00bdb570ada13a11e0a202e7c2abce05ab9554b9d033151e83eceb1dbbcbf9a190ee1991db1730a8b0a3e016019ffdfcbd18185fbef126cb604b1f05c45f59dc38ed095bc8bc50eeb3d01002396aa6dbdcbc7acfc37a3f5f237f5dec68bef97180fc61172955e635485bf35951addc05fa6a43e98a9064e9ab1c69ff5a7bc95f7194c94701a9ac9ce431207645ab454ef80d3eeb57e2585a302d631c73f595917b20544b870c1d32e59f725db886cd35269d90a200927de3f56b616df504e12c5545dfd0edcbeffa7d72f4bb17c7247377a1903e21b3d921962d12bb0b731762db32910a83ba95d561769ea2cc4c9459e1aee94c5aa183d85767e321e71339b54f2d1cb27c996ab6b3e5b8c9cbab8a3bae4aedcf3f4dcee8fd48dce3b708fdd3b8538e01985b85272d5c9adf8b06a79e0b5b9aa5aaa506f67b64753ae5632762f9c217e97f4ef831d7b82c0a53f374fa66912c33de95286b9872d0456e2b028ab43af52ee932a2d1a773d18e08ef5ca24d2db9ea9d47c940ed91d626624620409d39f07d7fa8adc55a3e65526669b8b0e23f605685ffed6a8a38156a796db50fc38beca7398d4988a174ece3dfb07900f156e2d996c0beaf6808bd9ed74b083abf9ad181b6e69f9ac69a2944abd2f6a7c2a1d3984900bcadbe31893b19d92a37bf088813a6360f45798140151ba21cbc8be2fb59dbbe21dbf09fa461281d3396c58708b120b87525b4ae8b2c5665b57620a7752c61d9a3a3b5f194d91e83c6e8a5de61de12a4ac28113d7e04eca82f4b3fc7461e5b9f6a808ff46f3ec5d7ab72fb3805270e3867a3dfd0b167b3c3039beeb9241e71ab426e7158dc62fbd88ea07ca63be9088c3eb46132f7eaf54d2765f7f259deee2db43f5ea9f852f43bf4d8a90d3d2d346960d689c6291c1dce9917ebad516764f73f7b4dfc4615a110dfe57de3fc374bf5f250977dec1abebe073d24f531b69abb6139a4f696a05920a2b7f0ae8245c72658df183d0feeefc86b5604705b18af6f430d7675b635e15b547049c0f9f8d7886c4fc15a52a5ff63a96775c3cf171b1e98ac85cec26f4887409f8cb8bbf1d3f968e0c81e1b3a2e9345aa5747a72cd24cb9a8800a11c81350ae45d90c4863c02ce28effcbd0501427e7ec5fa6050810adab7499174a8ccafe16cee20d976b63e32f69e315ed146d8ca25e0035ded7574c439f6659b8232a9f032dc620ae9f23f429544286b6127b648cdb6c666b9c53763bbce4304566c39bd6a23eda17b765b0278f68533e20c7434e874aa6934fe5c027d19350ed09475d55efdf18277fa66533c9aaedfd1bbc7bde1d88e9efed05fbb7a298eb300151b0c8e9e06081db120ce3aea96026cdbc485cda941c082658dd9deab58e8303cca333c1e5c46dd6e186ac850e7778f820d6ebe12216283aad46f6955c17e2aeffa3b0ec023dd8c4ef05fd3fe4de24a34adba3a955eee95c0adf31fa2cf39c5c5bbef2ecd881ed3efa2e0e0ffffe36d2b244671a92eda82f0d7c0be17e76adc3c15943306e0e8a7384b50a7f6883cd1d89f740e8a018f1a5a5227d2e2e39cf57bd88f4f2917d0a1a90356fed84cf59662e2def1cce663af6f4e3488bed7a775229adbf1964f41f2031bd2f44aa847f1ec8cb9bb55461943722d3f5a37e1a891adf45e64c1cea501f3216c4cf80e47e2ac661e0744405a083919b912c1ff199d27718c7ac800fa4b8870ce40df40fd5bfcdc2dc771b85d23acb9537a7b77a0b403df0f2bb7fc34bef5131bdcd81a08636450e7f49d14d692dff9c116d9c1c50a601a4f36a40d716114d955339cafa1498b97cdbea3c68290cba064226a1bcb279fc561308ba9d70d4ea97ed7e8cf9015bccdec64c97b2e04e440cfe15d52ac0e65c3926ff4d092e155ca4877897312b0448fda4882f82453b15f21b69380730910f8bb2c1304cc4405fbc642768722586586b8ec20cc9526725438bf82203899321d22db0011be0fdde9925a8e2024d3ae52ab801b6bad90bff339c51040974693b843f7e52a55c232eff0223ce5d7d47346f005f6e00bd869a8d24fd4bc96670a869724323c2787e1c83c6b2628768eeff25a1d774a89fcac178f827eca971aab6b04665d24868c26b949ecbca6ca9a9a2770a3a0b422277f468d72a5485b7cb213992a08bc6a84349a7a28cf3cc85bd8a1d19def3d5c1be2a32d80323548a3f706eefe0af351d486a0c17ffcdf3daad1058f3e68dc8098d2a339b32abd4c77c3456e8c84042bfeb1426f0f2bdca5a71efeef2df375beb2977b8efff6d4ea23d9fb4e6668da50802366cb0dc95d17210393ec6530fb0e98a9d59eab9a4ee3b0810826740818b2266048f6311d2650b76789c3051dab5f2e4f4e9e83dee2f70cda46417c15f5bed3a53ac9c09a3f1fdcdd6ba02193e5fee413f1e68127b6fb56351b48b0c7573c72f2960c172d94dfaaae96fb4aa40abfd728df1377db8a6f04d6bab424173f9356709a60a5b54775d434f8a252d9bda36d4c9a2da79db90d9481a82b3f5b04cc2e1ca2a18c95a3da6aa1e118e8cd77ffe677aca404de428818dfd0600623a51a34a25febd059711569b8dc16934c03f84e37ed05f79f431cde1deac6c9927a74d24590c10d2a6b0f23437a3085bd1dcaeb1f21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf6f5924c8860e38549d330d545e71f3b1e79dda607393b12c9f3a26baca96eebaf7673d19b3508a065c5a7dde1f5916ed6c95f603b9f94be5636971221d653aa21e62cc13e9f154f4a77952ab886f60900359e67d1d9317ebdf715f231f6bb7789a238522fb2fa669be8b5116d4225daa39e3de947c45d916fef46004c65529a639621a705ed70c02a72701942964159738addca431e8d72b0ef6559e4fbe57bedbda8e794f20534f78e6e342cd925181d7e123562c7ff9c473fe2fd3f4fe4bac966de5433cb369429eb23e7bf0ee78ef8802a28601e461cbe9f91fd57ee563e8f2d56763e6a3325c154d187980e6cb1a34b16e8020be16bc2e3ab2a660c1f3581bfc23f0bcfe426da1a1ec35289b725ae2855b937a9a79a8692aa0db8091b47e05b7659da492bbe768e1b7091e3b1f92935fd5bfde2fa73ef946d1e22c5b713af18adf803576141d86071323ee6ad06d833fe60b2ea682eed3008ffaf9576091b04ab0c70c408b0973ea662c6bd9038756b08b3a5c49b6fd1556f6dfa358afb3cc1d0188b2c20c2cfb03050b696e0c9a27e137788ad6972aca08d88cbbdea165e7c0dad1a67c643185e04ada721b7af4bc66ccac6806c540e0a7efeedddfa87ee2dac34b229efb382787c0c395d74ad4bb24ea2088843161d16d5a34bfe9b4e5b9cbc6114ba04dc29d867402d443caca8783b51f350a4cbb144bbad43d9f07cdacf5b173af6adb0643fabb5c188e9385c8abf2245b2317b13267c7cc7ea1f6e376aacdcc0ddbd66577eeb67a645c43c5185adfa88093085e14396b6b967bf107263e90d9f3b23b5b93e3e0f3f25851772a50736449cf47693e9174010ab9e49bd01c41f727bbde75e1b613709817ed495bf4bb12c464e30034f25abf7d26c1dbda6b13e8049a9aa9ece742270558863d6160dc47006837ee7d07474d1a9e4f80f5c193f0ecfd0316f413032208d1f1ab2095cd3efb0547b54923313367ecd582c507521bd3f8336c7de196a8b55b5c1039c75c07ed3e6de642e289fd27c7f20d312ae7b86cb3b816d65fb477588b70e970849371d28dd0cb4bdba7d18dc9a5fb76005426b3792777e138a37599cb5b7784fe7f1ac6dcec78cad265d11911a0fd42edf2f0242c0306efb695c1f8b69ed87e6acd85c86750c6c2709b75b0302fa6e9da0f2f7e45d23aa2fd16052309c464e9a515cae7306d7c43144d0bcc2d74900c92051b4de7b7a53723bf26ee4cb25e72de40727c3f523d328d517d60cd6df98b71bf32b4f1d14ae2be3f81fb671bfd75634197383392b2303c997fc31bc511c03fbbf83ff9603a3e240906c5bf4216c9aa7d387c50ba108792091cfad202a81db56118625a56a3c4ddc9595493cc2c3543bf559b930bc189c27dcb069331d77c812183169e3261585506ec1022d479e2d060bf975c4cf279712d57caf3ffb1cccb33d980d5bde1ae1293b11d477f55848cfb8289c9710873553969c112345b576b498b0e9cfb0ea34184b3fef572bd4c6211e4add8ea47f2790d266e292336decd81a696e5e6801b44e989a5aa23e1b2c799c449596c2b1a23a8b350e3b914c0d5f7db73c847361ad3dd33e0e540eb6859b581569631ef9d0413e9baa9060969c55bf9820469c45b025023c83a452d4ae17c84924dfcc2c76ad65e7ec10fb0cdba5f8f2c4855e34f8c5cf7545fc89002d89bc90ec5a727bc465d145efec58a68c292f801902489425c66fe4fa3ec3954db92c68546f490baf956f4c70019203b0fd00b38c389ab3973bc73d2423fd03870bb49bc553500dd2931d302379de2b39c210c2b996c3a5a5fa1c6c3c39254fee83fee7c414b16142181d300dabd3675880295eb41d3df22ad38c2271c390a3c54c5fc47d975544ecb0311a6b456db73963652174b860efd73d335be7d8dca0ea9eb8bd4be186bf5f96f8027af3dfa76cfca8b4da93c50b3794b0ae6e653b85b2adbe7039b5eaaff28d8c354039747e921ce8f94d38fbed847f1944e5d7950339490d821013d4c56d8270fa7e9fff380f31af2140c1ba4332a32f0647355cd6a28317ef2f18ea35237f148ef4aa960d76e09a7095dc9004be813c0ff0f19fac810d901eb0a0fa7b457ee581a4375ddb67438768594b051a8209d49cb9b38712e17f6fade5f1ff1aeb825e9d5e7fc061590fa145679f07f5bfbfdc4a5d1211d95dfe02d854d4783170543d67319b55368368a4e4bf69fb371c394533faacbef44f075f695881f74e535e29505502378b45ed931d23cc747f8d0f58610e81b99e8aab0233f5a32acbc415a1250c339f31a05cdd2704a0def655c639dfc4855a7c60b8bb9cdfb68b67d26bd74ae9e089d8ae58bac5464de1eb5639be59dbde552cd572889ff57d352cce245c6c95e22bed753ede8233a3d18fa21d3a8aec46da3b517a76a3610f573c77614e917941dc976c8409183b2449e49aed46e7da350496a1a5dc87da6a0587de742ece95df40e1d642ae2f150081c79c981d7bbd27d5a4c6121675bc368ca760848e6997d3ca44769f0707c3cd99b417392dd98fb26d3ee5f64f2ac908ad431d279b53e2ff44ae5ab1898f301ffc932f0d18f8041b5358f93affe9fb6743ed92131a85bd67bc47b84d79b8989377e66a6108f89a481200dbd5aff0b271dd695eeb41d58fcac08efa79f476d7821ad05cc70df41f989ee29846ae63d8a1d81560864025f5bed7ee1f52f00dc74242d6d2767bfcb0d137cba96c01a919deb9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf93e497d222c7e5584dbeb4212a71aadc16702e8fa2b3dfa6c124fa23340b641e714f10db3ba2ff967a86f1a33dd677ea5b2f43903394dbc7d15fd5bc2cf5cb2f3bca65e784e0d1f6e36b6b95cf75397b19eb5bee2e9718db326dec5d2698cf7dd81eeb7bd6caffa93909ceae355775064c30d53c5729c64ca163907246260632a8fe9b1345cbda8e11bec21ed2cd26360427069bedd66e9888552ff53f02a0daa2dc0095262eed715c086680d68234b0b3a09409fd4f47d4011c2d79940a845b2d36bc7b7857d5c45bb81176983e3138f38f7982357a08e2cc12e3a30fb30d59c4bd91f0f9a95de4ce36a53b3842e283779636a3e5c3f1892a614a95bb234657ab4a9c61206671dea396ec9bc89d87bd1cffa8840e14cecfba162987dd1c67371360e68624feb436b397f02ae416bc2d50ca4974e75839d92f0929d5430c88d1b4973b83db42ccfc4b61ec06ef3a0311951190e674e159bf8c24b6936789e46ebd5fbc1ce2fb5457fb1c3416aad2e1e2c6c0f59add8f20c2c0566df6269b54658bdb876913e1b3e99819bdb6c027c9062fd95ad33ef101b202f0b678b4a2c6e830fd8da09e1393a369ff128add932c69189ea594df8e8b064a24c93425bfaa9483a822a5ae146219245d30348e98cb056138c32b44550e4440fdc4d7a0f2cd47402c4d84ad3d464cbb71291f45867de1b5a5a0f1b52065434b757c1c513ef758be540f55b266c56f27552ebbd870b54e31ad04b1844c046bb641c34a98ae4f252398352f59f46c54542f774bbd85635d0852fb2dea8f7a3f351748052ec00a02ddb4980bce1535fb358d723bbdd6d2590628a6e8634a6fb5cdbc7ac86e5ae57ef6530bcdcb2b03b04583a397c7d97ede10e808118cf706f8899f7bc9f75a6b62194a1f0d178ba9b8f41a9a6dda3b212aabd38409a5c2556cff2cbc68c3f4b08ad9d36632cfaafb90b5d6e82a4a3d87695093f973db935f8dce4c52f30541e4bff955a3e64691da57e0f6de31cdf680f1e62aa90e2a073ce51921e43d62cd33fdf0df15e225606fd25e4da8f0caa660b50cbc4a7fe66079fa7b395865f5f20084b025d27e6b3132471c92872b3326ac72d0935a8196c41348a38ee6e2b2e8a290d94193890a449867577153343a86b3b727e82d31cb3fbaf71a5454a98c7c8419c1688e828c78d62ecd01ac16bca3d177146c7267687f26ce72facd0dffb845ef69ef6b01b463eefc9241f1a628983bdfaa2d680102abd1d5bfa3e4d08b246e49c5ff64968c4d361c068f8bb99260eb8aa83e9b55dc8b4baa0632bcce6960837f7dac0f0c3af6f1b5422caf42498678d59bb33449784e9a6994720e7bd836e625d79506a9eac86da7de520c965044e6f0ee62915faf744e48ffca5d184d0c9c6084f67b512b7343bcfc0b1c83baf26137f3072a15b27a3d1ec04d22c4d130ca713203806a938bb6eb5c5670b0436e0f6a3c7840a46b89e6cb90e3019b56b763e4298c0165faabf74b8d771ebd39af34f397c64702a31143bc624ce76aac9e06ccd5b61d47f40b27bd875d4b894274a2c669c648f85fb146f2db0fc6615039e34cc764234cf94196db116c0543d7173bd0a83140335fffb1548ae1816f77b2bbd8b23b1be5fe46b91e67ef8a41ff95bb85d8c56021674ebfed4fa8ec8893a97bd16b072d13d2c0d0ec6f226a82b9c7d11573337343c494b100212d496fe73f3d03bdd58fcb30b63b9240dc59352104d3fb8240f0a7b92afc46790a455fcc4c9056e0c5b6714159346657ee1bbe482d0e108c1cde36caf03c40a1f9f5ddc0f034bf8d00e0a70ad95113c8500d53e9d873e8353f28e8d15c77332b60124107e6f85c2e2d3b437d7a017866472f9818dda5f1431c5fa0e0fec0aa2d9a5dc2acb49c6027ef51cefb30c010b75355bce532924c3b72311c4bb84f493da4f32ca2969f8f521cefe85dc04b440da10e549522cb3349b57fdc21266531f430e9dce5f61742120ae13ef928a5a5140fa70eaacd2a5b77e1c438212c7aeedd885a7473a02c1183da890cb7da2994f1a791dd511cfdec0825b2ce82306fe2aac9b15498ba259644de51c8e5dd0c53f258672c382197730ebdd2390dcaf031173dc701d7d99d88e335824b0cfb0abf4dbaad73ae843aef5c912e576e4b8e848b0a3c349a97ce91283640fc759cdc0ca9ec2852c3081855d7fd564c6bd525d1408adb3c80b1f9c123accf62c36b004534cb59aebb80cd1817b81eb8ae1159f8a000ec19d6584a0b833264f9bde91b5c85a17064225240c4a63474bbbe38d581c807899e4a4923ec813689c858dce072e8356b9815f77daec1b9c30818fb71cfeb604a60256c79226a898972d09d6ace337fd5badfdf8eb2d86228aff0b2435dae2d8b37410f85447827de30b320bb19cce65ff69379d4596941fe766513b80cfe40da5823c4df08dc46e1ef23da740372230b84af8e49035a93f14f5eb4727f970f8be7285a163a34ffe9a4ac8322d3029cfebdb9387a43a74ad2126f1901b8251ef5a5465cdf7eda8173e778367fbe6b54b5536c75b87f2909017db156febb64afd2a408c8c750d507356bb5330ac99f491e24541767a735a21f97578cd0ddf2f9b0d4a18f3c328282b7e6b179d7909da1e4d9c5303471aba37cafde359ded46825e275814312a4422ddf833ef11e34b3fad004605e88df9fb9589ba9e5f82248e06232dfb2230e51253078a3d371035e379ae284a025a21ed5bd4b7145df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf78b35de313da570f333692249d027bd4183222ff1cfca071b35f0f4318fbf449719a9753b057fcfcaf85dc222c71175c622623dcc276c587730a5cb4c77b0c21888233305ec9917ecc61f49927ce2e7434a02b30e13ecb6ce3d7443a2c156651ec1fffeab1b2a09acf5331a051407106934e29091770d43eccc662d0b2d0a9402c3b48e6c524af678eab64715f54dfd70acc827a7e17e0823c76a85c640a5d3df2bb12b02c18d99d5c16f0c1295df565673b691d3bb3baf3e5d82277a324392644d56e450287509f2572e3f633b8232af89c6301e6b0c4e7d9bbf6d2c33ff52cdea40a4ed09bda962f276c62a89ca7cd7bbc2ff594f62aeffb5f93c3bf2e27df3c8d7bded494e5a85ae80e80bac1b44c36f79b2dc3d9d4648b079eb3dda20dd3fb6a02cb2697890b39458222692c883cf81172b87ff7b2c6b327e38b0413836b87a7d8d866161d3f7398891024fd07c249319ab40aa430360f70164110056fb9424ec0254ba614fd42b83971512f27855a2ad08663f0f23ac800e7e689b3013f2857b7372f06a1d631872c83eaab14044fb51b91a208f7d9690db2039ab2d8a451757f112c6edea4e3920af3b8ce03d9e557c0bce3853b840308b1bb395108297f8330fd7328e37257bdf640d96988dbdcae7c49cd622f43866878f09d3231cc2e3a9500170c8e13a63b3d6caa739dd18de83918a22e7808e638a309a4f15b92e584ea9fd2eaee042b7c780402865c9f5fb29b6541b91408199e7a780ebd40e7c7b141463dd3df79ce08c3185b075904c779e3ed71406632b72ce21a7cb2b659b33f62803e92ed27f4c61250ef33eeece85edf637aadde2d073ba97cc255e6689a9a48dbfaebfe92632eb8638788fa753d635017bfc7da6423578d5d442d1bd224d00cff2bca6b9a650ca0bfb95672d4ee6800d214343e79c944f121b63ccfc45c576556b3b3273d5b5001e731654b46799c8da9a10388fba165a9911ea49e8cc181b01435a0fae5b922e950ca65466f805749dbb2fb14905ea66fc7fd949a695c0d764b3378757211c8dba2f3cc11198bd9d8c92eeb21db602160e3cdb50095db70c7a5cafd7ccc165224c4a1c3d967bccbb5d78ceffb6b237f049b24609ad528364af64971d951375090b9bfc9d5d80ecc2e8e476e8f71dedbd1376987dc07ae7f3c651a4642421936c2d0537670264cd307e610a936635fffef5b35e69e0381a7ec3193774fd2fdb8349c046bd774b4064c36b35fc63fe9aed3c9435a34d9ea0c52f7c502cefd2deeac4a6e3524fac894808703aa954ced4afd52f65ba9a243d1e13a0c8df6d491e34521019b3f795593744e9885e20f157842bb409d14cade961368db2c7fbdd9f5d6d541033de37f07752676a25dac618138cf9d18d95656f69124eb5f77d914437e8858eb3f6c88ebba78a152e5dd96219369d3c10609ee81fd90de655e838dc3a5ddcdf36324ab07c0c24f4297594f298a9aee2880ef71dca6f71b493e7df549e9992f0ce80ff49ff6fafd17d76202d4266fd6178d3c5cfab9ea82ff73ab7bcb861a0c49876f90ec0afc94a883033449bcc2570d47a575f6ee28b41b97a4a9232c370e2e38f81d47742749b025935d51693bc790dde6b4cf5d9a37cbc1ba827b44ac48b738e265209dd0453d0dd5848c50647ceea5480cea3f0d60fa45cda4ef2e66cb6482c3e5bc33ce74b1ceb6233fdcb96952635c737ff5826a8f136365e09f4651fb217b31c93b3ed6e6a268b568274e8987b80b5f32227766e7541dda6c9c8cd8f38508f58cceea9bcd7b59a4dc79f295d3433bf1efebe909586cb29fa2fb720c53466bc540cfd0a918592048506a5e51cb1e9ac94088abeabd15bf4fe9c309f751d330a315adada776f49d3265dfa58abf23aeb16baf3863f12f4dbb73ddf53e65cc086bc629cf2d6652d5549608464f833ba500eba8c5aa32d29b21da390c92da312e2b4260b646f1588e083b39121a39f3713ad02e585387bec76b811bced2e295c2d52e53a025b108136e6793a09540f4957b95d0b391808d5d4ea4926146a551557477e9c6ce04591fd7e33c459a5b19f712e4e39971ae00a75e5a4da61d4adb64cd3977530cd760b49d73cb4cb6a4418eb2e7ceaa84b99586d017eb046b1be9ad0d5ffd49afe650ed2035d8669205ac19a8a400518fbe44b88852267389a469937331bc2c5a09de9f24095466d3b92a44fa8d3e99385edab017591417c0c7d9b8acc8760b9f5d67f8c23e5635b58b37ce299f0b372d0f4c3f2c7dc85be3b2bd3ed0759724dd4a91279d6d7af9646d7ea463b11f6c587f0f5aeba132bf9ead0d0dfd1d43eed3f47d873754529020a4cdb29892b77f4a9b6767a25798635ec278c554fb6d55bf4a81a7be9779c5cd70bd98fbcc3626e98d6f302961e48b5e56f22e5a196c56ff25428a73073ee6937358916349ff2eee2b8f75b90c80c11742eef166b938566063fd785ed9cf95e98b5dbf41251277142ce445e5f208fa84b8fc9445a0dd9b40dd92038abe11dce4aaa3ca47cb81c8c7e879af7918a343734fd249b03b4aa1629a60506af9d3710c4520d72bb2b2dbcd6411561f07bd4e162d401c2f2ba47542f58158476e58d48e3fddd11fed227abae6c37d8fae00390c98854549fac8fe55eca791b42451c70064f3ee02f7a54d57eb17ff1e4a484cef5e89a2dd7faa02bf1db7507f628e11f68c809138681e7c56e321716e6ec3e57a6f7133f0ce5d92e1531c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h88e80839d2cc2b265e21c920a2afc6bebd049bf6cc1db9afa36414727d43a7809601817b2ec228793038b1702684739893e75da32fecea44cd197fef40b2592650c7ee3353919c357b4392c45ebac62997e312d119ca2f94b55871f0f7b23d78a411f4da79afe7f6bda9c1093f87621417c4fd3c6601613697e847bb07bb21489511e21acd3eb9440f9861bedecb6e6fccd6667a361dd605b28ad40608c0616c110c4e404324254452568a8fa14d75140db180f7a6528e99cdeea252d5efa5ff9d25b361976b2d47d64374ef76679060cc142b94ed33297cc38ecb9fb8956773935b051534ff300c2207e011a753ee0dba3057aba8a1685939365d2d66d5e0cfd1cb83b254fc2727124b5cf8e2ed80b628af54407577b8dd502782f5dc4d729efb84c7ec2fdffb10502a627031eac46d73bbbe31d2dafc8c63644239c97b46955830cca23b5d0d36b1b877fe08a3a230fec7750eaccab95b53a2433d2429ca96052d8b2b0b930a0c1483e899ba9891b3f5f47ab63cdfd3c93b8c36bc3cc54ef7561402e6791025efda140974b6fabf201e4f8b575566c31c84a5cb7602397f9d127e5360dd2e2698be8f8f73f44047df71829d2b9bbd3cac87f4101621da36338f242727e0ea65df656e890baaa64e46244eda526920de87eb1c5712005b233e477c67d825320413fab8e45bafa2afbf64d2cd8b2fbc6a3ac160ed723c04efff55f54775f17bebadc39bf9db48c6ffe6ed4c8e211c7d09d63147e66e125586b3b9782f7eef3d1239a8a6471b2469b8ccdf850ddf24c9ca359d9252908b7b66e78eec87400860613a8e628c87ccbac3a98b40e2ea92d54d28603423b45813122abea288a6eef4f17f9e4d2c627e43f6d4a9b562b797ab2cb4b23740498e9ad480819f057d3929d2cdbd663c7ea95a9b0cc4487bf236666b6246a1e29e3fa83db563c18cd84430e1c910900bedc5cc10bf40ffcb4d8c0466dcf12e5d066e555ded5f00dd10a863ac25ef7ea7d08a2899d2ee0394e373df6151987e7952daa855e996fad0c1ade98d7b249eb58b7e8db4716b5eb0e41904ffdb02906f9e2d5b8c93906fccc658cb086ad14e4161e288d387ae48805c21f19a1aca00c85805e7db6c31dabeb0706013a06dbaff0d255be307f0e4b38909f4c434950089dc45efdc30f155d20769366755ed17ba2b1da6e19c0adba68683dde9e02a41f7816b5e3da15c3647a1d4a3818b649b702839b6131a4c084c2c0d8c318887e55066ba859212405e589bcbb55c48e2dab0787804b35057d145b046e020cbbe3ba2229c5ae6e948233cf08f888596922308ad3f05ff322e3e0c400f7d384976d2e455fc01e06163821c6a38c0684486d38c68acaffae40a2db39dd86df12280fd07ca6b2e3793f65affff76ad75aeb41229aab7439bcbf988b9956f31c255576826346450c490d6be4aa80994418640d71d50f8d1f640374315c8cc8ed21cae71d2c8058b191a65f9b19835537b36870c2e7b22e74d2419f8e809fbb8ffaabf3650ea013755e641c9375da4624d9906a1367a2e3d18b550903ba4ccf6923c78658e6a87eadfc0e7ea8e39ee1a916889fc2b601f9ae669bd0e57659697524811f0f934706870d5eb447c5a754d32827796da29480623eaf3831cd88c2d2ce87663e9e3ea233981beaae25ea6e36d88e9a00d6821e71ad367b05fd79daba7876024799446016bcb4de487d9681130590cf6bb53ccbcafedbaa53905368fea6837a53a9f2f6865e4a0a34cbfd82e0eabb4a492a203bb71d85fa441e6e25b04b4ec64a01127f63422420f51cdf3cde4cc4c79bfc73f9aaee534d351614284ae30447f03b3c9b3c150d56e4252638d624b8ed2cd26f4a12712302b75951eef0d49709dca109bed60f0bf295c563da3d75c5fe3c67e7821b788b0080f223af77d4f64f694696ab9241af53930615ee92cdbdcd8f667cbbf7f0eb138ff674f445542befea120d1610d00029c7364e7101dc74ba190d88d286980c0a4b6704457af9d563ad0d98a4c5d301dea11a05e44bc8215db850cd42c46e6e2a7b77f568404fca543a9ae1eb072a8f61af91f6f83bbf813a67a9345854122bf988ceec8f20dc28a5825ef131441b9ec156ca62a3bdbf4cf71480e021537a69545cfe914a2f9a982546b8829fb305ddadd31c02c40178f34163592852c1fa1ed7bc49bd160fdffcc32ffb66b62edaf79bbddd4e84a59d74930a071ea068547e6c092f40019b135222832fb7f2a7890180f211a97da9c836f0d8503b42094983a0d8bb147cb1d61be904649f7a1ae3751445b81e1ce68a480274f87cfec01c55a16197bf404fa262004224823b9472443d69948edc8f76dddc98e7952074cda63786bb12dd82cc8264dc3f3f47dab52eb8ca52f584103d14c0a4d4f1b31fffcc793bc19252d074d3bbede69bd38bc0f1a0cbf89592189b5226390f99aabf577c86940a8717a1f9dab8d88d1ee017897ad1b601f30a5f06398b230f1f0e0d27f76e91513d313a4d184cf23140508d1e421676b45ceea8900c91a0784ed05061916a862d2743d586767bc813e231f3777964d50f5184bd17f3fd385f8fc9d8e5e665083d8fa767104b93a4cbcd7fa7e70757972fdd11ca6faa66312662bd37afd43de0043499c53ddc6b4b16d578fad4a45253aed685bd59790ba92358171b345d55e9099e8ebd12e15b5a2873b2e0548a8a5623e4323333955d0503e661eab5fd21c201a72747172;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h714c373c61218fe257d1ff4b5a660deea86ad1dd22ca60b65aa5f36f28ac63b54e89a88d34866800df081563debd55f0ba8e51b1ed52d3cb4ad2b1b7bf891575dfd1c36e13de6bed790cb78c44f129f7a79a25b8ffbf8887cd40c20c3bbc409b347c461f36043dc00dcf293e79c0d0cf1357c9a25600ab498b7ede9e73f225c7d90f157a2aa24d2b0ed6ffdd4af48c8ba46711180f37e2513c59e5a20959abe8fec3eec069efdec710121fcaea79e3fab0e2655f4667ec78e54abba0056a0f9ceb0eb560ccf740006db13bf1a14b204bf0c2964236432b6a125f15a31fea75bbdedf4ee0c4073784ffda1b642ed2043592684227ed17f894ff9001d795ad444f13be297b565922aafbd6788c0085ead2700b57e75effd8d8ca82dd9bf71ca77654d4296e9ece57ac7784353303b22d557bc159e478ac185e1174d73de0ef2c4ec246e7a014eacf9736c11d6033f99629a6fd838218033ee3fd17a1a7d4f776b9589d909bba650bbdf3d05bddab746dc4950c7d2939fc255b20ab777b7d1b6056b6970e163d21aa9498f3c8faae734fffec9240003c3f8377c307f5efdc54032f9c8a0d67f93419690c831c742a7160e8954b71132500d8914ca16761b4dc4ab68a72a2efb11b40cd15f8488b35f8d71f9bc0089b51cba2c3f13203ead1311e7ee8b91fd495bcd930e1b575093ffb6f0f66918962cc44c03514ecc9907c4dce823df0e293cbb92651fcc5e043fc6dbe65f2f7ca37760ed597ad590d556f174e2cdf3803f74d965b14a5ef1d0f30e18ce5516c817cf11c3bc51db1acc22073cf56ff1faf1d4aab8c2bd761b445fa8f9eb97b48f24b3f4eedb04eecc45a5e46896c6512083452e91f77361a1464dfc39696f6636c36e11b988d0dc963d4881d77fcf15612d0e0584f2f49ef44ec94be31f261e918d10cbbb42c58f12c1dd7fc4857a1ce1bfe1e38a6a42aea0c73132e334ea1fb6e37a03857c90d3be3b338e2f04110d379e9f3877d5bcbbe810134ad09c51d309b5e387138a10aa34b63831c263f3ea76d37d1782007fb5af43a7144003a6ac5984853012c2332a16551c2056c8c68784c74c02c2ecf1a078517629a8885f80ea92d2fa202b1b565bfa7c1f3122be99d45037ae6f848a450b6f1087f81c8c8a3d891e7fe4add020ac077bd14927aca1e1cb46997244aadd9d7ee0314063fc44734e04e3b72e26b70ad928b4c333c0bb81d8b4bdfbc5e1cc1378785b64a96ea337427214cd363848c2eb4a317695e29cac5bdd7ae90a0918ea6aea7679f6f20c076e181cb659dee078d9d7670a38dd6c7ddf60c567460ae9dcc65f1241c92e471f0655859d3b1f43126d080c5e6f7df072ed0fb71190a5049a512e969dcc70679ee2cd80c4674da6babf3b826b2bae6328a8294f0530202087ce518779b10d5543fde66ad53b5241e1edcd2c631ff63505ce996536dce95e4e5e4075035b0caa31c09002b7e8f8a2bdd5a6ce6920123009ef2c8d04c2f8cf0e0f71e4d878bac6301fac8c99372b3d429746019fe10fff4c006be6126c520e992d4c196b8b9003b8073e0656fd22a5ba3e665041fa3538f2a5491de9b17195933fcc37fa8a6f2e4a110443696cf62bd0bfc5d8880f1df19f1ed1e9670fa2d66777e4f82569730c085992774d01c2d11f59612f8b1ca962db9889a1dbaf24496c8b8ae00f4722954d58f2be6bb1c88fc61bc5e975be0a3ba7a9997e5b9181c1a8801526317b6227310a0c0c000ae85fdc8d3483d0b6c08ad3b7d780fa8a7696c5e0fd18e62d0ef1375bbb2f1eb3b714079a10e6a379bacd064690f2dd34cf274abfbc230b843bcc8c4d4de79660a32a58c73c564185aeb619ba28df4c2e31b7ea515c22ced421fdedba093e24d0b54f7c66ebf38e684eb1a64cbd5655ae39a5ad6f2b8f7f73a944edcda2697bacef3ad1947994116003cdac442bdff70ae2a85fa18fb2d4572fa0ebbed81da47a98ea4ba626db603a76a7921ac22eb6dbb0c9997c230c8d9672f576992887596b3213cbbf647f378c431e3f5cece0943d20f74b4218285eecfb988815a2854044187b3642cc416d3e22ad73df77aff41e8af789f0992b56a1fad75d92bdc5f028c5a9387b9c18b3c2110bc04faa42ed04e3409b458fe57d8298c69eb7f9fcff9be4b20f39bc626fc3be1f092cff1149a1e660378f68184151e892a2e22d33f39d840bda527fdeae5451fef69cfc6d67e1a62bee8e2422c4156ec273a4d7d725c22a92a632ef2074d575dafcb89b5ac0bada501eda6ca7ff8c9412a65a094315cae8da5d29c1e344411d29e948b4bbb56a1f1087195e179abe71766051619600e98feeec6d807bccd3590d29296562fdc249961cecb2e4f063d7ec0942038370b1ba01becf13473b674d0b451c422d189d8ca4d930167bb6f0dcd17e1e73d6819fc497d2548b8a79d0089619403cedee0e8517f1b3a94d1e4500b660c4faf99c39670e6313a1164d535847ab2b231c0f9b193f2fdbfaf865da5ca907b85bd35d2e28d485d4cfacad23cb262dda569e3d7cddc43019a6ccbeb10fc657e52fa10b5bd6b48ccd22b44c66b3c0be24af17377bfc739f45d2856845e303baf77ca0f23b5323961fd549dcdda24487b83ce0957a27152a52c0875f81d9398b70d7808b3227bacde6eeb4ad9756750c2ea02d908588d96df4e7001517586bf5c1eba739e398993989c567ab1b7fd46585c06c15cb6c19a335346de0d9e2a50f725c4de50bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h9ce4b70d5ff7f2051eb58cf3e7e2064e2323fd71c3085fd975bd6c9f8bd3adf74d41d5e34e1355564b13d44cf7ba6ba75f0d386c8da7db6d779aab69a0e0afae35483771db3cf66ba42d20cbca1b7bc385ceff910a9c38a2e7bf6857a0bbbb94141909333c63840f5010a056eeaaecee59bef299f1978f9533b35a098957953af8a0515e8caac1f2ec98c397f47625db236a98eb078f97bf94f257ac1cbb7a673db27df750db21313a6d4ad5c27fd93a78747205b2ea49e9feedb0e6449bfe727b87352515b40b75f37a3bd28561ba1309986035a55e0720cc15c1c668af94b8f204ae172ab08b4f899ba42e5a3d76e14db55a71e072ef33163103457128f0a97a95b7d496a3a8780d4c70b1c25873d752d0c24a931b57720d2d83822717fb95fc4ec18ffa08aea721f7feb54d454123417d263543c290f76a4ec7f5ec96f481eff769eb9529392d7f3b4e7f7cf0b95a350efd0832ce92873f9b15c404f94fc2f3de5d49bf1571db4b776da268b7762d15f7be4007cb3adc55f2f59260c92e0973fccfddf7262e125c0ab30dbb72a671fdcabc432466d4e7e7ccb46a1da63a0df609b2fb7995d5601fecf1f49a7d4c08b6bca35c69c2adc9a63424fbfa1f2ce23d18d8ce6c8a0814a98ae367e589b241aeb4ceabac41a62dd0dbbcfbaee58aa66a30a54b7354185c409ad5003bf5936c0aa9ef622d7c72f4b4754a85ae8e8e242b3065de933224afe0466f34b8ceec91df63e5bec81f88273c8ec2e463323a35fcddc01dd40ed3b781a55dae5dcbc8043ddfb0b5a9cf553f29859002904897e08d02f0c723be3716a59f6523c09da8e453c7536bd7439154bee87edae859344a09bb5be651cf3b743ca7308c6595b2a93064d6532a54c336cd522eb5c2f8d748fb835ad747858235a43494279d695ab6f1da76ed23a9711d4352270558ebad712d0c1a15b650fd5b342743efeae6fad179e5ddae376b243c72928ec6c148f531b0462a78520b265ba370a1c9e6d0bbd204132e89b0c890f112c08d6a83e3afbcb8e5623095169587cd268e4e21ca3143c206e33d21975c44db7d03057b64f778fdc3a40a5aca9fb8c32645a21dfc8cca2dc08cc9234754b9b2ed216de00577ce1ae2b1f9e3166dc13c34da652137296200c85fc462ce263fe0ba20be64f574ade3ac56b7b947d95069bdd163ec0ffdbf956832fa4dc48071a2beb8ab51f95b9a77736c51fc6d89f32d2310c52a100ee11be33c48d8dbc744de288c04a56ed4f1e4870315787abe3eb4bed5fa40f3631da1b2d5ec2350d1f9ca000d5178ecc8d1b269f589c136fdea0885eb4e9285cbb6405b4c8db939b801c211b2403ab7530ed7e8840fd16b642c844cf4bbed4d55c8d86b2218c0d24d85e98c2f5c4b1e0d72add1d1d4393ac6250cc966b5a0113233e54be5991985c9f17a58d6fc96b59c879b2a0e3bbc4619ed271c3d353a71ec252edef17a8cda1dea8040625438170d50cc771e2bd5f2aad2bcfbc442c16ca96eb76301cb53f4a58d3ec788aa491de19f1b6020dc29d1a445a1be2d0e50ae7e69e21408f1ecc3b503da0e4e740e6969bce32b47458fececcddaae377ef7ff4995169dba26cdd2c43e971ff031d7537edf993d818cc6dec381470459c9c2dfaa3d84d31695366f68cb5135166e4488eb8971abcb86c6b5cc5e56e2d4b7179fc0a243183634178afc2fea24824fb06d1180d1465de05208168a79c655ab413034a87d4cdc2041a1010b254213423872848b4256af39f725b0a97786b71019e051e188ad8b195d39381770d186efd4a9a53f444804426a5c2477b850b62e22ebcb3216805081d293c683918ca8635d43d9d4828c830725e37c0f4485fea6fd1458f4e65014faf177879b0d4b4a823459cdf56a167d8e8f2c4d000e5d8622e1e0f7f7d738c52e7fc5d107a496d889c57cd1dc34dff5ccbc38f8ee45d836079a95963c72aba88e22e27dd952c35f5a0ec5a4201a45147116e6e9c92953a74f3cd427bec183fe8765f1aa359d53f4b3f03f96d160c4f7f8bedb75b84b43c6a2b479f1090fbec1fca51d753e229fa6bfcce0a4cd991277644b06001a87257c8302b594f81dfb3f37464baf83060bbc744bbf53e1321f4e2b9a755fdd74d91c63c9c87566d0de80161848fb2d840e00fd4a0ec45dc3fcc5fc5a94c0ad85361448f4efb7cd82b44003597f57b2a52f47dee6a9bd15694cb75fcec3b0296f2337e11e83d744b1a02a979dd14fd18e89fe94ba536c5d9e7633b437f8d7038f0c12d1a8c830394f02060260447367cbe397076f5daea5e37ef35620cb3a195c4ea2173a1dc52993d17db5b3e25685a20e915cd7be3f693c8e96c8e2e42cc7db137e6d8388e2eca67db5daac417f1eab6f4a83965f2c8c5f482383757a8de1ff74917e3be4b7fe8e5578854d3f725ca138516bff7d4c8defe271489fca11fd86ce15429276727b9d0e2beab6eb12aa8638c3e7c48e3db4424330f6e4316064fcd04c35bf018f54079065cccfe10e4e58510d9b8d81993394b02789b6b283beee013eb67d2e616dc96a3e521111da6f245d51c8e9c709242d7dc058dfee0f831936b814ae55ecee2c11c98123e37b759fb943202f0b66ab436d8dd0f472c75f15a8ee280693a57bb3d7716142b19860eeebcbffe9e326413c09799c84efe52488c337dcd06797203d5b75998b15aa793819a60753cb034410cd28e8f22e6e6512302830de4aa579a8de72dc3c75a7c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbb0f31ebe3938ca069ed6f46d772d229d0822817af45704841a973df06fe058375556cd442eca2b5d8e74669a34cc77607fabf1d85d1180599810334d277d20bace5d3e2cecc9f610a629b1ab4268822d3752bab29915f7a768eb441e3ed40768f2226a4135f8ab844244385ae701c2be8ee27d1836c2540704858416f9dce7eef1168b567bf3b8a1edcc1aed34d64a264dc238efc59d0c1f54273c411bb33e637c1410b140ee1b4027edaf52626188d0bd20402840e65891bb3aa1922d9e650ff42671c0af98c9c76bd377feb9e4ad00e2ebf9a250841c554fe03a1b1bb381b76017f803e042d9ab8414cf51355c97823bf307ab83752a77be61bfda1ad0271ab885e675d86fa1d4f44c2bdc7d2b089519fb3f379e1b957f258b845de6591f9563f8d52af0b19c4cd52ac1458d3d55066c44506da5edabc9681280c41c5cd57c106d3d9db71c478bd011e8558bf331f7e070932a3e733c8dc31a3fc88b2dce8b02704139a313f475405ef54cc33dd3b20189a42c8ebfab334ba44dcfd2a011a4ea33d369453963d755d303f884b9515138c23db17f987a257d9dbc1cd2a70b386fdc4b3b56aadb7336d6b4c7dfb935913d77e5ab55422216b5cef096c21a24bc964403825d6ab310336d3bebf522afe5f9fa97f12c2f59e8ef90481b6134da43e2718f8a4d55a409e4d4b132209a0aad9218f5014e5373f46da376cb580491fdbdbf7f5d9bf2351b960c317cf2d3218c8bd695546d7ccec3e556c36da55b20f6b8e4e8cad3efba8e7dc6c0aa1ca63579ade97d7cb8df18d4bff81da8c491e52fc73c0d141e66e5ec57a8f2597647453547eb17533bfeaac9f7799fd4d90e13a8ee04fb4f9a0ba1044d17fd96308407c93279714bb3493e57af87db9d1e9b1a5b173a76dc72a692f661615b23adb732e9eeb7e5928d8efe19dac8ccf91d1860c7a02ccdbc17068c215e51a103e426fc677d305a3c3367ee98355c31e0cd7acd8cfe02a2cf8f809bdb4519e4fedb9c48f6705d0702aef2ccf507c5fff5ed53956e2785674192718502f1f5784e99d7d94912a6bd513e5d8feab406f46366c3f81af190850b2b4c4db6aa4f16a669d4f4419a1cb17d48f1b5dcf896f5dbc51bae84ed51d311eab0f2373f172199d6ef8c07f624d517e39bffd246a580be758d6d7bc2f27c29db9b646e4a293f829e49fa215e06f1bad4648f74b34fde6b38fa034a8b2f5e497dd5f54660d05ad61a29f2b56e8da6854d41dca8a550064274456154f597c08895b1ade187a07f36e13b3b9b88e1174b1db6321106851d4502072171e31b2b31d1191006e8e3ae611055dc3580a32f9ea2428b225d7ef3898f55f93a6e9e389d27ab433fa544a2d089a3639e66fb643160d9fda33ff0d32c43d53dccee14ab73d85f03334dc7bc114b14ad2f317db0901cb91a228782f1604fd3d58495023bd4fdacd44498dbfd652d21aee9951a8dfca2c6a611619f88a5dec4ca0fc80e8cdc0eb2f1fd9771ba471726bd32ea762329e660970f1b0a0924bef17c219280c61461258555a8b6ee698ad2dea693529c7fad52b26b872fbba3337614bded4282b5b3cee3c72133461f606cebc61833e7e938dd13abfa4eade2ac4e8f12406c39f70783f38064b08e614415a755f9c9119ed6ed8834707bca2d6031526bba262c815bba9f5ecae9aca4c697ca0dc089ec4b020c28716c6ddc2ce480cf575032da202774433ea8dec3ebb99e1b1635f090767a431e33939c54586d75317d5e15f398b7e8a681b583b0e727c71d68433b59ef2527aa240c22fd71f438b5403f718eb9a0bf1915b147b604a666107ec8c7250867481827b663b95255f84e2b88b83d0d057df098e1c53263793381b6f9dfbf883434593d62b0a2095bd0008ee8b464e8150679c839e0e777c116d7ca5a9d7db81bcd556680dbff271e05c45f80e4ce53fa75463eabc1bd3de83fda078434b1b622087b858b296515bddc3c92aa8c78b3474ceac3c894afe45270b51e902dc6081a26599a133dd0cb24d10696696150d93c2e01e2240d4af40a0830cda7fc869200cf247e5d082b9acd99f6c1285f95f5c9070f3c22eb1585b8ac261a46f7d275580feb194d40343d9add8c88c313b2347aaedf8fc64dd4b7136f360edad1ec10cde9c97fd225f7a0371b5d8fb00b009aba53576436035db9cb8eba07cb930bbec863651b422163b1384a7b27919037ebae5e8fe268171d5ae1f81442b745347687f8152f674a3f066111caa352966564032fa4e5329fbac7dc7e53a13df788d6183374aaeea6e9eb7a2a909e065fd81645a8b5b4c2b05eac0c7d53a94a4c9096551058a8f60e5ef14f5dd3b1cdadeab9b3bf01177d93ce769d9d47b02802fad9e2aaf03f12315339cc2a57834705a488e1d7a9900b2b828798996eae0d8c2536d4d2f659dcddeef2c61cca82703a601e037ad83202942c3739ef493d332635d7052d93cb8aa67fd221cb1f658bf3779e628de9d2176c64b2ca865925810069ff2c5479b76a28e6e0365e4f1111ca55c42b257270e84bc8a8e216bf216e591b64db8317389df94c81022abdf3e53d2bf761e4e0ce6c29c5ce628ec25607693f4ecd1311d63f56b5c38fa53e8ac281730570550f74ffb8b5785d0b6583d5a635b382d8f59f2fcbb6395b0d8e488d17e7bb992979f1160ed2d827f43d106f795eb2741d1ad9a8e44ef02b32bfeaf5296fb48cf5078e4e4cac146dd37d8b1a0a21ff0862fc0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h186b80dd70c9566d44823efaf13a7de8abe85e8029104354c6d72d1447a5e59b59862daf65bc0a60b923141b895c2b5d8424d0d6bf9e0edb06a0becd41669af926a27fb33b72f2653ca2a3744ccb7d80771bb5b5ef30024995c5132e2eb429e8d9286510014890639269562fff1503ebab26c4b8001d7b203d1c8ae5a4187b5db221e0f5eda59456bad8532ffd9449f8878d0613b31e4a41f8a62d8f66998fa6f822e22ecf8d941708fdf13f35abd93b40398e8165670c1d1502b0ad599f74656a78539303df1bb8a72382bd65773272f456589aaa19b32e227891aaa627ec1c827654a9f408a5f79735ff7ea45474430a95c2de1fc0b1b14f7202bf41ec5719d77a6848511905606a2358cf4550f19cd7a2b460d326054ab61e8470cee17f8a15c91556f20b1b535436566fdf060a9a868d9cfab7561ab917704a120c19e603b6a50754d46ca615329a29b2148346d726940d045d55aeae308bdd00c0da0a16c9e425bd4027fffba17289cfbb8865614016fe1cee3e375f025693f0b1f6978413f4162d7e4013da1c583645fc2791c5170bfdf350c000ad602d58924b0a6ebf4899ac346e32f6fa30e44faeaa2c6a6247eaa3518e096283150204c23ef6758ccf4cd67078357f395f4aff6259e9cdb0a0158fbf898da0918f29ab8cab14a926c5f345b65be789efbfd6864b80445f8629c01d9f87697920957fa0e2a341331adbbb98b9c8b83941c1f2e2525b521248e8e8dfd0e2ecfc3e3ef454c430ce27793fb0e81aa0bcb5fa2aaf06334b1c8f9ff3600b557deb6fe50cd45fedf2ce624b68f2ce845267824847d4cc8b8617b9aa84ac6054c304ba91f2a068daf2f54ad27ff924309132ea21746bf8c753cda43069ea6aaf34c7a13906572e5b51e5c0b587d5870c0703053d25da1b01bcbd70bbc9b615870f955491aa998abbbadf302c57ce24298a0ab3b8dbefba91a791d34bf0327a3ffc49b52259a480c16815002c3c3a9cba9ad7a7c3defc77cf055ff44ef0d82fac08032bbc19a8427edcc134ddb5fc3d4c8fbd9939229d5f0fb868c2ac6d4435c7047bf1f5c7c94e4626262a77ac811f20da4f8be931a426c3cc54d8b51bd43ec4ce5648fc7d95be65d574e07130246dd569e6eeed33a422e8c3d57fc5056c0cdf1de7aec4a52f437893dce723a92d61557ded330085620742a07e1dceac6964f839ab193af2c5798076c0120de82e30a0e27a0cbf6766ba8bed32adccfb3eef731f71be32c7f97c0024471f861cedb716ff16b993bd018e73597cfea1b4337a80393a059d59f14f497ff01256f6a3a20b83db84bd488235649d87c3917cd125121ee2a0bee26b69a127e9799a714942757a5ed678ab0a5cd115afce574eb23ed8fd11d76fb33e209289426d55fe30042140a6f3650a9949165871e5795fe7c6b595d93369054b66630481dbc68881507519553d3438de8a29981f426dc55106c3a9cd7f84d6bbf30031033eaeb25f01256e4b19c6af233ca4eda2bca3cfc714be5973598dd28f38f9c646a6da9951d09475241147567b551b97590fd2dc2402ab4e2872b553ba2fec2c84c238cb39f8d2b8a7fa8fcf7502ffb94047c17cab93c973ed5b296f5add903bd593c28261101cb608fcdb30e43d25bc02e2e6bbe152e0d7fac08b2f0d308854450f72988758b3129d3e5234a4d525a525c319fe47d3c5bb9734fcebc21db00ade9753154c2becd7e31e85a7ea2909fa385fa1a919c417cb66cd290f15cf1f6e8f22d6a28872958debe745ad0436b2e9f750f2fc6e6f4b4a344161cc632ccec061aa170f0e42f855f3ca9fd6dd01a6067836fed1b8a4d0b9c6b782b11047e72f27ba18d5ee3956c2032ab14961a169f2a93e5bb9f04a4532f1d995d9e5533dbc576428f62a43d92440bb8416973220d3c980fe8344ca21c23bab6093cde3cc6b31cb5fe771a9238ae5bf0cb557233650d9db80ab70b278bdff4f0dc2d0ed7f71d096c4dfec8c7d75ada61e732ea9f00d42cdffcd8eb1f4fa797117024ffb0ee8f42e0066b695816bfbf34b9cc193f01c9e004fb6df75294460103fcb89545a2a12a10101900cc18a3434f04d73c1f0351eabcaca853de83ab9b5c55faf5a8568f88a148de96e3b1b1f938d5b21988397ef65711bdf547d5d54c5cdaa5e82b369654e602fc8cf285a595997bb435d88fce3b9e91b0d1e922d81922bb7d96b5f05904bf787c0f6f8c2aa2fb3db7a98f2d564e56417e6b70774eb6befaf97925e9636ac9726f9869ccc266f95631d2092090b8f759571516b3becdbe7b6d0a42d8009f3f22684d1da97923da95437df0e9e37c23aa7ab056287e05da9aa1076bd2e5efdd9bf766dc6d758fdf88a052659e827fb60c7dc70def5caa67b0a301c33af750a051e13863aafd637a22c7258e06c04559127c541433c967922662ae7d71a8a7652071882bb413b7f0556031afc3bcee3b22ac183e807777b0872637ad996955b77a01bf2e28620ae6b06a6a826ceb84e100519aa50abfd46dd153266aae7f8026b01e51992b10b960c858bf197663eff6ee011403abb4c0b6ddaabf3c71fd5471a1d7b7938a47c25c4aaddc9cb0bc54308eafb5376b171c34f56bfe52bc98b8795ae7b8130f099902709e3b9201c778d3ea3512b71063069580caa91df98e9c8aec03d9c0e147526b26ace8a9b4f0f04f9dadc3ed96c7e7ede5cfb98c1d4a002b26faf144f387cb03bb45d2917752a460a2a967496b097be2a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'he64accac29127068c21842b84a22d80841068e702081408c8c91a9b4af06cfa928d24c7b8792b39beb1d54788a32071785f63bd2ec63b8c36d6dc02bdc4282a556b537627d41700ca4f1ea1bf2a437bd52bdca8b76fda08c7dadb8b28e9ca102886393c4e63eae678aa5e09a1caa5e0d3425c1dbe622e0f112e021eeefca3cc1b842a78d8d3288447969f0425eac37ac469ad012a73ca5576d22ec909a464b255ddd88e91dc015286632da957b4e02b904f7a9516f488f7a2185d1aebbd9a6a3f8ab56494ee57a812fe926fa7811f95c6eb13e629a6a325bca92800e4519618dbaa34e7a73ff8ce5c70109a8b71b83e806c5e21bee85923db17293e4ee53d2ad6d6a4ec9ca9a7a9ebf79d9ec17b9bfafa19e3612edcb9e124fe09c9a6045c4a51acf7aebf536d315b6f6c84c223aee1f689d5740fc23d70eec0def42c70d8acc3abe19b6135001e94223a5488a32ab54d17a253976c323b01213befe0663984585dabe54523e7ccf79ed9bf8de027c2628e2cfd0e88d35e33213b6ef52a2d81373a62a3abe8746f47230d276bd8e50933701c1cfa6637f0ff2c32b87860ab2e5c440c13e7ef044acf1a1ccdf0d8f70a942f71f019c7e1ce4883ac7302a143f5faf40edc621fe3a18d702cc5a0c3854ca2be99c846e253f40bda9a119630d804c7d3d183c9b666dfe4706b5a967a0802e4b00cb083f7de8fd93e4b65af6f2294a9aab76f4cfd263bbda5eb0d416ae073220ec01d6962082b3a6efbdb6d2f40c9b4df665903641a5c21aca2adf1605962d11246ba45658c752dac3b250e4e7ba1d04a053fc28d61a2ae83b1acc6a7ab758954b94050736e3bf265887ac9ac25ddf63bcd4295f33ec5fe8033300c9a7527ea0100f32e1be5b1dd34642588bf2517e6ba52399f9216476f24b89d11a8985f1d7f728c10916bf8bb145aa26124d97fde272fb3af15a322dc83b658a69a964d201211c97808753047c45216e66ad39ba8abd2b6856321e638c5a7472fa3748e647228aa5155d4814e31dfd988b900dca48b4c88e9a1ce870b0ec9d6c168e6767d6638a3d86857f282ac87acada4215236fcfccb766770a4b8e2263cebdd89da6c90a94e1e55d8d3158cfdcac11a87f555b2f4a556a79b98695311dc657bd15fb0b995544c6e8a8993558d735ebd52f32269e2736795052d05c0d9412cdea3a07a126cf9d92631786d66c4910190748e5707bffc3e6cb03f850abbfc8ce5564bfaa10065da6d5b419cbe7e470e84e51ac0aaa2d441342b75e0cd20e3c2edd4b8757932a40bf4dcb34e787dfbe1af00e369aea198fb6691e7ba72de81208b2eb11f0c2b729b55e73133fd1aed2475cdf4c1a41288fbb68cd01436426a2002b66c5434b0c1ab5af448c61e1de6366d2386f9a6ebb02ede7f00941eb6791e76b6f8734b4aa46dd7619bb28cfb70a2e4ba12805317790250f38b3aefb0fba6a077c367159e5fa9c1636d6d4e4ae199380f3135b3c1b750453da11ed7ef824a9aa0ca22c24024d97cd455cc242aa9be56e23e16ef439453aff0c919f4f40a51c4721c8b8afdb2d9678dadbaff87693f66ed3aa676cc9d911c115fcdcb85d35ae50985b4a30c07a3816dfb319629027cf41653c81d73769c7f84d6b1fd9c392018a71f88fc08ec0a1f0ebc7b20fdbb1ab5afafed9d8366f7f7462f480975448e0dab49af8c5316a0caf1a0ee30fc24bd5fa7ca53a0d5ccc9ba859bdf424b474ab5001325742bd5b48b1350e5ebf85e0477e400d5eeee9a7831f999f60eb860ca1a309a0b3685add5c25e44f63888ba5895aa39e7040fa002da1b6707718ffc61de6c11faf3883e8a8db6096b4aff6a852aa38b0bb16b2d850de57c4c5c636b22250bf1932783cbb7a9be950fbeb79a29983ac4b719917587d3586ab53653be65b0e3c30db46c562a391eab746e88b08ba9b489fd244c08c45739b6f26ea20fc87b18e54cbb816ed2c911717fc438fd8af66316a01fb80c72e9ae3c16fd6dd1c5e4790b03fa035b6b86ed2c3d0b9f3bca84a36edcc7d14c0c91b07735270da0e3541ce2b7a5a3761c633a44101b81f94b5365820136978df0e4b55413697beabc969bdb5fc7381481935317d719f0737b0ad5d5ce262e15689ae4a4c8ce912c13599a23516b58c9e0e465db8db67cf1f33754554433eb8d1e24d6441b4c81cd1f72f8dafb738f87754b7626d634337b46de9544eda4b627849ac01b448052ad2d8c6364c90e95558d53a49aca84c27966d2949446f1a8231b6caa0424a19a5ada5677dd4bbeee8e4ef07828d5d0a3f5a3ec85aa692ac8a01581169a379890ec8472af5ed6196449b24b87ed78f5486c6b1d5e5f85700ffadb4f9068aba988982f8479ecd21b9ec8938e3a9ea91d7a44234c27ebb1983a3e6d89ceae198ee9876008bbf8ceb5492f99fea30d2dbc346e279e59c25131e329578975f6473a32a630800ea158896d683fab728bece0c2c0968ab67c26782deba009f575a20ac95270cac15765a9a3d4e58b112bc8f9279f02330f45bd04659133fc218eeb056caee2d409a09049e5cb3a79b16aa9eff2f8094be8e5ca50dca7931ea1dfd771a30c07a7d4731f69c46530c5c456163522c10ea24e51671d12b3838bba602ad857980e8dd60c368fde79afa06a84d5a9b0499948ffa77faabdf93a56aaece15516b62780d793d6133ffe5d6024a875820d4653b9d6bb38da1246fafd3ed34408f5437a249e4558dc15593cdb7a0b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hb21a9edc1ad7ca6f3678d08161ea567655481a6bc12f7644ee7739e0799d0860fc95b5099e46f0edd1a70917f849e04f578faa5d54fa778730103956361e39b67df56895db83debafc08cac781e1f54833399d9f9fc392975e3ba88b6bea53c046f3550cc14e66dcc98964e6346fc441fd13de6805d7a319b19893b8c73c12813bda64a6b858c8afbfc33150fe4fa2de9e15480ac522a7d82e77c466f417f81a272d207b91103dd0721a019cdff433ce9d4921ac95db195ef8842807fb5daa203c13c378f54f50c1b8dafe4cc50f31281f836166eaeef81cfb6808ce38068e2aca073cb79c3a9214b3e8274e063a34fa05ee5a2c8b905aa34e157f025ee9a022454300ff91a45f71f89a43eded0f673a58a66ac6944e281dcb5483a8f4a30ca670ff34b7f20a1c7f8dc9535bd299198f985b9316c39283626bc330724ba5cd5aba478fb933918ceb4ee3a546c0a72e467024b70d7cccbde77ee1b5de7dede984de428f069a9a014d4fbfe445b67cdc8b7ee8d0ef744a5d5149033ffe7dda82782d6829daf3291609d0fa9d553359bcc6b4ac3cc223b6555102b261da96da9fb99ae13421f7cb86d1333bbb3ffb37c93b8e15cc8e2a21a2135a730aa395bd9e620ccd9a7632d0837d48ec59a6717cd4cd5d8eac3254231cd99c874584c340ebc544a8e15081ebb318a4f2cc8e3ed63c8e895712a2b16fb47c72e8f508e05d4ff6e12551f03cdf2608fbbd3374cc8da35a373da213e488d85a49a9aab18960de3efedafa3bfb5b0f4cd2c6cd3a94ddd2933b17a6c83bf07f3e516d6322fc86c7d68aa644530ccddc1458868a8e161200ea5b93b138f6b5caac2ff9626e5e9540f6676fa61068fdad140166814f4817e8d6e84176e973b16a29d859512802dadc9907d4ae3b846db15b9cc8242c0d816619bbe5ef379a4f4fd8bbc9d55882d9d7ad5614c0f7673da5886b026b571a47ee839207a0d195d866b37f7a1ba5cbcd4750232db0f1bf4e4f16bfcf474ad0b9fc02ac6de5ff9acf3a01253f0c67159e11017aa3eebac4326cc87d0c75aa0bd59c4f1c560e644c32e43d280c161c9eb00a39b4ee71921757313db77847bef6f69f80d78c6ec3a30641ba48a0325a4cd7a89f28e3346b2d9d865cfac73308fa131b33207fff31d61847ab0ce01d42088862f8908f4d42e55ca2c091bf6e4d01755a236c9bc162933607e4c2f54dd178ab70bd7870c182da423ae1d75739a1da8ea57f5822e56a2809aa8c59517627516e337528f1636c0d935fe5c2e0d9a6b6b368b25ebb40a0163157419403659456c5b6de7202a1a3499467b27ca0ab664032092af7994e7a37b577d802672f53fa228ea20455082abfd485b8d9fa4d45b95ec4d1e8bb64bcf196963581726541a95e106a760cdbf8fdbb8327c95cda588ecc680b85826ca333d79990004436f935fe593d390b04277c9d41abeab8c3872b46016e7e8d016aea0ec2baf3a0cf4df45682aeb135750df630382d54c91fe04f216f4168191743df1ea88dbd98bd1150eb9109c569745202d1ac8d7a41779f85d4354f8d1321eac646fe720dda896fafaa2a84ba5855db41478d1671c0f1cc7ae77a6f4a30deebc0c6ad1ec79f58b7000be58cba8752cac7613e804ac95d2fdaf0c292fdf5ef9d56481032627c1c1d9ab9a41dcde51ab3d6c77ff086cbcb3401200d6e814f10ba9957174dd17714586f534764bc725f5ecc68c55ed7b809371b426a69a96b474ecfdc83cf8f1906979b2f4b9533c4976f139ae4956032fffedb3a4b470d7bcec05a83dfffd3c932087894495ad5dcc3f4185bc9e9036ae5732b706324b9e3e843ff624fb737ff11c8a32ad0fa7f6c86b91a33fdeed883af629aa44a3aaf6525eda73a80460774c978c54f24c0926ecf174ece658c910b3ebf1f06fb210d63ba2e89b2f263c27856d90390ccf8fa2ac83a761b32586b33e7267823f3fe570b5ac787ff7be4543738a415b85cec6f2251cd1a606f1ca77604f233771d40b31e70e10f23c386abd33fda7a04f39a98a9c07adb7fb95fe45fe799cf300dafcf3a7030a48695edde3053fb8b94ab73466e75e8066ab761c09796392f9496714f859df884678c390a93a0ad90d726884877904366dd65fa5828719fd6d5c1d9ece07d645f23ee39f6e8f357c29c0499a3679b4bfab5f6ae096c90b322eeb172aa609d967efb83bf57567bcaa10b5d0f41f65587d4bc34a13f8f6f516976eff4131e943f95013e49c0207c6302bcdd400b572041b03c5fa95b4855d03313d4eb120c52b7dc2d83eb2436e522b711079309c7c4a2c1d6f60bd3eb3e5243504fdd988de65ce6c69da576a1b2535265e06f67107a6d2f2157ccbbb4fe4eb906f5b80d1d14634e0a16fe93fb1e337abfae200f6ade7bb47d93b751291e1ab00595f9cd82fa25e220eaf4fb907d3ca300bd590355e0ace0bdd9a7ac831f65dce637392f1e761510f48f0b9f553dae02afd91aae1a009b9d96e19473d245401564592ada9beaace666d9a3bb12ce69d5bb0da8dbd1f236ff9ef827efbe90c17af23c4f6be5514f4add524cc9ec701e8c32415cef52c6925f57e0de525d969323e8abe170a9123417a8429ab5f830e8386e7774e983f84cd9d091ba21ea49b0e1f92370e5e3aa16ea2fdcb4d1a2ef3e7699ed3c4830e26f57ba80073773c3e46f5fcd5909fa5efcdf5ca94b3ef9e58aebc331822f98101f5d903d80eef5d1852329708485980567f23262bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hbafae66521acda4cb65ecc7f039375ab5115f687c17b018366c91be26fecd16cbb124e7b97e8b0ed9fcd81a8b93a9cb14ac597e93be24e71a0e5721d74bfc368b675ce826564b1c965e14730a1e7a7772348e194dc04cd6ad72a7e7f52e9843a3e9f8e3e6f58d69dd3092dc57ce525c25e6e4e4ff8be11f482c7f8a0261fb3fbc8849e0a6e70fd0d4db896e685a6bebfd62299efdefc7d89570ec3aa34de2ae9a78881d242aa6945f0ed77912b272a570863fa0c2e23971c3db499f57669a100c962d25d52fdc00ef55482775eeb06cea579394c7a39f1e27a20afeb5070d19ac84abff9c0686af59fac092856276c412c2212a0599d35ab915fd49a608e2fa676614d27a9be3818a0abe9910669f211ab30cf48395584a4e96b123ccc92dd578ca4a967e68fa089df616a873f99319191c668251d0f30880263adccdcab8b07691d12d93109d2bd68e5d2aedf5edf589369a9715c5d1b21e302e7a38013765712d44cf9f603e249b852fddcfc920295759f45193516589a2bab4d484e2b6bed015bb34e51257e095162e71dade43ea82acdcbdb3d2da87c85475caadd36e778fccbaf4974acef0137bc959a7a2d38ee5af9460d864a564403df6fcf1d9364734cc764fd6a70d87d7ed53b0d78ea593e1e5384e58a56d9cd29cbdfe4f1812787d36a5dfdaf54c326278c1ac1540ed496ca47af6205e91058f7953bbe001670a6fb54df028d824c83549598f47d858b07b04b814666eebdfa967c5402d242e20432328fc20613de1b625904aca7caff5db7184d5989101c72750f160ad73ef4026cedc364a954edac6b245e0d81170b90e0b21cd9a0dbb4d24f083be6971bfd8f1bc7433446569ac024a194ea31cffb60298cd8fafda14984d925c5340c4366307d124cdfda66c6fef1828a8ff68f616dac50ad6da8cae493ed376fe8030dc7e76afe5eb6d46482927c08f5f52d5388b283ba00649f5b066516c8f2d7bb9bca38190765ffbb0629a5a8e2307066cb21224b28ed4b026213257882ff361d0e7b3000adfe01d6f5fbe9e57a055099db30e21a9baeae0073d3f86ae487088450b069fc87a7e9d148940d75a68198f3ec53dca36d496eb99c127af1bd8edbcc757651ee20b9784ff7a953bc5553af9fbb08351fa68a70bc96803889d7f1d88ab9db1eb75ec9dfe6a1b21067a5d6fba4dda7d6bbcfb1225008e2dd830d83e73ac2fdd3519f33a652b8b6143e7322834ef6c9b011c00a800d00d1286de97b85a606b5473007a05c81b0e45183798760f1a7ea21eae2f0241e82dba75042630e258eb5ac183299d32b1fdc8bfdb513be0c5c2dc9bde0da3d8f7464e02dfca997c7339ce5786420a9bac6f95d5f5f521597acf834fa5633fe6dd267056b7e45f95c35c8af2b52f00771f266d2f9a1efd21aaaffeec696695d427f89061b5758b324d121716b37492c340764b87490d6ddee9d380686a9ebe53af83b29791fc9ef81066e7eceb1c03110e253d56a5e7d46973ee2daffdbe72c7dd0a4612997664d4f583e09a014df36d9cae69977482cac23dc22aeacfe4aed2f0c5a8f93470f775bda546203cc1cc286dbe5ec7ec916ceff666fb87bc579a8e1fe0d82d9eced2c66f2879908366a87b6dda020b9ad545ce9524f6c34ab99c40a03a178c7bf399e0be6935aaaddd015fd8c5c0e281bb33a55d5c1cb4d442078f0ddb622c261bb489ca722bebfadbb536b9eb605290f623ba62ebf2de9cca1bec1e39333d3de22a428dbad53c1a111c1d91aa438f610945c49ccd03b7d567e1bccb8c5e99d75336aa0b2adddc40f70fd358689a1fa4d7417238b39d5ba00b4aab59807a614dfa47d10adda30bb72417cd2ec057f2421922318dacbbc7dfb6061c64ff126ae3bc57741cee0d491119bd69faad06bd61d8a90614e7944e030c4ccf67fec0c4f8ad7a2a5987d325ed0b12927fee3583d428f90e90679d51d60d821cfb1cb2d66519e192c926da4aa1fc900a467b0a9aac35905716b0fe4bc83ab89d5f31b696c7c691ad9841097c65430255c0a5050d3e2d4dd1193ae157959c901d875a3d846c30545ab434c39a98b285c0c457bb309614e3b1300ef8bb6dfdd9bc56687dd7e9c13ebea7a6ca6dbaaa6b6f832510c85d23f442daa84c5871777b340d00815ee10dd3a96540dc947da07a3b96658aa333c33d6fb6948c9c9c982205a4477a5dada642662d7dfd217865891871cdefea238c6fd91b65f522e1082d7a920c3c83e1dd86e109063077f6a979e382b55f41264f0e10ba858161bdd2ed7a7e1d16cfaa99244e0b2acf4248e99300eab178ba949c2f51856028f4f975ad664c5e97899f9e8c6a81e4d172257b6eb9f59f57887090ba1bb5ae92d82a8d7ae6512aae0e5b90fe94b2be63009b631264c9f73aa86a28923c04e1d8f42292109374c162ebcbadb6b6e4d31d45d8dd21b714b00610eb230014b0f30537914076104a1abf926d9ee43e181c5af4bb2c956e0f654995f58e107b9577fe2f90ed59ac656e280106ff548f386565d75d11dcbb07500adaebf230f4ec4d47edc51ef0329a33c67921c52ef61ccb68a96ab8cd5c37ef876b21ac7da992254d7895b922e3043d65c2c644b535b8e24762ba38c1f10585cba2264a3e4451f4b4688dd8116e94a2cafc0bf2e727d6240bd95791c3de33c4fc9aecc4a50849d7060458dfd7754eabb8ed72f1e8ef43a52eb064b794c01e1733b0ead9b4d91b55bbc98732ecb5eacab4b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h50d7852c1c3bc7e2729677bcab91b01620ffe777038fe220aa3c332b6820755602dccc69697b14a2b3118a43b260af270df82909f388512989ecda3b3fe447421017faad87976c7385075035751d07f264eb9cb10ebf31a261c51a1f2e1716ed585894a47b01455738990fb37b55e9edc88a2fc4986920290ba1610551e5df78692d46daded6eaab92a11152eb07379a8489086e715ed67e383b2ac39d821e0408af324a0208ef70c704822b912d6cf4454a78297257b1fca331ab32673fab13d9c64afbabb17302dcbf1e6f6887d2fb604c4f2630951df488745130d897e1d0c56d71cce3d029013bee23006b3cc07418c5676bc05532fecdd422a71a91af79da51f42bfe7d6eafd4383b5c1a8727d1a7b429bb5496675ee3ece212e6e60dfca04fbbf34d952f5aa3f82ed3ebef36ca7f97d552fadefc198348f7fa169b447977c0c07fd67e914174e3d534b69d153b6807141c5ab43c27b2fade5d3943272d6a44cb4789be772b86d18769c21037997d1b3564f90cd52334464e5e44d0ac84b62bc47ea2445897d44c7c328746ab989a868c894756d0843fa0770acddce22d96cb5482307cada9067c806d7af06814e91357f99f947a71df085526f898392c4dec3946d22f3e9b9910d6d67cf0fee59e7d792ba5435bab9a31c9d82d0782332fe3b3d9369665842d73799eb6426e086e76cd3a404458cb42a30e2feba1c8339836dbd81837979e52a3def748a8eb6d014c99aa9f273022695810c547a6cbe877564a108029fae4ae3db0eeee06e4d2ba1ff7bcf567a39243f5c5a3415e3501791e30ec92fcddf3f217d97ec3b3782e0dc7bf67a019dd0387026089b54f3a6d7c1dc7e379424b180e2c131667c89e3d839e07d7bad6781fd452264d19e50d4fbbdbaca25bfec369569e847608cacea07446b7ccbd75af0307c43fd64fa73a2f246a53eaa520737e4c97e6d4f9d0994ed75eae94117ffbf5f1c200d4f266b4dcd7dfaf3a08f5b935bfb495f532360a45588fb0e2fa9a8478d9ceb1d62689afdcd3d1af17c720f540a48872d0ba0b58c791f1b3267553e6eea9c5a702dbbe304dd01ed1345349f38df89179786d69ae30883e30e9c6ad60aadf2f01864da850d7fe4134283ad0595782c103961029d01e7941ac21ca078591ef6f2eda7b0fff4e430f9ad8568c5e6c9cd3d4b64f8218736a10034da87eecc7d339664d9d8c092eb55b031f3afe6d6890afbc0ba0abaf538639f8651b4bba5823db891942ae915084f5e5e18b4c449556f602cb86956e2ca846e2fd513a61f38c3bf9843566223fd22c99c425fc75e78019c74b6561d1e6e75d073331a5f4182e21d6d3bf00e2f2549cadfae3444aa8808e94d61a0eb98eb4228cbeb297ccf929ad536a37c6fcca2cc93b3d372f773f5b5f2ec5cf9f5af910264e99afb984b38c74d24669da27495ec0c137133f4ef40fd621cb5811e8a9b6b4de1a6e8b59bce253cc4e2b84da6c62504ee83285fb99e5b6ec09031176fa29f60392ae5d83a56271e6607a43e1ff830502bc51128b06e35292b2807a34735d6fc6e39a0774f99df4e0690e81c857feb980e50a882ba98ba5264bb4f6c81db93cf72c37b51d3a0edac297e55488b07d45e01e216c72e719119cb9c2634146e037092ab096db34986ca6b2d0a47642e5921e7b1d6b9bdfcfa4bf0ca37903644b76cbb56dd15c8c12e66501e7419c9e4de63fd024c12b5a80e3fa144d9530a68acb2b959827935f59c4421850610da61bd2c7ccfe30db94c07ac7c655d10965eb86c5c026e2fc2df534b3f43d11a50c696469bcc1ffd07d35bec1582ec662346f405fceb72e0e416a5ef89f6968aae23cab51432449dd43a52e9d940d3e96a6a0ed7e0d61a9f062239748657dff03f504ab2127501628e832f2b324aa5717339a4fd6158b32cf1b942306312f450814990479363b174aaad07c0a525394ae98e19c34330c60ccd38ea255c7a772afa2c5860308f28dcb439e4cdd2368bc9143d22ce8000536fac0ceaeea9129ece4157153d77c1a09948e067376b91f032f20c0d2405b0479846497eb73255fe08ae002c6464925a51c1023bca533a2659ac7e62ca5d0014b52c2221bc03ec853620631db8c52b25298560681f3f9a8ecfc237d6d103da372c1ef4fb153d79aade647efdf9f8a0d5dd51fd5f05474eb4c70632601ab45143f1f2892994b527ff064dda9b4a83dcb4675d36190a0da5a6195c5b2f889467debb5fe941ef4598d188a754937e85300ce00bb7a788f8762dec251f1862f5ea997a76d48e83d86036943a6fbf566d39ceb2eed17db07f24554c71d5bda8192a8eeee95783c2d4f05ea46455ce3afea1837ac9530be6844ea5baffa5e5fb17623e22445937999a4bf3241656c265266c5c44dad82cd0365781a27415485c16fa0aadf53acd6d3abe95f0a08cf18c520121b6fb45336d4b331a35afca29ff4039f666513674bdfd195d9dcc5865b77d2cfe747a7ce6e35320543ee530eacce4a0df23cdb472d39da4f728e858d3dcbb1ff2bf01c194478ef7c3e07dd44bd02d2a171aadfa488887a31e43622e9dbd19ddd037ee01221a4fdbca718b95b1ddf6e775fb565bec37ca6bc5e9c503bf4fc6cc5fd26f85a822621373861f71d8e047b4dbee6998259905587e418639a078b5815411b4fba08c09f7e9ec9f94747d383597535992fa6f85e056e59d3d4fe8301add36a63dde5b23c4ad26ec6dbcdef0ec5452c5c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'hf2eede874f84766030764393865b8ad7e5b7762177086e2b815f7086c5bc5babf92e28a7da2e962cfd5251140480d64922425bc9b13f5c32c4981f035ae57eb3a3e8abf2b7f8d4afa42cadbf5f8cad9a5e0118b5718cc932697c7fcb2c30fee9d6289427b45d9a4a05ade5c732bfc5b0d4569cb4657dbd307489dfec8ef6f8fe521cd6cf141575fc643ddf2f3306a39f83049855fd3b9050c391fdd2978b7ea35252ec236b21a6e6ea6c675564eff03e667f566d9afcbc18ba42d3428ceba88d761d3c20eab50f80076b47f573b87e26bdfdf76a13e84e3c036f744c36f0d2ddd45ea13b5c81c80e6e8d8ee4f3bf3ce4f243c66b613132c4ba89f5a94c598e83438501749b80d6da31239d2286cb9bdb59a501c9fa0097a30b2f49241543b51728e201a35263e118ad9508fa175e70cf8094811057704da8cbc91c37578fde28eb24c36f5019b0a3502e58881c845cdcbf8bbc90418167b8216148d9b81efbabb855448b42387054f329ca718810d7b12c390d0ad77ef50e111dee88d0164d162af6657a40942ebb46926f23d448eb20ce6a1a58ad167422155f1197f3b44f08808e818a2f6c7ac507735837fc26b8391231fa56c1c52f03f819ace5ee957d2b4cc9e4a0ba40b0ffa68b75b89b1ae9fdffff7da07ce8641b07fd8cc7a4c1e2439f7ed37f8e1b212fac91e97fdde41a51b6d9d5110f78f207ddb391d4d50e1ab278a9d04fb58a3b54411f1700d092513ade57d9de02819976086b5011469fdc730c0f78167c961dc4ab1c0ad526400bcae8ff067def75e5e4a2ef5f5ab06789adfda5c08fc8467f207c3de5584b34b253bbeab7ada3546a5f0b5b784d6e565da1ad35d78f0332f0a87ba792f352cef7f5270094b06bc8d90ccd51e89c307bb85fc45cf5a18cf13bea0babdd2f669976f07fe4928d14b20fbe72b4bbff7bd2c14fed89a8ca3b8225996a8d01cea04147cee4ce839889256fd2d122aca15c62f8c50823d3908cefaee6fe99ef44e918e6445a6ec582ceea5d7df9301716bff8e3ad014dfe6a72395da6bece38bb6a2cf00607accb7bd27fdd5b133e51e65ec36e7f44cbb1594b13e6ae8f3e026b61a9a5603f41c01b501484c43843162a8eadfef1839eee2f6aa3cb7e751f5169445ea29aae03edb351871df127c75fe940c8a854abe193857f5da87cd476bb921b4037639e7007dfbd14ab4541b59109400fae5a78eb32e59ccab4fc36197e0d6f45d37cc1f7a02b99da4b073e66f82b064edc7f5c519e254290ec682c9990b29cf538e048a56bbb9ddab1f3b0eaeae06dc659262e47f01430310e61585d7dcbc544b2d7ab9e3d967ee42015dd63a470a4ef890ee151d12d69fc7d6d078582fb1d1a392129fd1856b2c1d5f57b8df11c83433064dda1d3461e4c9d78f5eb3ef95e4d6efed3ea90372f41aba9be188cb8f6f9d6eb0a34a7b5e84a7805b272cd9a8d5ace960461262d19e13b4e0879088b91e43a56bf38ea05dd70a25ab86c1fc02b7c550a7fc1dda0f63e5b5fb2c515ef64f7ec75e8d796125a4bf8b783b6c891e8d21b2edd282f4b736991d23800c4e52745ee38be57d45b012babaa5476b4dc23cceb9cbba7d0ae1285e8551b4eb593337785130115fa9901e3790601e2a10284e75d01982a4bd51e56c26525fe77c827148493281dc183e4058e24fa5eb80d7c6b53dde95809447440f36f2c9b9168d9a44dced51e2910a8ba8076ea5ddfaf00ab635d3acac67e9349bf387721dd017d23b86777e479bdf364c3a3ed0bc83b65ec429fd838f6120fc37ef43ebf3a95bfc54e997e0970b0483e5fe4f44e47ae17f5013a2d717ba4d9cb6c87160c56e365dd54a75b334b32097a80ece6ea1135146ed006fbaac462c484d3fe1af8f75620150773cc55329bed38fb814950f6303c95dea45de0e739a9fe5fa2ebab0a667332c01cdec7001ce3273c912bddef7187254dc7b86ddfbf7c620914028ffe5d0f8351e1cfdd3179fb17cb6b0c6e8a6c995ad04e1d7ef9b896a6159dbd5b94927bd69ec2d8fe0e1e23bcacc20e91436508ae4a1dabc2ccc532ff1429d8b17737fad9b061f191395cae510ec76c03cb384ed1f25e4f6dddf9f60bbc62437bf413658e9426953bbc9a4c1b53268ef19b5e69f67b6aa35375255945edd56458156364fce9e50bb62fdd54398ca822482d17afd7b867e58c175a1d6cd5bf7eea646e0c3d3405a669533c8565712e6feaf2845092b167251f1bbab761cbaf7e6767d6d2edf283e0907d105af71ab9731a2ca389d9426f9524c49d8291999c77e70e83c5eabbd448df95ad260832bbfc2c8b9473339cef66e12936bcf97c6e4b5f6ccd94bd713b7328279eb1393031fd794b762288e68fe0964bd952b8c0ef7c7a1132e25235c1ce67a55a0397b95da952f07cd2f13f981cd831fa2286c4bd47506467cab2f35d4123bcbc10063b4590f8518ee45bed0a8d66e3fe62bb32d87230ba33e2e2ab4efa3726c54ea3d538ccbbb3a2e33d9f34862d2002e8cd4e4425922c6ac6a53d2198dac24fe6b54b61bfca23387eaa6b4b45ac173c43ceeb36bf0661aed136b8a80410b06b51eb85627953dad3372caf6084677f2bfb54b39e4c3691bd34d3df3d0389b39af83a887706b702dd3c21497e2d1bd914031adc88e662cecae1d09afc01b05106aea0abd1161d844d7d641f6161b109aff55ed9b2aa14e5684b7d1783dbadbe302f794bfd6e65f1b1522d87efbfbb6e2a1e6375ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 15552'h951ecb9eebf38f23aae99298747f2cf99609177370ca9f63fcdf81002891c904b9efcaa9c7c0b09fa5b7a2d44a46562469c819f6912074c194ebf503b091bd620daade7eed0ffcf6f21999b92b037c7b2490ac68f9fb9e9dba9bbbda3a52bd00218b8a2e592f5e9e19d4b37078923f1d7535a82077f170769fec4f03802d623e0b56c0f2859b3e988e047c0daac92ab4ee2bff0bfc9128b64074658b187a805ad35e93da45de4496c444d1db5993c39893a247d31277d62aea6cae5e08cef439ac0c788413e5d6a26c775460cecfadc5c517657e9b26e4b464cfe800bbd5c11b12ca47f4ca20e0277b0f8a2c8d3282baa164f0c0b130d325d5c7a15f6625d1371ec847077a42be9cf9bd820f734fb46c43b1999aec7f883980cc6e83c0ceee6e41d405c416de07868cd4846e536296d9242bf49575d359eb0a4d138712a0261933ab8bcfe497e0616de250ab98d2de0ac651fdfa67c0102878fb1e8eaed47e312a948a65e601016868a6416f4990437af3046ef8db5ea759454635f19540dc7a6237600f6efec48c46511725bbc027c859cec7efd59b04e55cb858e52c326001fd176c0c87ae75991024de6a4d91ec686c40be187dc896d913858ad6471cff74b207c58861f86c4c673a1758e21a8f45ab43e5a53710772ea614ca9339a5e65f971f7e45c75e5b297a14ebe7daaf8c6018ceaad2cacf0c51426e2a9770b333a9339940cab988da976936bffa79407c0aeaf1feca77b94456446581fe881c1c3e576ae389762ae414c68e2b0fbb90aa22cc59ac33bc0aa2b803891b18847190478f589d8af6755180b90310e54b49be42a725a1d97bbf018cb387bd57f6a6c1f142a807147805e15c2881b8f7c4a34504e0bbd8b128e48641e9e829ce371244e8e047f84e8d172d634be09d12c26620f7d94510046817946ef81ddadc9d56a16a0e0fee6456fdff6d9e2139337b873af3c90dd19ef16f4b6b795288cb052c5d053c0e5bb29c9b9012707dfd0d687febcf95f20b6eb1100cbf92dbcd4ec6fccb543c4d8e5da286096934eb698554d1a27c69b09c139da15eb0e92e3f02b6da1e5f95edccdf937759006854d7d1039b83da2b8079c3576b6ba6bb6be821ca3ae752517d2f3cdff49d7c188ca5e14c55b8b72693313a9f0aac23b62f8b39d6bdf6179eb957760f2a249fd3f74003c3dfa876906dae2480ec5234bceef5d3616efda4533f8b7e727d86707e44a59684d5ebd2e96020860365d74e175359260b4db1039efb777882a71996067c6391e9960c764a18be697223b023428ce1a1f6b481fdfec1aaf4e487b1ef99375ab7e77e5b7e7dfa01804dce50218b16c6f67555f2f314e254748fb04a583cb8653b997a35ab382fa88cb2bb9e551f0a8413a6a14b15f752814818a6dbf872d7454150e8d9ad28b72e5acb05ec2f401e065cf6e0936faa5666d6c5da5ea70f1a62eef01d8abdfcc44933d0599f6c72190ba6138695f5a5e209ae4af0e65780dc84ddc85ccc9faa2eecc4cbdfd78502fa6e8a9c3149fb26f9fdaa0a2d032aa4cb5898df1362569fe91d35390fdff30e553cac46c704c2be05bd57614f7efd62471a58a15f83e43e593f8c3fbe379bef13d17ec29e5f1b823a87c71f20137be4929efed08d23f25d49ff7cac7eeda1837645ad3acb9d5432025f6ee9240ebc73c9871c98844727bda76b046324f9154e3910dfbf43f2aeae712d0385b6a9cb3119c59bcb393644c323d1ebdb9e8431b8633b3001d8c4fab63cbbe6d80421e828ef9d00cf1dce96054276de89f5d1f16ac59101ff38b5beeba5342c40ff6372a866c7d8cb87f6e10760b3d461cf0b65383327771f0274edfd4dad4f7d36045b25f09f2b530e1a3fa093de16f58a620c80cff9cc6eae1ff7fd1cee477383eda184006ae987a63377a19c09e045b00bb254a0b2547fa846f0b184baf7927ddb969d619acdbe296a94b7b643d875430c78511f7d2526e35b83f970d3a5837d9ad99385f8fa435d6ede1bc62c4ee9fb06ad96c93d42a1b2cc7b739d977e284053d826484846436dcc12e833c889ac7d8dc4caa2372ae3df8b92f79c36d92a05b8005f5cd8719927c13b4772d0318c27c8457aceba54e81d7cf4f2fae8a77517501af859a260832dff1b1e2b19e827036263c94ef463f2c66a489e43b51067e838d5346082561242400d68b37391b61bc5a167a0be252d3aa55ba8cf3bee5824fb3ce3681fbfea5fec9b389170933ba47b87f38801c2b07c4fede80e2d0fcfda554d2edb38e63c7aadc4c257a49c0dc3b2d71e3577e628db412add6ae823254036b5c599f670c6889ebc51f49ec9577b417f6cd5ea972824080aa8fbe3dc593062b5828514e9929b1e7d511e0443d5c2ed33ab09a6305ad738d2f37c260c4517d74a08e0d896d726efed6631c2aa80823d99710f1f610e43736e83d711f3a0dce28a22aa917a27ec7efcb0359d743958e9eba389d2ad33521739d7c398b0f866260e8eb09a5a76a022ded9a0ea99b81378317d537ff6350c712e83b3e261d2fa11e7a75bf7ddd289857da5dfbe57cd0ce16d4189daa31354f6605334c4e4e307d8c746977f5e2705521981f34edb3c8a97c4775ef7035e3ee6e0f0c412da43adc2b7ad21f30c61e0f0de7d2ddeef44054aac8244662fd63061b3de8dccd3c8ae5fc986930ff4a0901b6981e158fa774dc2ec66d7796bd56f2a701ab28830365b866e18b673ff189e0bfe4c25e923de107f93;
        #1
        $finish();
    end
endmodule
