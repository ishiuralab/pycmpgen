module testbench();
    reg [22:0] src0;
    reg [22:0] src1;
    reg [22:0] src2;
    reg [22:0] src3;
    reg [22:0] src4;
    reg [22:0] src5;
    reg [22:0] src6;
    reg [22:0] src7;
    reg [22:0] src8;
    reg [22:0] src9;
    reg [22:0] src10;
    reg [22:0] src11;
    reg [22:0] src12;
    reg [22:0] src13;
    reg [22:0] src14;
    reg [22:0] src15;
    reg [22:0] src16;
    reg [22:0] src17;
    reg [22:0] src18;
    reg [22:0] src19;
    reg [22:0] src20;
    reg [22:0] src21;
    reg [22:0] src22;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [27:0] srcsum;
    wire [27:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6c247de462564487de29c3fcc499097cc2307efb3ff8c57d14bb7236627024e697107a3edea27f8355f3f75a326434e97fd9b58b6c923efc77b8a14d303cd52877a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2a2860e51f5f0a2809f32f91dc2250a5efe8ac64b451afd709102d00b12b62235e21195b2232b0bf936697d58b3caa286031d9e1d79402b7f8b024704063a913c1ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h104f40a7b60cd555000961f313e0310530163efd018e31783122e294b64c8cb3acd1f5ad16ccd641ce60a6af9ecbb97c1ba293515a3dce021120fb8c0b4188c2cc4f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a3695fa790b83740bff1fc43eb9594d488bbbe64ecdda87ad84b56a18f795215221bbb4b97b42884ab8d199358c8a11ff623d5d2c59bf6fbd05356b695ba0362384;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e75bc9e863faf27053af7e1d533dac3e773f1f7fc9a4ee3615472828d4627795f8ae5ac21f7a3bb57f1d18c2a92c3e7c35b81d4ffd469bbf2527cad4ab23d793ba3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bc3386924510f0756dbf83afd9bffead95e0f8333b1a1a506b13bd234a0e75a83f3bdac29ae906c6c0f6183816736c07aa79aa27e9e6dd4dc6f3e4b74bdc87a5b0a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e2e3c443a5d5d90be1a9858a622a5ee92f73845bbaa78d97dec4cc84b82f9c3ee877dacf81d964f14922bd5f1c761f6c09d6aa60aad41afd3df92f60d47d18c6c93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8721b5401766cdac134062da497d6df6baaf44434adf39f99e76fbad69ae1a2eda5e02b7b575383d54cb13591a52c2470dc41ab5a644d2e5cbb1665c2b3726e8e7e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e27997bbd3179cfb77825d2db7f7142ebaf198bc26b49dcf269875bee2b289547d9d5f819dd27de8b8c72e1adf2548748e069de089b6be7b8581e9dde0bb86462545;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a47d806c045960f53290d4129284ce2ebd74ebd14a9d720c8036a635ba0b3ced359752fe40f33b568ac257b223b9d113ef30442f22553fe882b34bd001085d454772;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143bcdeb6e37cd79bd5779b7eff43af2038a635c707643c90976f06b5c2a3d8f749fe939e8dc818c26ab482ca2504ad857d1d6eca98726c88c2675836ddc7011a6bb3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3ba6aedd229e8e72a0a42af79b82cfb220150596d01b9a4cbc5bf9de342e34c830832027e9494e5abbdfbbecea60caf1ec07a712710c668433c464cbbe76337a51c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha8e35842ec34efe1bb7f6a0473e70e74602cf58ba6db9ac8a6d263d99d769ac61a80534c933c6987d1ce2bec58a0caa7e1649733c8f1376a6f457e5e6f226391d66e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cb299accf0156628191ae0a27fc1ad2f681662280c8dfad432d22a50665b78092ed815116eec91d133dba52a3c96336ff49900fbe57f8b01922a50b23dedc371c181;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f5f6fa668e369876e017c163d2e2980dcb665f7e7b250f77002d3bcab6e5ccfa9473f16721d9e263a40264db157d4e7801bed3254a3510c946c2ae58009029de97b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1053d1974c3d11455211983dc5379aca758ed982e9c40186cde4714972bb8ba7621cf9e938d3e922e6546a491e8ad0603b3918657b656395c226c3f51eab78b1cef61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d00a8795fd99c47ddd9965d90d5889d0a80deb8dc8ec90002191c1ca1ba8a7d595f3eafdd9a5b8a3ee52f576c7df3537bb11fad4d30818bcc6665c80a085c0228cc4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hacb14ca49d7f97f0da2bac31fdd7c951ff26a0d541f23087ae9fe36b166dfe6bef808b6c35a64f4077fac3dad1c0cfa3c1e1cad2d7895aeb8cbb28acf856ee793084;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab6b2795e99fcff9ea888ea55e7759332f3dbc8494fadda2e40cd45374326f21af7f33c1d3aad853e3a983c46e128e2f1e47ee8dad672aedbb2ed87229ccfaafe6e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfec41e0800f8954ee3f2105d570eacb0bdfa5725d3434f1313046b523030f6fa2f73dc5ce669332c50f15452699b5dfc029c5e938d97cc0107234b7a1d9362f04a72;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbeae4dd72190c53ae70097baf6821fa66e937b55a9a51f377a4d47e4793ecb5caf609de92e0c19f0f3e202baf1756de5573780ea80d4398c0c8bc5e187cd5bc79d53;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5045e0d41e89c14d7d0f16cc23087c7e3b82fc98bb6daa1c9f32e700d2a61206eace2fa912cc00b3a38d465fba47e987c64d2bc2d038a94b9d6d4fd665b5147548a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbacd926b80dd48ddfd631434a5296ee9a05e264d0e9a15456130eae15ac874c8302023ad57a95d43a89a9a251716bbeacb4f346f244406cfbf67f45316d7b0c1c94;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6af84728aa9ef261451096208107773f05ed4d1962cebc9c7ca122817926bfc314fcad464f7d9d01c266699d70cf6580fe0d819b33e68ab0afa6166e7de06181a911;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d0c20790c5694e28362b31e3018653335e7c069a6f9544365f5e5d451ad94e6d38ae4d7ca31a0d30938f893c64700139a75e981a07bd3ad3fbcf77266aeee2ad0a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b8e70edfdc22d9975469603e921e6d3a99d3ab696de0253c6d07b02c2028384ed42b2f806c1b20705c9c22e8bb1e038b6e4f34594d1b180bbe87de8461201f7404f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6299d79508ca1ef207cfce6ec8a9c58398e9adae296574ccf597d56e92c9473ebc413e5ee50ea0173dc6aa47e0ce03fec8bbd41c03d60cd7224a93d18699a173a3c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d52a5a61810dee3d3903f4d3587f9cb71c65acc1553905a3a161f646d6fceea21698ce707857fce79a7dcb9a0e146a06e091a6a806d6f616f04d29c8468aca5a6c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c03706feca44d192148108b399d4f134bd60975788d806efde90359b577bbaaaa964f2ddcfe60a18a3799a7b1ddf0c0857158f72529c925531055f117abc4b93371;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hadb1bc5876f62e2fe0bd138ce23f494efc744e45b5323224aaef03afc36d6461d3ae958d7b18a1b93e7f1f7116fe3ce9060eb73d7472b201baf231023c3b6f0746f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h123475c66af4ce6a06499510433197de0fe3b518dc9577466339a1559e02d9dc806509f4e8e7170af5e211637ebce1b366a4d7e65c379bf610468dda3683f9339c5e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eaf2f7d35cb104783bb3f24b463a76b38c37de8b7276d85633545416196c50eccbd236ba914b1e5e51c63796536612e9b83ddf3eb3cd7accf10819c0996048bbb4e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e3ed78ab69e718124529da80ef3742bac283a925cd5ca4ef8fec30897eb3db9c04bfcbbbb8d29b9514ad1349b16ca09d1f711c267e69b1bb477bbc2c2b5091e88b17;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eadc141ffdb2ca5de4113d562879b5da1f1980bf62dc7efd742d15f4b9d74e389c0ea385c2bc94ec35212ae1b51102395dc5e5ee6ae100b0d03903c6c6831a03fdc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cce7049b9bfb2d42dd5e965d031be8f45de51d9c5a9d0b814b46a870dae8da842be0862ee3c47c3f93b9cf75887a065171e2147d74b295d2fa6cb4e5b5e09c226e77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c0f4c1ff86a396b296d696d538e944dbbeae2fb9631c55fffb92a4b38eb24151347541638fd68a7de6026b9c227588835ebe7f392fa59f2ca197eabe3aacef8420e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b9c2af858629c6c6fce25274cd6e6cd78eae799afbdd69e145f8ab9bf0f61e27b61a99e9da927ee2fd8823d7a36c99b55ecd3b951d0d9e38a4c16ace661f3367bcf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0055da2a1a57fd0a217a39798b6565c2cd1f9da8157abf07fcde7618384777501c8e6556c5144b675a6dcf2297753d79aa52ba1561ae59e08e9cc9135f2871cc9c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13ec49b4244f246d54423e0e7c9be8952a8f62f871d88fb371a414705106de5a4a6e24f648dbd932ec3178dc0618d3d1be5819dac684c3fea0aeb241735779dd47b73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a38fd069a6018dcd2ef3bf12f3d5ae704cb2e6fe0fa077b93a549984088d78cdb3e77ae049a33878c541f72b960ef51d6d869da5a9f6e58103794cede90f7e77b40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a859914ec3576834f72aab69aaa71437d5047c93c0fd1eaca1241c495065e6dac4ad17d0bfa0c43a0e0777c990bf0ed3a88c4ef94af5b20c1a5a613cf12bbbeba6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b6a15ceb0126b6373a95a17ae934d60229d2bfab7131137b43fd712ed23d5a0cd0494a2172aaf3aaec53da7370cedd6d90b881981c396c43a0242b70cc58043e38e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc62439190e79d56b75a2ff7fa7f799a8a3df69167c6f451d8f429a7b34f3fc505facce0c552c27516a6325233592410af3cceb6b1d38472a24dc8b32bda057f22489;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7dcc88ebe5733a263c1d5aec73e4f9791ae4da077678f4b9bd37d961e2d3c3b5a3845b057d2182eb782ba355b72f15b0e1019421cfadbe63aead5e83360722165569;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hff8e8fdf7cb4a58cdf89b4476251522e8095305b10c9a16d3903f19ca3f8f69ba1d04f41ac7d81051a0bde4032a0b720fd460687ae828aa7dcdab8485e25dbc89f9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc901e1f15777fe30736990792127ee71260212e8b5b57c68bb903d96f079427b89f6e2a21ae551c348133006b624991787a04454819426616d7fa4a53b4f490c0ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61e8edb43702345d5f44983d632447760f7052d012122248319772c3f56bd01c054fa4a67e402c0aa9ccb528559eb3e5fd45bcc3c991460bef770245f9186db9ec70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14212cdff77884a1ac35e4380d7582ce676f61077998d2b1099c3ddfa1f600c2bdcf6f36eacdd78b5862a749cebf60e2bd236949906ee06de2c54b736e1c620a4a6ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13b6e15dbb85e6209b95775aebd213ea3f0fec61a38d46aa37c8b0ea9e53d9c16f615dc8035117dbdeed9b78dd3cf624b01369f3130eb0f016cffcf8893bbdfc7a3b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5120ee6a213a83a302787e5fa4bdee3680b8610d7c06980067c34b493995327499bec79b505c688bcbc36f3d4da5cb05d081fceb90fe25ef9c59abe9256fb595b2f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1489225a4f30736f5df3f45c001fb17424f6604f7a8189256fbd6ba826d505c188e26d3cf6716926a3800ce5b743da1cefcd82c568489f126543ae49400c851cdddae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf5858ec7942649ece55d1edc9ddf582c8c0dfa28871dc4eeb7f447d2b8e363e6bcb5154b42a006f68258a5bca148d432a0608fdc3b9f0a21a14b2d658024f860caa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a66569a7b2165e06b2caff63ea8a707a95992a702690c240dbf21fcbf13fcad82e0c7fabf9e3e2671d63a5cfd9fbb6e105c305735767028853b4c147292de63318dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1585cedb24892471cb0c525a5dc366c7f0ebcfdf08866bd041a0b6791d864bf5d1b4aaa66d814cd91387c67c4fcb4a8472dc070eceb147aea13795ccb6363c0b431a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd53e651a418806c2d446eb3c1d96143e8a87bc5f3ba7a1cae1eedb0476690b1c36c7c3554aa74760b15433e8dbc1fe11a3e5ddd1d9697ac7d476ecd327b0d7724f5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'habb641f0703db9dcfff97f72781ce73c5273b8c3793af5de6000ea7c7fd8aff417acd938f864d1b2b66f53dc7fdadcb2a380fb8b5e3952b4391bcddc75b617484c6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c0f45988dacebf8193269533b01a8c51b67edad4dea55295ac3595bc33bf76d20cde9117f2f0a5b2884dae15e54e76a315e57909f64b58dd6239f3171ff739171c24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c6e6d74b155f966d9ef56f2f313529691f24c1a5ffd067a26d2473a6551c2b7e8545c0347a227954f73e2c721372f2319a694bb9820242abc85493f3241264b8a5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h75909f8eec66dfd2cab1795acc657068b8eb8de6701cdd63b02ae8af219cf45b24fc8b53be663c8859aa2cddb5fd861cf3eb84167a806debeba771716aa895727137;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf5bd84f77e8284c13cf605ea5e2d1831d4075b6ca468e445d1add2b8769890c70d2a67c84c21923f1a730e871753ce1b964cddaa5d0026c909ae96fe7bbdc7ecedc0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15fcf2c76ba0673830102df32935767aefdd2dd22d732e47bc1ee9820584d2bbc3931ba57e594e7c3ceae33a889f72c4549ea42638e5652d0a556e7d7e1a6ab3b35dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha2248b5ea945314d9118fc05c9f7a8804497b7e627702564842c9981fbac062435a316daa0da5a46abfeea36ca6f07f4dbefde6a00a11fd44ae031692c2c0e1349cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1711466451b212ff3851bc21a36fc8f51311ae8f06885d01d8b259405451a4c710da7e9502de3e938dfd11a5451f4d38a5c46766909342154b68a1ad2289b3acaf87b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8525164670dc9603ba5f4bfb490c474f29e3e86e701e0a6d307b865bb792e28957a94c1769a2fc7fd66265bdd4b678fac40a400b641e3109666e82c88088e11da8e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd651343a65116db2d755e5cbf2c51f4b0c27e4260f5f83b17f74f7d7f6b762360f7ce65fd7ae8e72873339bccd8ee568ff6a149dbacfc5042e1d975501c7621b7222;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cdefe0b2a66acfdefbfe2a630ececd5e6d0cb26c8274939281911ef4d8005f09ba0c6c45626bd6f34af0902aae012b1e3d13aef2c164da3174da4cb45b407f77835b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90c7b4a8660a33b821a96cd6c9b6b2f93cf368dcc21e09e7385fae532e54abcc4c5bdfa4b79c3803668265409275ecad23346af54f1501357419ddb0b43157b775ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha63fd7d6b2e3c2ff4ead88b90a27cae15d824be03e59458fd272a35cae1293e6a02dea76c7272aca9d6b95a4be2e31287779b8f9bb6d288b7f604f6fd219a87635e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ec7254f51d8e715a85913a8e6357fe58083cf783c0672101701ddfc8dc733e63b9c4b2111fd8135922d9cf08e3e3f012ae5e0a4d78f52782ba4ce3cad55a1be2ea3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a7d9be706f6ce8491914236be8545f9a98fc12eaccaa7747b1965b0bb12cdd99a29d213fcaf095419ce0c899f1cb3da2e8dba1b28514775680dbf907a2be786ca7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bfe874fd88c7d1d21dd46f806e569d03223f31c8f058ccb6ba4745df33f0f7a3170e049585182466220c89f44246801089fc5b5f7953154dab604f6f5fd015844043;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66c1dbab7cf5ca20eab0e0e6952b9ed610805024ae64ef34d702c556f5cbc9d356214d98da1dbcf7586796467b92267fd2f2ebe1e1e02e1bc2964cbb0eacc8bf8a02;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h46a0543a4248eced17858f7145c1849d9256ad203a98f6c68a8668c3f35dd023ba1f7971f39d8518bf3dd99a8d07233687982d3485106d1b57e1ac526fdb58e5fb85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h45e0fc74421b586a2ed8a1a169ab2c2b424067f751c0d6ca3ac1b7234c044aedd46df9503202a056838f6fc21d333e2ee6f583ebe0625290a0e730ebf99fd79bbf56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b96c81e90cc5c4f4c1a8081b70e7d32443e041b19a20fcb31b94a2bc9fc1c213c7fcc7a1a8750a6f350538c11ae57a95b3b2b3c0f475496bae71c594d3adfec3811;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e47f956e55ee0dbe80bc0fc60ae82187e5b35b604517a5ab44438317dd52983e117d653e7e1252a3a32a83d2da4ca2d642d4b7c73464b8552480c142c9b6255e23fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11eed927a3386ab7757c60cbba5cb591bd0c4670de1c49cc7b149daeb300dabda5a6134891b0dfb3795896b3b17ea978ae4ff8bc99fd900b89bb6060fb0f0bb1a28f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b87478f2cd467366dd3c4af28e6983fe2b9540872d6ba3d8e732a9e8eca050da800468d2e777a3940cab5cb2c6c2ab3d2ebe1f9706fbe0004f4ceef6d50c3d841ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67a8a92aa74ac93f68a8d147de24f947cc7e067824ae888091b130c736b1d43385648150c381ada58c69124e10085cb8fac847a323d94287667a16e2e5ba77001459;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h776eebf69fbc3370d5787cc06d649ed393d29e94ec119944da39c591dd8193860c947c8667d7a0d14d6b81544010634a1a0b90e5ff4a6c67f357cb4d71769835d3e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd2b4fc67211ffc701a8127d704b70f850306e3f9d8dc819e355970f3d6a78b6d55eb7a9132ffb73c2283cf97aa6d5f7827cefbb0a18d714ecc64b11aa2e06b2c4eed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he208af47ab3546c2e8fa6e0360c2f576fbd4c6511f10b9422debc3f382ece928809c1c0f15414f017569e2dd3a34828f7f8d953bf3143dda1b421dc860cefcaffe20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ba7133e1b794e3b1bc95b27a6c58343163a1b543e98a88c1abc499228e984cac625af2906935973d92c288abd7f0c08f0f7df6b344ea41ffd2218479fb063a3671bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48a34646ac8554b2f19e07cca3774666a7abe8c40d9f390e8427891b8ea222c7d975073518a55f10c94a22135f6b82be6b57efc64bbbadf8bf0af2d7a659a8de120f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17996a749fccca1e780cfd9d504ea71d350a8c0ba5f422685307acbfeca0b22248b60c109a1ccccee4d621f063b09cf26f9e5d0d67b9940bbd0dbdb6f5260aa7dcf11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194b0b1dde73ffff873b28e0a1b6889fc0e916339da1bd2e0a97f64483a2dc0efb6bc44b7e7e93f991a341260acdc68a8d52f14d97ee5dc37bb8dea946196b33f1932;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h678ce629dac30f2007773c9af745177ef317a7868c543f054ff059fa35e189a2357983d28ffdb88114bb6e99463eb9cdfdd8e960d708f1e5e542eda4e3f91073a3bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h116db170b1fc113cac5cee2418d9a4c7b0d913f00ceec0816417768bf7a356b8ad5e34e80ca6a424108631650390b82b3f0c922fa769f6c651731811421d88627c5e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1978a08d0cf4a0fb126fa007b7b5d5082cba4f390335a664f966931eed9b8b8ff94e6ccf08d8b3aa2e2a707fdfbd9a1f9c52b2bdfcbe384df053cf669440d581a6f98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h492d14dc56810b69bbcc6eda80c8869b475f43ceecb7c37d4d14f54dc1514ab92fdb30bdb922683181254c1cc4f0a95941f56242edf835e048b0b766bfd639ba0613;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143061bc075283e39ef2ae97041cbd124c470557082e38d1255993e5a7b901ae90b14511343ead38f02f1bb3d66a96c6676303aefdec2f1eacf9c4256b2e183bb7056;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61ca4e8dddf32ed72d2d6185c32c70bb229a792912c23e9d5a31a7c2860c5759fd8da19fc3d433f50b47fc26f42840fb1f27c3b7432435aa26192737362652f1ea55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bbd855450003d26cf1a1e7df71435a0e1d2d7fea745419d6d87135f3a6f77cb7c3784c361d513f81264f4b61735d3ccef8f766bab4c08f6d736d8301bc453367e679;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c6f9d8123e272555b3050a63a0f94953da7235ddd47d33c5be9021a350987258faa57dae703379098db343f3e316eef28b57915a266393d24b0a19c3156accae2dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb115c892bfb6ff9ac0a03e9cba602a0e20b85d8fdccf648d3a608f6fbda9d7762cdc0ffeb7e7b42a4b02f5bdafd9cc7e0e82d8e35cc51141bb0a2ff36e938e90e819;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12133efc8a667408e1e0c8db01812a38ead5d9c280604b57907faf53e7b370b2084e786739e6c4e1b8b4bf7c370c9a1a0b76a7e0397dcd926726a58b4a35dba953f0d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ce5fc6e7ba62eb70abc626d571847cac661f43c8ea51cc1f89641fef7d4df16ba78a2be5ad39d5c33ade667c946d2709bfadcf3372e35e65c6b65800feb0b90772f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b297bf73f1c85d44901f02d14f590b408b17c73612e951cfef0226467343702470c65b24151ed6825afc6c8f032720c7178e1e3b0f27f4217654944a45b4cf1f3e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbb33ace54d8407b3de47dcdd995fbaa347c15ee1ff0a2a2003ca43fc41d6e786c20967dddf7fb3eec4e8ec08f015a53ee2a51fe23a87f796998600b9776f4ee78b39;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h179a2f56be11ad204867919e9b971a07d7ed2e0319b4b46c25fb42b96844f6a59d48b71358ca3bbec0a841f698e24ae8fa2ecc070f709b3b0d5700ba59eb0372382af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b40bcd992d399bdff3ba1d11b55d9d0b190b3358bd7131756a84a4930cd7cf8433c69682e2363731473daf16233355a402739657d4f73ec540d263f897f0bc4fcfc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1553efdf0a7a96dde388f78c9c23d4e4864e37d492bdb76e5f559e3048e533657f35727b87427a024961d73f9fae41a3f5d2a591de9ce24b3e3772758ef4d324fd31b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193b07da704dfbd72621e40a19adce56dc4c60bdc558ce56b6cf58916d0dada295577ca5ad2dd5d63e87b9798af02a4738bed38fc229f603375140b7219dc09903dc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cebcfb4e3dd26093e0c5ae1e1f00a9d82768f50feb2d2a94dec75265b9ff1e70dedf9725ddcbaf300ee293ae52c56ee94c1f75799d5ecc61afd3ee643941abfb6612;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf61bbd81c48ba5e6ada79abda5571c817b3d2f8374c7a78efd3f58a0f9a152bce71a6769ccec633f4e8ac0f3b5399a5c4c51524fb00496869aee94631d972d9ae560;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6be5def2a3b12f93bf47d5f78169b2c75b23ba3c24c62e5582390fa735462e2c1cb81af1c8d263dba3a5f833420bb1d4d40fe81b2568ef240224a282ddc081b2401;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb598a3e40bc8f29ed5a9ec031ad6f03537a5c62cfec387b9ad6adc19bc22dc7e54ee7de0d9b0a0968ed870310d55edd8fa52d9eb10b1b2f38a03cb37180e3f5772b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9e1c7725df07e5d1e51e82b3087196f0d3e02f96a2a56c10cf506ec9519f9554f82872afdec5c9551763148b3e5e4faa129652aebdb90438a4dd824e01f1ec7fa198;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd1ab1077fe76527af470c0f7923d1d2f4218f64ec16f8e0c0c945b271894306512d40847b62f53a7eebe839486e83ccc8f04cd2e2369fd57e1c1ed17f862596b3db9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18fded58098b8c656e796c3444791a0bf991f9d956f95aca778db2b322d9d0899f85de080db9f06f06874303a37e2f09645a68d683ad73363fcea03e4989657a7391b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fe830d188b902f5ffac055b5aacb484f059a190d0ac202aed9d4b0968a4415be2ee82585975f4e19ed305bba719256d10b470c4e0da31d2d2a93ffaf0698f10e44c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ecb39de29877c534f2e1b10043ec249fac656ad1f431f90f2d911100603a668ed67a32bd08ceb0194e9f9c2084ea4753a1fc8ec6838b8126a5f9d68bfbdd0fbc931;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h321531fc734cce7bff6a303170b753c7e0776af7165065b34b11b9cc7f30c27fa9fb9730c4d5676fc878fc59d1be0a7b9e3177ea137f5e1d95a2b3dfd22ff234d422;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4421bc978857884ef338d5171f234c3890890921ad0462e3893932ed52864c883bbd28c80ac2c4378668fd4054deed48914fb4652736dbbb30e5add2e49c2fa09fe1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cef074b566f019eaae2a0287ced03537409a3bce8aa9491ae5f729ea07a13ba2f94606766b450e061b2cb06e9ffb9db1f93bdb7e89c5d58e77f9c8a00be1ee1c7d16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1913bb271fdace2290fe74aa664070c10cbe8f831ff76299c9461c95a3e684596cf0127d0cd5a23244c1f4ea52a5598f8a5500dd2efc2f48fc1574f64524eeeefead2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1387d24bf495da85c3f70194b36a6e83dd256ed8b3c08fb0fc5b858bafc29e376b376c686f16a126c061174d01dcb42d857cb1000681df6cae531f0170002720ab47a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cdb091ee6d49acac59566728df16555c8974bb2c42bab9ff102ac290139f189384269b2a2fa7647ec3211d8ebf58d9e40f05e16163fa4c25d9186b015f52d8d1fc89;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bb8009abfab5e3339db7426c4372a54063c57df44494a8542e5277795733810d836a701da185480ffb44c23a6d1ade7c333d016032fe5692fa59fd449f1f369276b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe53292fc6ace8e08aa0f59fda3a4f0cf3ae6023fead86518cc8f652cc2ed9715f092c4b2805312d08e43a1bb325ebaf265bce025a749700df6be474baf1eb0f6e6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he861854c675aae847eb09267fdd9394081691ac417a4483b52bdea8b743696e8978077de8178c7d851ca3fce1bd91d7718db300858d1fb5ade8235a1570ff4724ea9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h785312303e8cada9c98dea048efcf708100303aff934f503cf8ba0ffdc5432270219389736d27d574edc07140eade8a098c29a48f2081553dde42bf3e34a55c0dae6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7ba76e4d01972569398a7a128a006aa08740009b6753860cb053960d31e22ae4a5d5f9c26ac2604d2ba50a4c056011ac5f7c9cfcf29f0aed408f6546a3ef6ab094fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18a54c2a5d775707fe3a3da0c8bdc61c6d8f380e39eebac56ad88074645be47aeb84876ed43953db67ff8afab5149c6768f31cee4314fe68e40d82b55e86e9d17090b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb8b73b58734291a416522097b2bd50f4b913d94a8cbe16a2a3ff8b38f9fb6b88fdcdfa0105e567e8ce7cfcd239c66477a0e31edf77864d392ea0559b331309847a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a6e724a820ef17ac5af44ae60c6bb761ae2d46ac646e0566d06ba3a792b10d8730810b2d50c102a37ed34b38927e62f207bfa5a5106539d64ecb590ff7f846be74cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cba96ba3073c2bcadebc8bbda4ea32938ba9d651967683d0622309c2ffaf0933174e900f8f3eb0d316bb6246c3a602d2605f999eec56849f1b81f3afabb07cad9e3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he56de6147f59cec95402bba37110a3486922d828a72c6e2d714f09b36c22c9ad76d7a397b47bc5cd565dadce2778006219d759bfec8ca6c6453ea7ae2ae654df20a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd77135456bfc11a6c14cc1731022ca30da735be83d7cfde6aa8c929e859a0b5140ae58853a6e270657b46d5902f62c71c171f871a07ef42c7467308dd42bc10999f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa7d5e9d5ef0bf26d334bf3b64d9ec7369ff67083287ff6917c943e76b414b9be9da3e28e26be09455f53ec29d3fbf45b13998c46617eea3dbd8a76c11676f0528e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f199f91be838f0dee19eee62df5d4191f7bb3adf6a629f8895f110be670e7d39823014e90108f6e458a18abf01dbf52db14712ffc3a44599f39d2cb9ffad89f5998;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h76de9195c5ce66ee29016040c3056444f983f7b1e7bc95d924ed68190edb6fedc92a7a831b4f80e2bdd1265f4decf261f4a7379396568248344bc4c24a23f7e13ca3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h668cd390b26ac7e2e435fe8f801425231e0ee64ec120066c6eb4bc1cd3fa7db7fa8660663c471b3581dab13544d2131e6ede94f59baf7f29aa42114f82a7f37360d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf228d52f86f3965c509f643539980523d1de737b7fa61c18fd47b79ebf1d9a0a9b3aa3a8a8c0129c82ae8bbdf127defed773680483be0b50dbdaa0a7d2d815f2ac21;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h530230a1f6958d48f65cc71ca2064d135cddc690caf6da68cd4849a494f866b1cdc79ef711462022acdf361438ea383e5b4176296499175249374a6444274d04bda4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73ffe936f63b47c7f0bfd2bbde3c243e535f9c5e23965f1cfe105862557a7672666dc0e5b4257d0cd2f1e5b3d4884a0e5e2c6ee30e2070f2c78dce3705e729d971d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h541c4645267f04cb065983056eee338d1300968532f0cb23b2227cb8ec8e24fa1a872d7a34f9694a2976d9dc1e64861f5ab65dfcb5ea4a8521b6cb45b2ec226dacfe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1589652c9968a186326d47092daceb0630f251ab090544f06b19320d8a5191f114d06a2e7650b7547d9a1aaaeeb964d993eeb95c0879076a5c1151a61f5c4866eaa5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1008a6b45f2bcbcb7898ddcfbcefefa3e1b4ba147f2759b780d69bf7ce6d6cacd1ec1fd5197f57bba79974842a5a33cece459b2c180f524c1ba9d9bc51d5289afa131;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h32de9703fa057ec709a26712b137cfdf92754caae97e66ec63ccca9b3ed8596dde4d3e05bfec6f635d626d36cf786bd6b47a2f7fbdf09421595decba03131e8058e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8fbf9ddaf44f93fceec0262c222d7a2b1e0d13dc0811fcb474b4b82514d92e37271b78bed960c4198be1d6bac90cbbc6b114d25780c22eac8a1e5f127000319e95af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175f3dbb70a41af43f1b63df3c42ac98ee5847dd27d53a66f568b4e6a099b653f08a2214ccd2657de3d2d002bbcc4e7547ebcde8aac2db02e1f76da9605ea214e88f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11c677f5453eb52eea5db82ec25b96ed8935ec5b4e59c44ca2bb6532b52f54bd58ed3404e0d1688fa1950b2323341777def82a96ca763da260d14059d702e0fceabb8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1508c724953d7642601e5ed8d3e18887b8eb92ee95b65c27339de79afbd7544bafeb617b3bbdc8a37ce281b457ff16e490dbe6349cb98b1f7343cd3174b6861af64a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h897a6bab8135e36065c76e63062d688411ce132d785a509e492589e047846285d3b6fb3c773f10d684a802e6436ec58314e5851d2229cb1738397ec4dbd2c68bca2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ab1fe0cae0ccab059b31f70a64cf8610d7760e8c3521b37c746480540babd8535622ea08d85471e09155579b26507cc2e89b9431fe7c66008ca8d2ff2968e004b6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e26294569367a3f9857a9d484b8dde7af3872af8edc918bec339dae7e61d426475b2611cdd34409ed481acded483080e06ff3a28b5dcf33e26cb5b43cb74d6a995b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4d6d0f4921ddf5b953198fcd23cadf493059bf443a0479d25f918857e1edf7303011a44eb3ccc7ca18b92cfebe025ebb7efb74db17e2f273f5b7de7bb89ea698a92f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c1e4d9f0f64a2f9ff024c0cb306c8c597d2212900b4ab8ba7afbb579423c3d8963176cbaf371262fd6295c47e1376198d360b972b068de7c194287dc0aa1cadf9989;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4f685049541e762307498244483478f06fb8c0f8ccc8f744a93180e01f4cc0b9201926391715081d5806979fbae131cee505e0e622da13410d4eca99a219018098e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h147733802c8199f452f9708a93b10ec562ea4d4bb8549d90838be7dfbce97acb70182f6d49370aea95e827370ada281af96d2773ed36505c14f01fabac5d0c1b87e60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c936180445f6853e15ccd2b3dd0c8424c7a1ae5222ab802b6fc9842981795695650a21db401b687d6013b73e64bd2b4449a4acae2f23103a063e5cab196573071f9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11c462b787a2881c19ad1e59f73c38025df21478d26e00b5286beb5ac2d506dcc243c48ab44a2b1327c6e75550a3eaee631286b3ec7a7437b1b7ba408c88b7090b44e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba4c75a19ff68eeafa318395973dab9837dcaa2f6b11306c230d27f4e46e47ab8e45f6412e0906168bb47ece4c6e73749916a94d6702185c5bc4702cbdc8ac29cdde;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h45fc9fbeecde8a4ee1a8644223bc089017829cf99073cd97f2d1883e1dbb8a03d550541f9c18bb288089dc8a8ce00ef2384a97e3efa14bad273b0676c493ab9d682b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa128b29449137a608b0e85b7df114642f9b19f831749b4d32b10a6ec98d2608b665517b8064f5af11862d21f51610b6243fd46181ba65a486223eff7c5f4bd5a51f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h131e82c5f2f3d1ddc2c7acc5bc986687e99a5eafa799a06b8a7e6aed5d1e64f2d5abc5ef715bfca30b964ba30813245954d8505aad962695cda7dd4c325f8ae6c1f48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h390841dea4a5a92fdbaa15fccd2df8021411b96ac90b45a82373f2aa4300d2a60b7d823bb15831609b2403d920e58ee12bb6c9d9ce260142251def4228b0dd51680e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc166fe25b2cb20594a92242d04b9cdfd9c625f05cb9ea46ba9fc02702f6f14945031a25cf9741d64b542d29707c4576611c7cf94178b1f137d858bfb1c724fe6bfb0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af365fdcace34eed7ec3ed5ea3a47cd4a45a4ec41f0df38ea642a9c4f6810b7549ef56657f857c71f3b0ec5324806e0a2c9078fdbb412e01ca381cc5df75884b4940;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6cc8e486d1323b0b60394ab0a16a87ab05fd12b06ad4163b067cd6b89086d4e9a816d725e727469a023fe1e68852bc0f782f5fff80826b5c4c840e342a880c72cd5b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f8c0cb24efd13ed841aafc9d6614498ae32e57232e7bf5eef1d6ba683ccf265901347fb019106056f3e872197543a8966d1c0070710f8ece4f4b4c5290ca7414b73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h174179ec67af7327e0edab5e47774ca7cb90f1df0dc3be13dead519477457d57ae5482ce385de809eaba3a8baeafd521ae47df6cd68f5b140546c6c004e785d583123;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1198273fd1b878598941d3b50172979fe2f3fc7ab7e187caa8e03ee5e4050be3a10dfbe2a163926e4816c97466146b413c78d48382aac5b9487467860891c775c569c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa434bd24fea5eab83aa6cb93cefa32ef95f1ff0e052eb4508e2d12d0e702f4f5e1f6ce064f679af2a67783ecfad892f669a475c8b4d636bbc96517daeae043ebfc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1752456440e1fbcd3dea5067e06e782e531c2e1e219b61cc7b5ff6ff153dfd65500c46b0d4f68ebbb7a0504772065d4b55197a8bd6282aa3bcf758bf00a4fb18bf0df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h88f7d7dcc03cf7e4637a83257ed308702b2f7fc06da7ec68121094a0d374b4295e5af4c9e540fe2463a6d257c7a1d030688ca1815540d90f8b46d5b721fd4371b105;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c5077fd53c60c38e051728242fe713087850f31469e97b6463c2832fd626a98394fd2240d86bbe0df23cf54f7c1abb5afa3942504f0459612299eabd80bc19ce744;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca3cb3c1508b4d0e41ec457561644638e799094ac3167b333a1d6520b3ad2b3ea55dc0524f398cc27ab4c38a97e8014e28da8e5927aa8f4ce83081dd26aebab8aed2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha662cb655f705c726dba9bc68688767d8d7c2b8848aa7c113b68375a10099025d9590b776a25792e4c2e631d885bab6616581507690749d910bb0a2c2ebeefb0f983;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c32c38244100a42ba5be958bf0d1d67e30ca27b4a8ff89a7a84377459f0d0650218f448de605b8b4b4cca75b07a1dfc271c891b3bfc6049c5cc82c1ec9039ebf45c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9e08c09cbf68d06a06eadd5518d7e0e578f3acf91965e1923957a96c670de7d1091fb9948a84f23482ed4b99a7cade5f802677efcd21869f5ec672337cd9c400818b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcfdc8ab161c20fe1748d5cb4f4fe6771b3bd332fbad00ad3ce73359d6c11f62ab035ac9234e9b22f190922e7245e12d6efa9150619e2b4881dc18f6f4af473c07960;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7fa389cad5c91718e92d888d0951a6fc7fcaa1dba0b47b00674344e33722900bc13e43341479d06e03fd19706d516e0db6db4f443f88dc3733b60388889e212e1dfd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b787e9176b768a51764670ccf1c3139109243b15c354c398f6b7e9bd990c9f2440d7c806b0bade0051d09fe1065fcac142f6a051ba2e0b6cb10399d4f06e6884e2cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c0d197b189ac44e0badf263c9604852b24669629d47332227ad1f89f8552dc9d1a3cb9a8dc3390bb66b9999cb76145ed61ce7b7aed74d7df8cbea2cb72cc365bd43d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffaef0a46c33a3db035a188e7c650b65f337ab8db7b9d0c5986d9c6d194370e5048a7369beebdd8f66765f8475bfee6f0199d2902f06e37ca969b6bcd0f7e0dc3a15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1846d40d98c62e8db57c1974504c61ef6151be368929f417f335180b6fb3fed9785ff1c1f5e0093d99d5e7f48faec114e1b45e0118dc57cb9d9b584c0d1f4765525d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e3b3058bfc8b445722431623ec6a7b9d8f753bac7af44a370b9414a208523f0f404a289ed96440c396828d8242e0f70a47b0023c8ce224bc8afc05c6da3c2e05028;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had554a7c726aef8d25ad0237582556d8ca593d2052e6d59ffe99dd08f4703e940aece2a6c61f78edcaa393db1737eab0388ad4c4b5f930064c9b3e98dc83bca6f6c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h357f4769cd0b3652c94196ac06de7b4a8ed2426dfa49c60a8d48d00bceeef18ec8c25431794f8e1235e73f45b3900a0f16e1879d856d2b141dd237d6b58285f51c05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e87fec166a12a150c6458bc7ba4662305f7492dee7b886a19f1f605ebabbff16c7b2f5904ac91ffaf1a1d78537bedca384e16cfb9dbbb69adff57fe5b04e0c3e9ae5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf18b30f152a116fc2758fc6c300d7dd7ac42f519b7ebb6fa85da8fcf8762a0d0d80a8633ac4e37b7f163e09cdbc27c929ca637f4310c7015e7d746eec8747b607fc0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a8fbcf18ccc5dce2737a8c3bfa21e5c4d2501e1f878afc502c87b513752e3927d3f403cbef8349b53910436fa64ca6090e3b8122ba379bb3ce4cba65acd90f404fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfab2500b5d57025f8a835b13ae84d6b32ee42fa092f9dbfa781b52efa631b187ac52cdc5b2a71346ea906242050c5c37c17b55a5686bb50e5669a5f0a52245893b47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef78e5f17e02342f6385db125a8628c4a9637e8a8fddbb65c5a29c46ee5a38d230fadff1bfb7d6875662bd3feaa88944a126369d3d1379b956fb1068e632ef6f0a94;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h49ce0b1e0db4d7526d9618f94e4728e049b038d8ee9a7bb52be69d157d5ba651ff196e89cfa98b141a454f7158a41bc3aa8a38d35fd813927ad560d08b464fc0679a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf2b9e5d596503c586d4530aca60bb170d72d9e52556728f8acc617513cce8341ea101cf615d411a7b7233f603a56e9c74d0211a216fc5691ebdc289e931784af1add;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdabfecaaf96ebb2b7d93bbc3176f232f527b7136cda987b9bd4c8913f1b8878b06428e51b7c1dec7b00b8ad97c5a10d699897a0fb2f9de0f3b6926549da5a3fa7ad9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h891ea3e8ba9d67296471ba292ffd53ad5ea2aed67d68abf0fce127c6b9131e1bd0ad47a29c5720240106a7585d94110fa26994b6fc9d4e205836e28ee80ab4e325ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1be38df94e3bc246199e0871cec03436ca093cc78b886d8a0b1951fabec59a45dfa253d90bdbef92da69f2587c1668e75903a3b0aba7b64290c79c714d4c2f32bc03e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f18b41ecb00c5493f22e67a7a3dfc8967ed7036d2a772c781b875751aaaa6d5041719a7eec872f36ce0fc343f0c690b985a17654f735fb0591c9e7d12f8c3bdd52;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90078938e1a0f37260cac9fadab644407de175bc6e37433adf28cbd8d28de36f41dc51c85d70676ed8e71902c2c9c61dcc15aeb23ac1f51d2541a7cd31c7227d52ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14eb0bc028b81a5dd35c394d545fe2b848b08c5fd7718b91e432f76c994724c726fd8cc346070f41ed26a41f914d9150d957a2ba68de1de28398f174652caf24daec0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66d007615f3f2ff9b6f14a35a47176dea2e2b902606159f4ba873dac31721158d3b18a95427fb55497d47635448a935b5ad91bcf153514182bc0edc6ff85e5e2048f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h530a08cd26daad8f2db2ef18444257bb1ba9dedbebf998aeda1640417f83a7bbd7a6f3e32cb47da9c34dba573977470986eb69139bbf953cdff56d619c52b3bf1baf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d1cf277eb232e2a8679eda8f3c12229f4e5c0b6f5bd22d2f219597e48a6ba659e6c9fda9ee87e5c131f2846cde5a5371340db8be66353e7d556ea01537d7af2c8ca6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17af214b679958c0020f09455af46eedf9138bdc6ee1146df6bb8b87071c505faf795b0763cfbd55a3194db49de7ed963ef3faa41941ada5570c46247f1ad795f7458;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1db5c48adfd4baa88c3b07741b800dd7dd479285dc45e599e3926a82807de58c20d6fa957d8e9b03f1ea3d00f8f7f0deaa34adea389e3680094b1db6b7b80277dc184;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h156b1858a9277c3f4c10d6adf9c2cac1658184e5b2e63dc26811a33156d060fe18d5fce4f44e7c2e50d2ad9e4d82e5026f4f58ac33a2bebc1b67e03fb6811466421c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1093ead6631cbd0b3128d1955bb1ab98509258313fb54b288557afafdd1c5ffcc3d41b0a4dc0773fbbbdffc644c93806c779c9bf1fc5742f57d7678bbd2abadb170cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcf9f101019c9c2d2282934cc48b65d5d020337742ad6cba4747c0e27d6a4c8b32ba5d145fadb5f86930349ac23508dbf30ba1f05b98f6fbf0dc5881d2b33ad1abaa0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbc7fb4052f6f095bb70dea514e5438763a6189dbe17e00308fefe45736f760a307e65c2c28d7ce1cc8598220c0a3bf453b20822b845e50d31b42da3164a8db82d02a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e21aa1a81f82e2954db1808622e727ee17c45cb08d92994f9c6f841f4beaae807755ea8ed518a52661a4fe05d773c878f3a63ca902c9c41fadeaf033b4ab44e5f40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10924adda0375193ffdfe774ddb887d856d91cacca142ed228a77e748d5a9f6c371c7ecc2955a9db2dc52ed3452a8798ed2606a0fa84e8a31c79211a2322712775f3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dfc11c7e2c4b71cdb84ebcd3997de593d6920db77f42ddc55f8108e04f1a732478cefaf964ff7a541c2ee50d44253a0e7b6d2355f6793f60b2bec5c9d24b692848ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19bd93672c302f508c3990e3525d2273578852cfa1a7489f6228e737b89a8fd8c38cd41b57981c33b785639575bd301b0cc43abb6dc3620f70bb806feb007fdbcc74a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c65466a0901a484a5714c2be1c83316a06c5353d5a99e7ded2efc694d063d35ef902ec1bd11a0ff66f945e66bbd83953174475d58717b3cb4909e5ffa229d235619b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha662556c859e3bfbf6cebee14fb15d984575337335fca8b16bd3e03fe639b837e1cad0202d757e2106897837cb513d981fe504c03fc81705bbc610fe786b8e6734c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf4978958c1bd74c186a3066539a8ba7c304b8100be6626bdeb659a60603ed09f0cee3be253902d936a3723dbd82e0eedc3d6ea7bf3123501b858bb01b490f167f8c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab51877745d7018517f3e690964a0a6ff5797d2e9039a6857e7facc9cdc0147f0bd4405471d5dc898069bbe748fba382b5206a5e174573c500c37bd223d34145c6c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15f0a213b2e26902ae646d32028fab14489ae26b611bb890d4c6c392f367cba3cff99a0518fd439a7a611ea23f4de8f2008aa31446ad42afb55ba070ecbdee7c3d266;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac6bc93c656b7dd0b1582d0dd5294a4884a2749d92c81746118b1f26e752e56eb9e0f84b03aceb6d029793e51c60445273ab87b07d9746c301d307ebbb2d59a842c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6bcc3303c9d345d0f82d4320d818baed1bdc5a019154e90ed5b63b1d40b29ee071739a9c68c4ea201bfefcbe93b502c7d1ee243ad4a36586e7360578ad0f2c8ed1f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1741c99a436847a260775c7f3aec741e2d7107adc83087a1c0b2f971a738e579906b414a3c6a88f67fba1f588260824a9bc2f41f10408e399d20933e6b82c6199b2bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1949307909c97f80150aee4cbcc0549ad467354d4b272c3cc809812c69774c4f34df1b64c6f7eaa6c030439e143d144f1be21a4bb50047cf0c2cbc3caf31ced094cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7fa3e6086e9ae1eaefff3d32bc3872f71ab2689679460d99eca20e862a7f673c0ad3232fd839aec1ca2597d8c4004cd56117cda2f6ce21527771667f38424040120;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c17051d05918cb01ee494b2a50bfec23f34df4cac8f8784a5b43c679b8793564badd76e33fca3c4d69e0ed1b1d422958ac9ff4408dcb339d016e814d76753001e182;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a70309f60c24a07cf79c333f9f14b5257ce0b1beb6834124b00dccb2b613ccc69b37bb79f8904046b9a2fa924542606f966dda011a0ddc66bd5fc9fdc82c6a21fad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d13fe64e7d2acd67ee130474541e3e084520c1f8b87dc11b79d539228c13f18954036ba7612afffa11cee07a914a3419a771d9d257c0b923cc37c97f90db51020c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a80b6b1743151b3955d23cad607328006f21b5fa22e9f9c5899513640150c6bc4aa5da4cff6aa459f2d185eba5dfb350b4f6e6f2bef459641803f004414f19d05974;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb859573a4823621c7f690c5c8f247d7c839ab8a8466ec386fc6163c28b7dbcbfe7b8f804b0905899376b907d6a594fd7471cdbdb5289b43da181a221c571d82d7a5f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcae5d8d1d493701957f36614c0dbcbe7704f406567949d0409af762e283169fab15eaf380a7e77be72ac53c8a55f4bdb497ff475b518a64762269880e4ff557db8ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18eebe2df94401870d171603bbe68f1d58141b6b0975d961eaf4f4d137c73d725aef0d4baf347e15661bd225e4facd04287f7d32420371ba1fb2459bf80e6ad591942;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f357e2dc57860f5536a87a26bf146b82078bd50f92524f4e97ebdd2260d2e9ecc996e0e9a14ea2d359bb404a958d2ddb07101125a9cf59bc8edfb6397a40602819c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d96f7430727bbb659c28b822782d0eeccdf2dd23dee531eb1de363c0b451614e2c37a9d8dd1381c4bb9e93f173f13ddbe807875754b6ae06f2af03e710d0b9b38046;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e763441d9a356f8db444b290461aa7e8460ee3b2e40ae270a1158c54b3c314e1ddad2dfb828878a9f5535ba6235b7447d6d0e5d66d6e94d88a9bdc22b76c3fcb1479;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed17a637001da5eea8dc6e08358eea52049c020c9f0321699d4f0a82a55268f5b311e1a057e77671ef4c6e2256b9ea2837b919cf705fdc9cb80115ef9f6b4fef4ce3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11adc74b96bfb1e6f4e9244e72230be4e199a42f767a311bf0bc5513e9caf93494942292370a1dfd2aacea6c600a092f985824a71640f42a0a7e44d45c60663466706;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10d69a68953f9a121f222c3bd0e8f9cabceccff9052b40417f3e98ececcf8a799d54e366837b31e5d91b59baa0e3edf949eb52c2b65a17a28d3f5157345951a9569fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h45704e4acde3fedd1a2f3907f54e8dafdaca4a679b2c6db14aaea3f2c26bc6842400efe3dbdbdaea095a9384389b3aca98bb235b1bb542b0054b5331ae1f981dc365;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d0923457967b35652b3acc3c26783383656acc776a32e0e5fdfeda8fe50fef664e264095577be53a6561a24b34a66e66f7640538b731a14c2609578270d27144c1b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1caa6ad04514ae17b894eefc4ed626726a3aa10d5a29643bd8e9cbdd140c75d447962b09a527d2f78fcedde5f21af6349c7f27a238769292accf43515de9eb549839c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3b7d2ec707f83bf350d1523ad98dad170291cec14a84b67d33e36c9c57c14f76bcee60b99a6256ee9e21393c9ffce368d02a6bfc2cd6ebeb02c5ef9b8868f12df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb171aab208086ef33cd6fc9ca23fcef6e2b44c7c609e6dbe811f24a3035419902d86972eae9fe46401d63c08211d9905ccd8a73edb3b9d60aba6126641b2f68c71fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h72ff7e9abc00a23e26c75248b2b73c6c9a647f0e2ea933873972898a2f99462c8e85e0d70f71b8b81f87bdba937d9605820e8f4ac4ce56a4820352ca00d936cba9c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h43840e97bd1d807f946b625791059c4c6467f6de38f638ed8a7f0363bd13e649a0dc280db1c9a3d858eb0fd849afc1315a6299090306882b650aef7a6d44c270da83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9b2d5bc6833af4debbb9749c7e3760dfa694ad842adc915d596d85b912255f7c4a50e9e664952247718037991f876b7fa88e9be00efa6e35c810dd0063ea58b0ee4f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1198c39f1d80a536b01a10c8f72aec5c99649c9f0498a3892f4e151779200828139e7eac59d9d24073847dd8a2592c4c4a1ffbfb437c104bf84869430e38349ad33ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd5a751336662d02a39e076e6c2ddab67bf071a565d1bdb0df4b70e40c7482ecb9efc7a0129b767410cfa0b959850d535c365137057c82e3590cc4710848d74ab14c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd450d5d7f06d0bdd8b2570566c1bda475473967b02ce076a89c29b53a4d40883a1beb4d2b7cd586d4f089b3e8e3b4fff5c632762a40cf5f4d08f11ebe98bfa23568;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9de85391797f42a2a176cb03edaf999fc67fb6733a34a929b0f1674071c44b634414288a013d048e1c616590b68f875600e8c4d9344de31f2f27bacb725fc3f8ba87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcb4dff9c234ef34a5852668fdf694a78c2d9bb46246929e5e247a58c9bdf4bf6749316dd35036ccd13b22628afd75e0adc5e5f3179e3eafb12f21526c8008148a4ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h347f4bc796337a0b667212b4fe39416ec87101b72af09555f2c80aa1cb6047a9f2b68e17871d1546648441b71202ec61d96b9788daaade6beb812e667bdbd04053c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf7878623fbe75f3237d6a3bcc3a161d0c217955cec011c6ba11e5f2f81201a36100abad40c0c306d4da92cc4167d8bae831029e9c05308bbd3141f7dd180fbc9b5d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd86443078ed52f162afac69bcc042feae2efa2d20d42432c807888958afbe4d1a16e031a20ce5eebc480744d60ae2211f2ea27dfdaadc09b3fe5d0b362d3bdffeb3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aefb35020f0d378a3c71d838e64bdcdfe37de5f97d19eb1244ba2fcc3b6e6e91a3f85e8576594afd72c74497e692e677d03605a68573947633cc4a309330847e74a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103d7da639589dfb44609522803c9a35d8c8f44052d8d897e6c5b706432e1bd31ef0a3d9200527141c9e566e17d53518cf170da84884005242ed7fa35cbe194fdc93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a78317680434f8a74790c0ee1df2827981828d54395db01796d1fce4822dea6e409e963d686d6c6b055c2553729b882b2e5b36c3a738d8e346514173fdc7c0d02681;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2a30fc2e11ac1621fc6de13cc087023fe73a614165783b78e16ad48f5838a0cb706138cc5b0f89e62df03af260e62ed00db84d14fc450f369f2795bd203664c21cec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa8a7e45b0630f781d5e5b6651e14b56814e1b30075d57734df2cf5618b8cc4d7e6a4c33b3a5a0c13fe20e417b467efaf2e9d894e9ab5569889506b49c7a4d528766;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h142e9d800135332d42441b845b2dd0cc4c98ef3d23560f11657b47d76ecb43301e5e9265964ce10f5de9f478f9adbc73cdb44b523fbba96562bb1f7929dba5e90430;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dc9b02737814667c4b7c2181c442a8e428ae28c17531a5e16dc12029dfe6783586f6875c4d48c8a8dcf9ca2e80892db2f02a32f647b0986c3ee195fde849613bb024;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9a7758a43aa96c881045c4123a64e15dce3a505edf414a2afa70915d6b231454d87f32e609969dc1559aa7deb0899ca753f3360e865f229b9912d3d4b3ff3bc7bf1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a0969baafd4adc0a27227d2c8a3669e2d78ff54c17ad919878c34d96437ea5032392dc75508c5ad6c1192f00b8a04d6eca5f2b007c8d3d3ce5f1b517da64b740125;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ad5086aa0d11fe008470ca8a98e274f9b51fde4b2f3aba7705b30b5163ee10d12461703ed6b4bcf4e9a065f2cb32e145daf760fab35fa9a4d570ca602e82346e8d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcefdbf29545e7c9a86446675a0c9b2331e03c1c2a30b9eed5d23b27c901de801e6e29d2566c0919db50175d4af9c9a1dab07d95d39d1939863fbd25b479a5716f0ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3334b43d52a1e54b4ece5092558417387422e27630e6d32e94954033c2a46dccfd095d0c6197e640970aed859d95e231f325d85486aa87fcb96cbcae76a9c14eda8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c0d668a4922676a022abd62483cf3630a18c9a0085fc73e92bf4a340264d3d04b1de758fcae078718c0bf8ffff8acd4028cd4cd1b5b06de4512fb7877df2b48dd05e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16dd1a7c00e20993c6dd3b704ebf1ecea8146c64daed1fa2e58905d2a541fdc324e191e32548873efe77f16ff7401a1a68aa6954652b864dd5d51addfebecee417120;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67ea336bc00f035d80430780f885f8cfa8000677a3e1db085ee8c5002a9adc57d5fc4a2a62449b12252e47b5ff714f5ff6167ba6dc1a0bd3f78a41bc06a6ad9660ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h448df030055b9ae25c767ffe33b79d843b41d6a835e408fe7782bf8f01b2397ac16292b4bd968085ace36d9759794420837ec19e851f58ce4c0edf37890968e229c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba426f8336678dfadea080c31ccec521c5a1042917b7c1e734ec376972b78ff83ccd31bbaf4e9b995572a30e8805dc996df779b4f114124505fcb22cec0ae50c771e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14e56195c266487ef90519ff5f5e74b5e41a3451e6db822d18c63d7441444cd2a7bb2fc2644c83bb7d2b2cadd8b1b4aa969843146d8ea604612fd00727bc681fd1069;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ece802e9d7506464c9f14447e63ea5bb88efd81b5c4bfcfcf043e47c5cf4199767d44bb615800a13bb63440d1985a6d86bea6af8adde22b23a9f36192639c38ce5df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f356471a610b518e7789145a29a771ff8ccc5fe131edfca99c76d07e0a4018666c5472023baa23cc2cce3a2fe84fa8b0bc3d602bdf094c6e4d1190ea1f2729482bb4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfd3e28dc66786829e4c595bc5c5cc624f633343e40daa7fc1a22b0fa052887a73f4a5d9f104e36a0a0614031f171f9d637a4b3c26ed672f2cf58b47b12b07aa8324f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a5b8de984b59868827ef72287673588f61ff567949ac53d9df880135b0e2eef610cb8d4879106671118e93df5d7fea6cd75efdc1924ff9cf71c2147aa64c74680ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e5e07b8af9e97c5b6bab5b65c234189688b47255bfc908833ec2c195b5179e7184dd195068af4e22124234f01a9eaa2018be00170d3ca78d79c8d36accb1f8adceb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h179004f97bbc7efdfc60deffaee2b83cc70c27ed2c89c68d832f0f67ad3657f5e0ba7036f1132a78949f2bc3686312ca721b64c06c439b37b3b2146c41460cb3f0412;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf35b8b4e55c8ec27a89ddbfcd8f26cd5ded8493095f9eceb1d471a2c60d316032d1be059f33627fd2d90e821e1bfb23ea92bed403345a842f7bff6c7b6d1b902add6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h123f3b4df090446d66cee63417a2eda63d42e67e8c21889df85b1ab7288353bc6900e780d195e8d60359e73cf7119cb82a6dfd377f44156075049c17ccc582a71213b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h745cb98a7e5cb91b3bb198e49e0c43fd229534b0af4fc298dbd56d66e569543e0b83e9c402a5d896686a6ac236427c091286f94a0dc58525e256e8402172f7bb71c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfbb013f4d780002fbbb8dba5e0f7c8de0957e2275846fae9b601b118c1621cb1a8f741cc9212a0ac3dcbfbbacb9f4a7bb75e0607b859716ecb66bd426caa3a9693a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f40191965595fd9d8b93fb684af77f2a0e3bc9bab51c28373cb8c0f74e617cfe92ca7f02c4d366651d8a33c17421886de22e05bef0cea7d0bb42f77a43ba5c005c0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc42b0661bd138c2bd8468de77f48e899cb9e26bbb3cad79b4fd8d9b30bdb7aa5a989051214aae4a0e3492cd0685184d1ccb563f61189367ba1c6dbf21ea675931ea6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h122fb3dc962ccb9ede855bd2c7f1bd214ba421e452b7094efee731797ae22a9f2cb7f303296e13e28db2cb46f85bd6eaac1491391a109c42986b3d67288d49470abab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1219d0d29d4d56576630c3cdf8d759f073b340146b061d1a4189cb7843160d84ed29d0d0716332e1c127ed1b2f3e276fc4826b36b1fe763d861c8c1170689ae32a384;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15df3f128f124a31b1f245a9e62f6587a26ae9abb2bd99638f19895ea7f638bebd6b7ae434cae1c9d67c804f84d131bcf585003f122511794255d7b290a383c0e16ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc68c37b9136b4af3baf161e19bd199484e7c1d10bddf779e8d6fd9fbe6a1c3722c0bf1da3ebc7ffa04ef5114f94d1986bdd369d8f741439b22f1109ff69ea7a092a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6b6d9521ce661a2f76e749af3ade4c8e4a40a7980d411a1a255b297e95e1530bef8d82b8dfd53c906a0feeac03da663c2b3bf321bb41d1f96087bbe13036cad11385;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf28b69fdf01815b769d0c0a007de7df850385ca6f93dad3ea0fd8f1dc3557889b4e280d0b4b61d5908d10728dc236830f662e0e1b27674143acb9012c7273a4ba99c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12eed52c42ff555cf6666bf340eba212d486bbe3579537115b2019ab5f85308583566c2f763a887d61e7e64d9c0ce8af509c091595b039e13cabcc57c78e88fad14c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h158d1dbb8ac2328bed84ddd4fc744185208d0b25469298484c39a33d3d2c498dfb1c4b7fc011d5c44ca2a1a95e14194dc72b0671e193b4e1805cf39b785c92ca05c85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1359bb23454e498fda0307c16a5e2b857db5dc48874f96b160301768dd0fbba89acf108acbeeb0ef2462717ed068918b53c8c1ed1c56add81dd0392b5c3632ec9c741;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d42b9d7b523e8a4f9449a22305229446a31b9a2ba87f3795a2209cf9bff4c6dd7aaf5b0f6e8328579242b92ecca0146c3e8a26ffa150606b1fea918876a42538c1c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9a8b62a9ed9e088079d14740e0cf49f257737d7cefecc06643af60095f7f94a6ec580ca487d503250655f8f6393240036fdfecdea227519fb0662690fcd833b05ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b59647ed898de274733e255b5678f420ada02da11edfc49c8d4a49126c00ef7cad6f00e320b9c970ede852a170cffc32f89054d9a11337eb53750b0d42a31889634;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89153104b73f72203e3c0b598578c7695c6395034ef37f344359e7f35098de5555cc68310799dfdad20e6530b73b90e4958bb52acb3dea0a44c9ce1643e32e691126;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34dea1ee72e8c0e3ccf0a73592cad1249649b7f599670e9c35937dca52ec461dd8924e376cb11eba844e2bfb58c9e1d1e8e349b238560ad7bc4e3cd1921725dc11d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7aff4cf89d6829ffc0d5070f4224cd872ff472311f0f50693089736d4aa8acab5a2e80ff7390880904fbc94f5b0cb684436814c896293787eb38eb312e9fd35de59d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1447136924ab3d4c27223bdfbae68515a353705c2dad96e1362b5ceace1f9c0c81d950f27d834d561b8e10784c0ead98894c1347d2f01929a570995e55bc46bf89fcd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h115df6a0ea28a7b60f96bb97f75d7f8ba5df62c820596e350412d81f3b5cc7f036bd88b7844ce842aed078c4dfdc759fe82602cfaf11014c74dbd54b4f3720c501be1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10985c04887c99f3e1fc4ba96a8ffd5ce10c26b466738ec42180dc9a01b891f99aebb98a1583bd5196a27efb5056799ec920ee2bf5272bf7eb4904f474c22e7e454a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ce45ae559b1d6eb88ffa8c8d8f3cb49ca8d4ee3d3f81f0c3c75a7afc6b7f53cf51984b640b5b5a3869baaab2017081de02baedaf329f16181fb6460d7ecdf9b46c44;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f8acd92e6dcdb61b1192756b119d396747675613b7d7a95eb5bbcaa498ea7d5ba8c0300b1853cfd7b8c68e5036010dd9677951386564999956b5463452b826a725c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h360d10665864599595fb28735a352f1e34782a373a2188bb97066d73c71549afa31f9196d9d107d920cc8c68aa2581f2177089eda3391bbda68571a6ad3214360bcd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbba199b981dba67d623bfd9cf072b155c05c007b66eacb896dbb5e49aea85713120c9654d6fcdc8d4360324b54e7c5965e9cc725665f0925ca7f9a5ca20dc1758af1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he8b1154470818463d5b5cff6dfea103f8a1017a1aac9fcd47232ade249ccad6ffe74d84cafc345bbbec175a0779aac259b0cb1aa9665d34d4719efcd8b10952b40ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a079a5e91ec2037fbb4e91df422353a6dbd72b5c6b7fe743fcd007ec2405ba2d5a2d84429fc611d2cedc9bb6d7a200b534b7b36db28ad1c0db2628fadd2b8305fdab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1179210909e0e14cd3fd57fb9feda164b29ed91ee0f0c9578d75b0cc0da013c80d0c7df22c03c2726021f864615ae8660cc5694bf28a9d4027fad4f7a0bf5b5bfdf6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12cad03eb35b2c1c2cfde5068e59659b1d4c5873ab581746d0e1b25802dcb98f6175eea568bdbab8773817b7d6ed37b1f3c06fd6b7e1ba98938e414bd82702ab08475;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h128ba2d574a68b4861a8c7a47c36721759998a7da1acab7e6e116339d67db425f86c571f27606b0bf16b729685b9354fbaf0de98d61a7230a7b6853f57f38fb5eb145;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f3258efd7b965b8b92aedd0ba75ef1912389eb3f9e62c91357d3b745210c4270e885733bc4894582965b7dc01120a74865a0986033967caa2d9e6a4b9f3ca7155200;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf16751ec50d457c10d768a034d609c561c6edfb16c2d003efe1fbd6eda40ccbd1ce2f2af77a4dae22eae14d77872111eb5fad8a97d020fa4b4c8467ce6d1be4ef11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14edacd162b0c6f1970c3c962e35b811383f748e7c5ebab4b1482bd6fa8b0ac3baa0f80404437d6aa9ee3745fd215f10560c8b03ed922e4a0305f960fc15d3e6666bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16818c4824fbd18bc286bf8dc806ae0bd32116de97c933cc14d1b5bc62117737b5c681472541031ba1a1ce8ebc2541e8ee014ca92eb5ae0859b65f758ea11a235d4ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f9eae34a9741390bec04ecf372f3ac52fdc8523dee1f7bbe1b3de3eb89304b914779f760a96e098364415dafdbea617ce34fbf0c6fc1d96da7ceb3b475738a6fbb2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a27970a3fcf58ff29c09f811587aa27529afb378efcc6203c875aa141d5500ca3b32c0be08bb20b1f0474b29ee4a120e08afd5d576f5332c23473ad65491fc8f341;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb93fd11da08975c6f46860c0aba25baca3a13f0e5a1c31f4f7c6a769832b3c0787fe0347f09d4b71de1d43423dde614e01f83e70fc9f63c35b437a3f78c73022f32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14cda1f4c3ee1a4b18baad8f146e182344914b06ac0ce2f58d54f4996736daf54b66fa091a873ad5050f0cce6d62b1e7b359e36b1073c3d43c259b1b67170860deb4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h52f01d8872e4912388041d17844e15f1c5950b16a0ab5c8754ed7637c12928cc1869afee73665fdc2fd5386b5e2dbb55e08531e19bf63b89a1d6afd66f9564a9d82f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9739e670bb8e586c58511c9638fddcc137d8e2ff6f6ade7c02c5b86074de6f4b4eea4172ec8c509f6e30a7d2c4413c42a0b11cbf568d0934fcdb6f3daa5bc64bba09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he170d6eb748a30a90d42a45f5cd36db4a566fd2c85d0e482eda2fac4d7b6d6344cb0e61a43b6e3fd8c5b825e5540c17af586f98690e7acb00461488d32adab1da66b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2f8e09ea77efb2ea535f420f7576c0193c36d2819802e0edf691891180b3925e09869cac12156b6961df1b2ef03731f6a193fae3165125e399e99345f335c8e973b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b57005126f730f5a40f65c9ae92676306d89d9e31bf54d751684af51edc167d68d46bb51ff31f34cf86d3dfd6c959aeec534e1bae32f6f9c1bc7361e883ddba72a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e1b4a95651232f23b73e854f3566ce49f1078d04e02b785c3f3c1365c4759880eb13f74fbd32d17c9a218c314f022e98b9211567c7c2380d49277448d02d3aedcf06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38156d0b07cd0f9b86c60428f530c0765566b90a0d20e13466ed6d54681b863b3e1e39b2ff326b782373e15dfcd5e6308b769bcba4c76f88bddc0ae7d64ef4145f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdb4d5db6720f650c310df6cd9f9ba7e3b8ee805b8f68fb3c76a5264c9ef116d8587bb91b7dc71f8eaea9d710907af447ff51f8d9c5a03126d0c076fe2f1196446511;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13a1d314c8a3d3ed863a34b916e0d966768e92a7e1bd17ac3b723fa20a3a189c6f904e916f9bfb3df48ecfb0f436554bdeb558f10a63abb0929e50b80054e1d548a8f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha626172f5d4b27cddca437378ae68c803f3a3af84f504f149fd9810dc0cb4c8d6e7a18b34539f2c990892ebae1845a8deca222c505d1273cb1f1fb23b297c7cdd23b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7b7c129f8ab25fd1fd40b07aafda181b76579d3c24ab99564065cb92f13fc4c6222416a95dec51be9186eb089f9343b56b2bc54fcfc765c0eb155f9240bec4ec7e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a1a4bb659c87a200f0deaf70eb3c195ee1b6bd3783f89ccecef7bee113fd1d75d3ddaa65d34c36ff5832218fcf2cb20109dfb84e7d33a2483f4b28b05b2d8eaecab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1038672df489220e0f0bb300db7882318e7687b607cd91f412aa22ca428f54e39cf8f7e5216a3959028794ac17f4e943bd92aca3acb0dbfd8fd965fc883f7c2ed60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ec4f624bb87b9691cfb8c6a3dc725492aa116bd8190945cb6f1735d3b3974519792a72befcd913d1dd2daaf75fbb68950d531f3671c289b6bd684bd81fd5238e8e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h153292b989117dbcf74fada3e33d9dfe67b1235e8b386742c98c7511690a168db3e816dbe7546a29dd07be7e31fe3e94f36317828b006e51f049c95d5e174dfd899ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17fe34628bc9e2e28f337048b18222fb39ec93e3c52ed1b9a6142d2ce704bbc884defd7f3356bea30fa62dc4e5bf6171efd2bde3bc3e5fc37c5eb3e96151e41364f8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1858ab0a6d3311fad6faa54660cc744d5d58d6d597071e77810af41dfb08c92385f7a38abde7d83794d5575279cbee674eb090ec895163e4ccd0eecd4228abebdd261;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13a625b603bfdf8ca63cb9a1a70c57ed8ffd142dbd090e147174547f42ab8ed28599e1a9e1286a3a5ab4fddd4bc66b4caeed61e091b7f1f99b318432093f34878cb3b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd74305802fb118542de77321ffaac5b38dbcae2d56880d16331c6cb5a026de20dd8c6f913a1a5ecfb949ad86f3c82671eca54f972969319046e948372e61e13749ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f9ac1142af7dec9bc1bf03eedbcee25f2ce48d5b3499bca4f1dd1382cb7c015024a28cc61c60f4c1a1aaeaa6c640f3f54a6ce63e5395b1aef24758d6637c33c1fa3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dc8e29e689a0426c5152f8cafaefd58c838b22846acecfcf6ff4b7529eb77bebc5e9f7b5c9a0eccc81b2a1e938764cefd82749eddf21e811844bdb1603203d8442f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ac223d1dff1b76a1781815cfa13a6c7250ad3a1afc9bbdf7e16ba7816b2af099eef6bd3ee5b54dd485c4d02d0b432331f2eb044ffda8a5f2843f832257747fa0cde;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h182c59cfddf4f6fe61a307ba4b6ca03c3437d6ec56c68050b126474520d7367f49f616c1cfa1dbd728afab3b3cd5a12251209a3b4421db2b23d0edbfcda0cc2bb1f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcfdeada1d0edb25bf1575185fcf1a378eaf1590c9b20df9de69622c9ec74578130bc73dc3c254ab0965c24eb430de3a59fc39aa88f8b717552d5649adcdeb576b67;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h126fba402d6dd962d3be8448a08bff764f96774d555cff880d21fb1b22a07d8da38694481f17ca0d0a5eb9de8b253b1e19883b9fed7063720a374b97d61bfcbfb8a7a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e914edaebcef0c0770011bc3eaa65a5aaf4a4dbd016fb45a8b5452d5686481ada4411a1ecc6209ff27f596957b3da422701801aba0ad4dc3c50007421a4aa3e0ab9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f5319a38e8ce4d6e0ec1b4d415f8c472e62b1dfe61282df7571287576db1bdf51f2901a006785d6c9135d9899d5f4d8ba7b001ea110e94829d5cc65fad816802438;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16be2304527f647248e1e4dc00b7490d06a9ad410c5da6bc5abec1843f8473f9520acd18f8ba27108346175a37bdbee347baaec9c7579a4f6a07201e1a2f67fc36659;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h472ff6d2ffc3b20f21e97c7091ceb20bc0225f3782c04d96da1f439dff59190b6aa4d1c73af552d50a858bde3c08d76a20542021a272868162af07e2f33c68581a27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5cf7cf5e3caf51a9bf375338c4ec5f4b0f34c4eefa3cf072b85eacfacda61472f3534c7db113a877e342be56b90330a8e4951ead0950447c1a5c81aeec9728a5fc76;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h156c0eb1b341a66a7884eb404674b811b6306a49dd8abc0ba893b83fa2992dbeb88118d24e86b08faa934f463048f3ec6c030bf8affdaca8cb4fd2eaced84a535d938;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h36c100d6db1eb3b2fc03e0ef5cb1d3be4adf080e16ce0d049794abac66ad61943a37937003c013986638ad4761034333dc8519410ee7382fd31677621b4eb3923adf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe527d4c733c490cb6ca090f334abde5a0477647f83eeba4dc6eac671854c04c7f86cba2d108d7f373416daba248ba304716623403e395caf603772fc8f6ed585c38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105237cfd7a866c7c20cf3e3883e29c9d6fd8cead177d3f47c03a2c7ace58a45f99619f77074b1d9cbbe89600114085d453049308d29f4688e61d4e696852cc03c93f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heafc3b9789f694b70992a7515420fa76213fc01fe65a0c83c02e6f80957772f917fe49c3b889aa0db3f8eeda6f90eb14297a3db8ca6220b1e40245e4df24aef5f1bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haf748a60ed06ccefe9e3dee0fa647c86828c50647de5ef5c199fd30fbcadc7497489bed6ea23617b9704b9ba864e0c52669d568befcc350ba016a781b9bf263edc49;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17574a99e06a2e668b8ccddb12059bb48014274e944b34057c40c47690b60929b2bb04e656833423c65a3fce4b6eafee448592b4da9949036b2491d998634df8191dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he63ec510c1783b285f372d174c68e664e235817edf433675cd149654c394be7df501978908da458b7410667ffc1e57a5e7ed2bd0ede97d94a03d0de8f85052118d4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c5b13afb724fb89b0c151fea2c475644c265cb468e8a5a7e02fe229c0368b9ff10d8788b61b0796a5bce89c98d5ff782deafced42b1525a17b4d25abcfabc6f561cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h715cc49f490edcda4236b783908823bd03f0c994f7ff11d948d5ca05ac16a01fc45ea5672585b83769eb7d6fd6ff90c0074f8613f721fd5590fa652fe95e3384244d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he89a4ffe5fe59d898e35f3fc332efec0406e809cb2da40ed79f0addf3fbee5eb3e606a76ab995534db8db741731a71cef5a45824136f172f9f3b341e0ab5d6af37c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h39688d9b236ae0e1783862d48eeec69d1266575ad0e33ed1a8e12dedc50fd9bb4f246a3205d33e6d6f3b8a6bb92b34e88c7d956caac06979703292983724245b7424;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h369c8a83091fa9f0239eebacebbde98884cb142b6cb364504acdb946dbfa48164514ce744a861f3eaefd28c047c93eeb6920eb06f3da8cdc07472b997c7477c0ff38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h85155194042ece8984a46faf405db102e744cd3e627167e62646e61c05151c86787de17a8d6872925a14f9c2e238dddf9c203979bb2f94a6c4a93bd0f6b6bd18c585;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5fed487bbf2ca7f419db491ecc35735a77487b01233189a3bef7dfa3371a3c839966c61227655792af055e3f47e43176ef38d9fb29d2fedd744065426019631cd65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd75058eb75f9b9c78ca7ee6ee7b755a535219ea93667cf3598fe1cc629267330d5fdce45ddc08ce10f9d050d6127337eae7606c21e1dc22480fb9ad7d3a2fae80be2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h94f4453e239ea8e5a3bd2c33e45834bc2800a2d7931071c52edc5f129cf242d41e842f30abaa0815534a63db74c98f96fae1a6218c0b1355db3a51af19087fc8a66d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h170d6704aa2250b4e239b7f80ab5f9d723a5bc0d6c8c0def13b035790a1ae8de877d5da693faf40e4c6b81fbedf0914885538ac53c4766f28382a75d650a537d8a98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha03590003cf148e37a26c9a89b26c2476945603839d6f5a4c9d1755de0c7335624b244edc7ee17ea7ab4f161ca9f795e510c37b4a4341c88c862dbc322fc7b43e8a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d705e5b56986d9d8c1d341f5c720be86ce6a99378fb07662e3c7e2b1aab128e1d88d852decbd441865df834e5577c15dc378d249333b1f63334a511cde3bbc53fa7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d17bc13e8499f7390cfa426cd58411e0dd52223e4f484d9fafaccdd9a10d5a2788049f3bd85f9174003b38d919d97872296ec4e89b563bc2f5c4006ee176e34e2dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d7a511d581d90e4c7d02443fffc5328ea40f9447298b8cd94d8448cd7dcd851bfdb3ef4f6d6456c008592ba641b42173fdb0f5258efabeac7fe64d895d2062b23afe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1badee73ec95a3246fa13bd76f61dd8d8f95f56b8003c3e6f09c2923983e95f31177c6a5200a623a831553023d6deef245aef8e87d2095a6cfef84a6998309233274b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h468dcf6f82243705257a6cc8e5f74b599d922a6718a79e0ba18455a5ec115907c2d25a56bd56af4f4c1c86697b5d3d4181e77746255827005a1f4362439ba5cdbba6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h178c3006e9779c1a3e41f052a4f9004d4be0251edfd8824a9e199c23cbe776a796ad03bc52e7cfcc8f977f42ff081ef02514203d09f5eafb4c0a8a63519ac42f16312;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c6559edbde90271f322bf550b6e3f5625c33f5bd9fe013989b3c3ddff93eccc8e19deae97cbbc9003a7ee14dd16ce37e5ce65d5775edfda7cbb5bc25880757dcad8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2173d6c76545ed78e956913636e6dd62e914595b35c967438020a1b1e1585c79cddc9ae9274babf678a3b1423561838411fcb233b30c88a32472b43c63a29065cc1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa897f3380feb518809a0569224add7b8bf7976794f4d94b8e7774fddb8272483226c1bf335346c13e0dc4fbbc5f1d15c1d9f136ee07245fd93bc7b6d3ff97258987;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb7cc88b675c88001901a5e9872153861340e9c2ab5e7e28d84e7b5981cd2c64d3052e93c45af993d9b7d5f4e9e483acc8d4ad2df8c4b438c61945367c48ef1395b34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7785b2d1bcdac5b1ee1fe88698163cdc75d860cf0ee4d7341a68dffc027ef7bb6afa4d9ebedb118b12023667f5bc225300f254a6a31ce3f3e6c5c9ffdccb1ab832d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5075e7a5eaa7973011513726882cb6ee01646290cf5b231f3182e6880cae864ae3f7fea374ca4dcff4952f00a6c48473241f4dabff16bef4c96a58c55a00363ed49d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e8a98c82a87ec3a28d09e65b42f81f80044591fc48880979ed718a67aa67027575b1425da390b960b978a89dcab0006b17e8a22298e29137712a171110ca9e9cb95d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a52692dbd3f0a1b1ad7d8b73d17e17d05dde66a8168fca94571a19fb20c4bc3ea36dbbbd6fc3f6cc847fad154e932e80f2cfe983fea03ad4cce78213032bcf2bdde;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h163fb3f1231b21910baf1714ea95806ccd07f9558b13829601ba9d524d36b3f693b1df33ab9cab9f702179ccdf8b4e41db111eb1173a7cb957e8759441798b8b887e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194e6e49f5c4547fa5a289821949c443a05e7aeb0bd7a54d24a6e9cb699a7b4807fecec646b675d65e7fd578c45892b0f88ac99f5aba10ac28f2c403569b43e1d8702;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8544a4aa6a67249a183569021b2adf2d8e125b61fd54fbbd8de73314f901cbc38ef96e57d94496dd90110f108afb69c7829c69ad75829a4972210f179402bfb14fc3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2d1e12e6a7753b8b0b1d0ae7e6a7fb030622d12e293d3487a2ce467f9226e0c0e95c4ef3f109d056765c15f63823b2fab4a48837f976d174426527d02d29acb78e8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ac0ed59dcf26e2c2538544bcec6f8d8b67f82d6c560f60f89a59dd0c0e90354e51b1e6151244cc023620c51b6812cc72f1eda720fc33e6201c125ff79fe4813b3753;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a0eb82febc80a83028484d1311f07a74b8cb37c7462f3547cfa7438fe9c5fd731d52f4fa4a4b34db624b1231a16aa863ab919e96111dd8c4548c3920cff354631f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc9e8ec30f094b683a1989cfdb58f28649aabfb1f908fa940b755ecc287861ff3af6225d5478b40d276dc2088fb283abce5b627110bd6935a24b2e5b1b4297c27c01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34111d87a774965fd6772bafa9bd1d34ab30cb530b792080ccd2bc0c0ffbf2f1ac69ebf5a1c5493439ec2197af0076fee14afe63f6d818115d860b2dd6260e91a0a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h124ed4969efce5678dfc9fabd6366b988a912616dc3d4c62029769250c2f4759b87fd295443df7477359eb561c2af9472b79840324c18ce7bf355be521bbabbf0f0a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfbd027379368e2b8fb5c82cd78dbeeb0a228230a09f44a58a55da1a494f1d3760c90a8925d962d3c6da7bd1764b3ad6c62ed0bec8cef9e990dd9b5e5c00744800167;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b3875937a21d6ec714ef81410efe32986d0a6a47e9f6a260482f1924f01ecaedeb0ab022bc284cb5ba4e6135caf0ee7a9b2ca6decd7438ece4db63146cbb23a1635;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1725abb127b39a96a817ea33e20725d4fac5d0ca3cf6cb028fbbd3e6241c6fe5ac9971321d6b435427a1eb53818c20ef70bff48ee5ce87ce57ccc0d901a3bf6b51bf3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he037686f7e9e0e2aaf486595918796a14b5058431bf70fd0476e13dcbb9f27c2a846c02077517aec991b9f22b66b0c2652f06aab4d59147d667f243f6c263db542a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9c9ea1d42c4dd12b859916ccecd5867df5c4dbad49b9fd3490f13acbbac2c254051922e949fdc166621eb273a7366c7debe5a395aa2dd2b16a6c208a03b1f096f10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha34d999e45084cd2502ef7e044159c701543bee0b5c88c210f8ec4b3252aea7ebeb91f66f2c78bd478643c78ec5bc7a20c8943ce37a81f64ef75065776d397146b14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9c989a7e4c93fe12ecac7b0ec42b20c1f1bac6e3f9dd43efedf5dce73be6b48b065de972831a1ed77af35796fdbdd3097adaf2c2b35d8991dcc59aff5704b131e7c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a7305b54f4cb51389e56b9d55f7563a7a27e8d017db013a5d9cc89b7212e05137f8efee1c05f41103e9aded88b19e3ac3358ef0c68ed8ba1ed216a1a182c6cb3d35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf05e0fcfa6d3368c8cbd3f651a37c58263159a36e76f68bcd574d294b0da84ce01da69e52c553430e5ee6532f8013099d2272bf1f40fe1f89ddc1b17d0e7abc4ee04;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139b1d7456b089983205a9a22e2d87bcf270a6e61ad2eed5c43d2efe080a177b88544180e9ccff4b14a62e152cae1d3a74b2d561d9d1959e1da56e12a58845e61d1e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf9a397c12637a83e2c2c156364c335d2a61d902c99463659384f775ef69326259fa07783d34701e7ca03a0e93d1cd62342cf78f586490d49034814acb4d7f42cb64e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143e686d1ff9fd043b5665ff87c976fc688cfa01c073671bd9a35ded7bc005629a5869866db718f544d19784701e2e3d314afe09f5064afa823dffb7e3886b0a3adc7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1999dca1bf3cb1ca6273d801123e982ebb8fc93b51cf23e750ef40982c0f693b0bd68b10aa0af3d524c8e6e5e5586270294cda7c1674a89132d30f835fde0d870a367;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89eccf70a10d4689fe9f0728af45027222e71c480a090a23b599792d061065b8e2e5f693826b50d1760576080b575dba9d001260b643cb2b1f2fbb709ba54f616502;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37774b3807f731e311998b81d93e966d4107de5f6a9308969d94a51fd9eef274526242005d83ec736c2b3b45c28aed73ac2a34d4e13297b20facc4dfc90df8990d1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12d0feffc6ab6afbd31fb8a2a67764c7261dddb349b1e4ddd9824686e0ed9857501dd7585e240d679e35f6b0e57cb430225cce092e3400063822754c29a6f5b6bea67;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h54cbdea4eb91000eb82a27f0f5b51e407eebbf82e5c2329bd82c5563c6413e771d73e6337637866858d973bd4edda390a2a729843137aa1204b17aa77fe7a096c33;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd662af1f737d042c06e90941856640667592832bee205b796349802e047cae988999c9ccf7e13034b432329d72946541fda152d691140ba9ec4919a68c0d9419de60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11bf5e7ac0f88033943e15620ede6950a6abed5d7d8faf6eafd1af441ad2fb97c6f3e0fff107394409daed8fd8cdf13b4aaaab9f467f2c6da326c645a51628bfe6fb6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61845a1a069f5b3f4fbb403219e0521cf879fd42753d44d45bc309ff8c88209ad549d9631357fc472e9c6c58d9ea2adcac6f323c1099e122909956799649e4955c84;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15efcef7a02ea0fff26069629a1a23fcacfe902d79d08899e230bf1b59dd356423b8d1458d77c18d8c564f350d4f7d9136144c8db33b03e8ea38cc2fa6c7359a4983;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f22e305c7e16f6dd26f39206406eaa1d461a1363375ec41aa1d01d84c858443a4f385f0a9d28e3dba7ac0d714116da385e1874ec5070063f3a554b1f02c7e70ca41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1750a262c6894f9bee65e5c8ad03786d44220341a099f64dec9dbde3948a080b319003588c4d8ec4d2fe438eb677dd8925659a7e72d2a889018b6a632885c235ecd58;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe2ecc7807506970c4fa5381ad16f8222caa9462acc4dd53be829b00090f12154852ca138a1e45cc4f1b8b24710caceb370b598922a7744bead2474616c69ebaef19;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80a168894ae9733149ca587def74a0349faf7faa42b50f0c08ad24e2fb2726bffb9e25015f73835547b460262014c1ab77b245e6cc5411f278f80741e679b81f91cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ae6d06860f4a51236b0abc89b608ca508639e813ae2368e606349370b42b6914905a7c1f19525a9a33ac5a70829f05f2890583408882f90644c8cb3c340c3e424a76;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c549a2a25e171b01bc81db0d01361d25ccb528fa17c9c4d781fcfa1d1c8a35d1bbd0d41e830b5d87197eaab3bf1f450d44681ba98ab784afc2c085c079e68d27a1dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h57b98cbea09cc2ed56e11954b4aa124e7ef7f6b7b3fad0322419579e7e63006a29b7ebf6e93c07407ed01778aae3e58cf099d22743cc8de6888436fec7c100990e82;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ebed2f18a063d89c7e5c8bb0dc57a4b8f3fe255e570a945c9873849f1088db133f9c089c2474c8760217fb6adb73d9d5900009c26873aa7778a52b69f6c9a5432b2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h888970dbcce25d31a77ca674ce2122dee053d59f05111e45ee1b8c0407663c492e7f19a3b34e43d8964840a843d3d84c4b3372bcad4929d6c19d16827d7daeec1a83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d8bd76200dc0d86471c7e5523828124ddffb24e14f5c71d44f73066189a65d4f541018adcb7d10f9eef7f8a3bfadf7629ddec16d5da710158943d400e44793e9ee8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1143b1d28cfb3a4dcf23f4214fd423fd8b2901669252e4976f58570b87fbb726e9246d73510cf7e4dce486f76f5d511b4600726e3ce171c907642794df1908c772a62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12fdffd01c8d736766aafc965aedbf4dff7c3aeb24a78023a67051a3342909d5264236b8f44de31a82390a08b79b3bc769ce8cac92f3751959e4e104981c0870528f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h144d30b44d9887bd0c6cae5c2d0fd22534e9e883483a6ff8975d67f6770cf0fef41d8e28d94189e0c4ef7893d48c45d35d3191500758e865f22f6b38328699a8f22c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17d523cbb160c1744133c687f3e0a09757e0ea3c71a6fd7d7f953d27da563504ea092a5ced4624a1b657a29f95310a1f51315524073e2c0be305c3c714ff8f9cc75cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h102be4d3e4403369a61f9060d52bdb1c42541eb805ce4dd46ebcb1fa3ed36ef8ec7e3e1339f0d031fa5f17a389c70a3984284ebbf3a3d6c68c0a9effa006260752f49;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c9533a9a633799b81f4a29aa09017d5d084615f4daae6a541b05099bacf76461199b8842da04faecac4adc3d12a44e5f2cc31c1a1d4fe0699ca47fe23e91bbefc24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c89afd7ba00ae0445c50c639237d47d0d95afac706cf1178756a6ba614d0649ee894c20162340ad6aec19e0180e91d7a0a771f7d0fc357bd96401b6c2b8a5c38ce6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cdf076d4c476510266b13485ff0c62e60cab27f2bb2e57e89558ae61ca3657c31eba6811a2caeace005bcf6e4a8b721daa6a5e2df943dee95fd8efff30a89acb4aa9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he25991e15a1c180c5cd2bb1c9b6d1a54b9e1fd02ea7a16c8fc7147c49892abd96b10990e7342be2268d3c869ba4bc57545e92f4f709cee9d3dfb410f7063cbbef455;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f272aa19a94cf90e49bc841c6e7a692205a70c36b2fdd7a786d0895fd78cd9964a310aea0f7585cd1f553ac368812fe5f23d3f5278eedfecffb0c40a8481db5c81aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd7c2a9ef34bba1f5ff651ebb246e69f8bc004791c685c192dfd75eb50aa6027f3359dac81f1282b544e376903970b2666dd39c624be0f22317c1fddeb0e988a9d53;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h229c9942573a31d848bd9fe5825eb5af89a0098e679dfc510b56988f472541fc8959b666d9c049f18f8b48f5f6e4f8f35c0eda71a3c274c318b1fc52197528a8d4ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h45aad9df8e4d231efa37bed56cd0207e5746dc570158b7b7f6b9846b89f7163cdf03ad2fad494520a563b19d3f3d5071a86b6ec9e9c42df4ea0a09521e8c808d2f56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b523f29f4721c1e0c40b04f9229d7a8de832d41001c7cd37b5faf01fd18d5983fe8c10daa9805b8eb4e0961da4f9d0fb12a40300301bc9585a658aac892aa502f488;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfb5ded8c7e879a8d9354838b184c09aa22c5310cd8279e5a5e12693d159acd1ee9288e66db02bba01531e90dd01e6670cdd3ccbbb4f4a89dbba9026bb31083db1c70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a04a14b7cbca5731d1460fc7a1ec46c93c994ba37df9ad6f20e36868ac88efab4d3a76e9a39f44f2941b229900ebfd0a02eb2026c58fbd316ae4f6ac8b496a4cfed6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149c4b6164c24c6b5a898ffc8bde1270ab8ac631ceafdfebf922bca8adb48d6caf690e889a077c097a2eae47de4f15563c7ccfe8f1a2b89851ae413f493461cc9f06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1507f894b0e9a4e9882aa7d16edff39818a8838858600c34ccad22e6858d105d9cb384fc178fc8295411df5b9e1b0f1c4d48eba24b2484502293c2907c7d4dbf82f25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hee06980b62ab895bb73e34b69ee5ba6e51e083340d641d4f7c744526577d146b20b9c6335972b5718bd5d7c2cea04769493ec76622b2b2dd043a5c545db532b5d965;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d01196690c705cd53836cce2e68fc689d39146be06862ac4f5159549c6d84bab6cb2d4df22015404319b97880d8b809f6aacb749ba12243c7699b5faea618f06c0b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce8b846918bafb9e68122bf9dd9bb66f6e283aa9af4c3bd6f9ce88627be34f5c77c9b2203f6f46c6b9ba4d0d12a8fcdabb89eb7bb9a413dc2b1a7600a033c3f79178;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38ab1c6718fd33c821aa9e367859e7f4960c82726e59a9a666bb8fc6c906341fc892a41fba99214ac2b444d3fd26dd8e850d06898f0dd21b42ed5739716936014c4f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce41d1e71c47ae60790441c654779b971d94a7433539a596068b27218676da148b11975fbbb9e984833b415f8c492c6a426aa5743fde01e7ff6dc89714ac5667cb4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h51cc4a2aac34c1d5b92247d12b30fa51812b0057fe7fd1ff470efffeac40a38e12246e5e34cfe71593bb8074ed6104020f435b2985fadddf30b7e9d90b2f4e7f441f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d3f662c9ba102bc0bb414bfc42b7d9069c0d2e9338d589a4bd658f0c1fd8e97dd468700c736c3d82cfaa56027086a4c537fa201ad8c2dcdf4a33b02b6efb4a7b1d80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1036717f7c1ec092ad12af482c0027b82c748a8356c47b96e359fac9822529f1c9d125b2f02ad9a132ca9d084e7d5bcc83918bfd0f9e20d7f580c73f327af1374646d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e8c1a775fd9146cdc37ea203ecdc5e63e8a5d50293a88a47a81ca8d87fa4e72d77081158df9cdb8e41c5962fb5c777d1d362997725150933fedba1135e566cf13b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b52203fdcaf8b55f71b9d65800c584cf226573a379e38a82895bb1343c72a5886a21883255a8ccabe50c1eece76c2b10297b033f7f395a1bd17975573f596edec092;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f7e7f722ae250efcafc24b121b288c4d69836d861098c45cbf43b432d41676a8a94dfd4a7ed7b9820e79f6e3d3757054db66309d551504c5aa7e960ce89c622a559c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h57b1f7dba73555b904fc82e4de911b9d2c7a739ffbafd589d68ac32519e1f65827f3939ac2fb4e27502d89aeca2ff1630de72b869c8debf61c2e5eab74eb01fd207b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d57fe7c70105da596fb3647c381bc365105d7773463dc868718eff2ff20ba4857b6d4b42e3b3df21cccf06818440e265b27f6012502795cc1b72c7f3ab121351784;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1004b2490c230e964a2ca345da3e3fdd88f0919e7edfb9c41a4f09faeaeb449b6d39de6b520f7191a424684e7bcbd9ecedb12e8ce69a45654277c9b48a8eef195ff2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c306d9e5f2712b58338705b0c360c919da1b90070b8e251a69826f4140b424c3ccc31ada637ff7407d6d1b63fb6cf5dae35d4931e07f0512c5e391cfcceb1cfa6fc7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5fe050c756de929334987b37413da69e560470f050090e4255bba386c78322d0322c25a1730d447b2b328fcb12375e7264c13372a63330db7d27ebf6726bda08483;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6668fb9a6e0d25da5352616c24d0d12fca2e2be0b71e875c0c4954b4801d0c34549e3dfd82a0093127e43b18ea1df0404ef257f8896a02bf42a2e46128f9bf1a1936;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h140489992a12fc7841b15a3df2aa475f8be6886efc7c63a25ab27d6939611fc87be27e5d417215c8c330e719ff0d40fad47cdc2dd0520ec4b5a7bf579595337a1b6f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187d50863a0e593bef22ca7c2147b916fbd070062845f177a75a817433625089149c44606ad7ce3cfd9c9fe7f1199c186854ceede1b463b235921b344d514a2e4b01f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h462682fc12649d4469cbc44b80acffc3098ed8f193a5344c82ad85adfc5d42a9bd9fda3c0be5677151e43d920541273db9fad1080c6927c23b3a289562d34d4e2342;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h164e4451e319d31ab7089d33ed7ad7422a75b2a1931d7664ce75be60c422c66bc62ced80fb6f51204ab8ebd50069b9fff52cb5e2f30921ff95d593d9f55626a280804;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9c88e1af36bfa8506340b114d0a246a2f0fef523e670b9208fe7c208350ac78a33a2915278fbcf9f63e2fccfba9669777d9f40cf2af089482463fb490a71a88330b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18573d864d10d72496e9e5b134844d637cd6249475a817aeb5bcd090962372261672420535144c6bf62ae2ec94aa88f9507dc579385bd0c3d5641e3051a61b5fac19a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc073ad17c6cd23798185d1b9033b75d2abd8f233d7742847ab440fe7bcd62f5d0b7687d56afeace61671869b3cba9f977e0d6cd216f8fec0146ebc2fdb4e918b53b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h333e751ecb7c17ccb03a10f911d6bf27d36c0105224806d2c91bf7e191f0aa5e47b0eadca87058fc4cda829196755aa22834c21dc0fcf4793a5f8563098ac0db50b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9dd589812328121ee3043595fcbe43f34d92ce8eefcddfdc20ecd3e777f5a8b30068352b0d174d3350c2e2f8b4623cb3386741d2162f6cb7cbe1531b4980ec2081e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14b3a179a64c92f4edccfdb1770200775849a18532beda8e0356692bad608e677e1fc2cc34d47267309089778381ae13ef4e4bf9ed33877b75634f484c638bcf0c02b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbbc7a3b58e1b678c472838efd69cd16b582358d5833790c2f7ebbfd742fc3d78fbfcad30da15c264eb36dcaa109857d2555df9d72ea18404ee2b72632a4338bd2afe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12651f21e376d23a31e1fc8d2037e95c9516ae9042c3cf01a3450683cdbf522b9fbb53bec8b60def196c2714db9f1be15ed7fe634ce2dfbaff92d5531360324fd895b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had12e6be295185abf7ae5213fc7430fd7d1975d2024b4da8f8fb197ba02273021bdb7fcee070debd15619dc32ffe4c678869da98f4cf275d250ad99d93aa536b1d15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a8dee28691909fd4d9e8dd2b4dc9bcca7e6feb69e278550d0862f987e4dab6f4528c7e09a3ac203541baa4500769394808cbd0ab3153e8a7d3ff6b45feb43f99cc6e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdaab1f1b99d69365cd0f3ed98d01e342fe4ad17f053cf286a4341388d1e1340b4b62d7ce36b549b079c9e8b14ec6b32406934e681d60e6ac24823f3d1ccbbc2ee9a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfcdc5631dcfd23e329d268a9d6777658a7a2c374de0dfd1043c2375e7e00ffc19f2dd00f518bfc1c9f01fd2fc12577c2ebf5211961e8908f8eac4184e72f9e3943b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb5daa996fcfdd20a858e5319b116873ba678ceb56d67b9cfbd7365e30b8819eed55a1e0116e71b8bf984184f41d49fbad2ffab1da83f7ab61d414b57aa8c9bfd42;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h128c38ca5ba6c40c7043ae2d98d95f2c43feea780088e506ae74d1b2bc484f47db88d91d68e62a6969eacc7b82b1b804daa9567c3a5e48a51d64755d86ad43f20305a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14abc43885b3f961f1c2ec8bc128a8276209bbce7ae8abfbb16bfe9fbc828ac8d87cbb160c99b2381f4ae74d116f43ca0b2cc2701f6d734918b88c0b4309f32f5cb7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ee46841cd25f0175ab3db73c963ea09535b0175c5e5b9e8efaaedcbf0e06f92ed9c636583c60c5b2d6f9fbcf29d443b6d7e4c9edc906265d0d08a268be5e7c2f660;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74a90bce084cbfc6240c114fa529d10ab4fb0daae906c165b6ca1000b0393c20f9b5e4fd677a8cd9b9fe8a921499e3fcbd8c6a82f0449b44e550aa1fdbc55a093c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd4bdb6a8295e7ef18ab4ae762e2201466b116cf142dd935233b206dbc5339eed543e1bf7d9d1d2782e0b8cf529e0eac3ff7f8ac351f0109f8a8845e51c9def78209b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19150188192f464d0431ee37dfa8c8aaadb72ba6d434d355887ec1cd90e7ca59e4214d2bfb31c8d2bb3bccc56fd6bd9a5512bd4272afefc09601acd0c016534eb700;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10aa708c4e386748241507a33d4acf29ae122f2a30d8b62b20c93842a5c62bcab206d3a5252f6ace1b86bdf650349eb5e6a73ea411e92e539de9bdc9c9f579d4ae558;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a22fa8f7fb911944d567007c0d05bcdca83427d5d1cdb5c3ad311599a401d4cd53ba7184ff03afce2bef6001299e2a6efa3238a828906fbaf33d64ae4ce5c2fb1a2d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc046cfce4d790244939930228051489fa3b9d2e4cdc0d4d101a9975761b0950e576ecb3f29c8257deb25479f1588557108bf965a071387333553d9147a9260201de2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d3035f2e39157f416358f6b2992a0f6d448ac9415ba4d7f1b1111ce3291762ebc970c8631cacbe195258903da872bfcf07c6a660d9d9779338ca2bcdf14a560b7f55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17b0d21af6845b64c5c562f40d7648cc0d29cd3c0d109ed27f278741bcc82f53aa60c78e453e26653e29e763fa19455c56eb15735a15dd9e2095e22450ca0c6452de5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4dd30434fbeed10ffd8e964ab38025131e2652f8f5ff31505c5dc2001388c708f862e3a0871f13aa358b62785b2d8a5abd23734e2769615c93695bb2e03389496493;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h29cf56cea3068e1943ed024a99d7d5d3cd406b20cc4186aaa481cedfee1edff55166d8f9c0ea4a248fae4404318180c8abb1244f5fbf857a2d7d22701164b65950e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h64f2668ec56eaf718376553d4f29ba31004bbd668a1ce8a74314ca948fede3da41a02f8da645a76f3fd2d9992ff347fceda5df9ae7f33bd0b47a04f90aeb79ac7c73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b6598261bced4885916c313d576d2bd894a16735b6c4d076bdd7cb460ae729b8731ddb4bd1bed919464bac6a706193fee3c5394b3d4d5ec84a3b3ed13dc9600e57be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h526ae4343a5293800c1c4b8d10c9a764e2661c7e598328911dbbf5c26a5ab51bf372959bc3685724947ba570130f740cda89fe3a6f34d29d01e5343d412a3774055;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1261f208a390436b0e6ef47b2f8d3d9c4cb1d3b438cbe8ee46587d848d3659ebe49c78dc48ffcf2c16e51125c89b678770c165998e64955166d233764edd36bdcc158;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h40fbf6b917fdbc56b9516fe4a809272a554c05e3f30798df9df18fb2e7f2248b3bfd65a3224c6536074d52c7bd2840d26bbc445ec55487ee00824775701bd15f5308;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd5e5365d2d46d20636cb5afed8aac299fbf2f2a95d76aa767dae1568be600711da2bfdc803d5cd51390a8074a818bf966baf7db9a3afd62aaef3e8c314d2955c5c38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13855b7376f129e6a4378ad47f8c422d41d8f57d7e1c487aa4f59af59ed3ea5519dec847b4becf864041e52583afcacc92b200933edf5911d9de8f6b7fb086c2ada6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15f6585dde3b9a3b4b247da7b382f8aa214a3888d2b24dd3b2a2ccb56e59df8b5729c2f4a6336015f610df26e30a88f232fb4d139d37906dfd97039b4e21523fd7329;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe34fd6975c974931ff9a3c2d30d2642f41c4a1de92921f0d0797007f73048c2e4044c8b9655bd0c685573355af91c50bb597ca866cb10834aefca36d067fe1e6d14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13a4e26207313014b404eafcbe24963f3df205f9b47d07d5be71c30d22479581b5a7726a70630f93b927bf5dc3613382e5083c03867277118cb2ebaa27a954bc3490d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1adb1f00bcf22fbc9f213100f4906703c3715dde1ea84cfe9fa41e53d63f60e0d0fb498352738176879e1b67400c47efad0f9a7ae7fd66113bd4516a1ea61c9c52fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd56f4b525809b5983f092ccc2e245b8f03b66a12712d4b666f3f5d9827ed81e1a93f805c0eaa126884b24b835dc5a7833f7bde20d080c2d740321f2379eaad938a63;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heffcd2b259a73c0a11a6efb488c51133e8f0f1831b59faaf46363ad71dcf0029ed61714202c1a4468f98350e6d0a905b7ceade478ceec79c097c9d4e7cffd99e8107;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h177a8781c28e110cd7d5c28bf36698b53023d3fff07ff33880d16375bc0804e08e1206ba07ac70690172993446b99e1b821f89d4e7f241e1fed46c14764b1f74b81b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18e2ca4dbf726f544821a9d9825ad4c6e64584032b16765a1d1cb8bc3e6692b324513b1a9855733c1b3725c635a2a6f5adc53312bb5a294291ba0c5b16f17c250f9f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h109d22e95764550a8f946871440a11a3360f8323d599a6679e3deee1c9827b7b16000c230c6e6f4e30b1de8b7d4dda09720e8195f69c102867b7f70880b14c83e6221;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h119ec3ba5e31ad11c434744d99930b341bd8b4f986efa45406aebd22fc59e922e861dc92c1aef96a12e1d1bf2637d9a45a6f594a03e26855d336614643113eadc8c92;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19f11cd83cf6f7cf69a095bfdc615d7745d87352c16d22f61e7acf16be8728df1c56b1e3e871a27de3525dd07b4656100640bf36cbffe945fea1d6712f50ff1ceb2a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e22763723202c147e1adf337ac8c517f77522f989fb4cf998b3d06a72e51a2384f6a3b032d249ebe7021496059241433c795cc3eff1b044850ce40258d1b1b7f1c35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha62a3adbb5b067174905e0a7d1b46e256ce07ba56d30283e77a7d675af4bece3ec1097e15083f3f116c1aaaa6fc7467ab3032658714df816d515f56aad4451f388f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haf6a7b835882ab01f19a1e9774229fd674452f137137961c299e5e6b5afde1aa617115791a869f77d530a9bcfd0210d46ed9d3437bf3e73aa835cc9e56c59af18427;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14fffe048b23a57f2272bfb91e0edc938046393202e910e53a66988dd24e58e821ee92283762cf042e091c1dfa6c0e0f8fa5d565df118673ed2b0e0744a2a97e08a12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf9222cf3fb12d7805b330fe02940ee5b14aba63de07abf09908a21280fc7c72d4fac8807e79a9a65a5585e65cd9dd32e8dfacfad713f3229fb480521092b262ea46;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcb2290246469ec2f39d8538588efe3c8e3a6ad740fd14a8fce141235e6628aa6011d447e17ad7a29d2813155899ab732b1fcba5c90d594a40029968094d32fe48fbd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf71dc87b8f50d553de75fa2c6a8fecb8bc336e5052186d7c9c6b49cc08a79c25d37b5d2350e813800a634302a2084aff0db034fc220683a6ef97cf52b4f67978a6c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h65682d702799d34ba5efd2d2e88f69638371a29c01dad33f9c495986860df0acb9b65d07d652974efa8bf6075bcd2d30a8824aae3ae5f63bed57357d82407c4383c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b631d13768e8e63e85796b55f6bc7105e1f0156540121986568769a2d3a5b23807ebf96b921106a5cf0f85aad3423f994362f5a82dc8ee7ead50fb2f09cd8439e806;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa927b836ab661273c5ec9d8c26809bcc6c0ddf88638efef59b042cd390999d5dcc0222d0f96b317d5ac9e67ec27d58558e6f79dfd062673f8a320f07ca2d77f3122;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6cb57d5c57f266e46fe2b93fad608339433a5cd99ca388b39cb9a4b6bb8c40c49667dcc2e3e3add154adde8a5164ff82d014cac3e8e712557ed8117879c817957296;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17641c9085456368b72c28134a1c3527806e151b310c1e8a57e54898fc9014acbc39da0e971e52b6ccc017bd5bd30ab64bc74152158ad5422f95d3b8512ae5212e795;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h153ef2c6e440a4cf1657a4be79505badb4ce34840b63cdf110192dc03f91baa4e3b7519b1736021fafcbfcec7d6d252d9d381ee8aac5f396bdf9e0d1c08b45072c534;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1adbd49532d40583111dc109a7359b576eaaa2d5bde562c96896e87713750c6025f67b9fcd0428d44acc68e8b958658f49b8a14aed69d6a66b161a7e35556e7d74f0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fe9bc0799641d171a9b0ac036f3b0bd3309bd6742c7f38a301b32b5fce5d499cb2f910462313323706b2625daca0d4c3b949125f5e061e2c1523f3680e71841e3bca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2f12af8f6da3a41031e5fd6effda6e71b7e201059663361b3a85abd1fe06db6e0ebae6a946c44ab1eff55e5256f60ec16df85725f1a8bff8876465f9d1d73970f149;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d7cdc211ec25d16bcc496fc50918a92a6122db7bae1e54399afd7c4e764715fa5ac1d8a19a8476ffaa8cca0e70d7ef8d121d5929117284986517a0cf92c33eed4ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5077fbed878aed7a143ecbd8f0ee6ba415cb950f8a6921d1b87522069e25efc5ec9cbf0a4ac85761ca7b4acd30f6c9c3436a2a49766b8cd6bf582ebd2d91ba267386;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a183d8c11681212e57ac797b0098a899cdb85bb578fcec21788d151e1f8d1b9a5d41c53ab6ead048a1150fa143068f5a865312659e5b4cc44fe8f3513c95be391649;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9b21e1ac8d3e025c9aa777a60aba816e17dd9f0ee052bf066365bcbd9ff370b593cee6f047c307fa1749d4a19b08623b0e95b25071a9feec12d99a136a8cc7fb44c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcda5df61ded82deb8981097a71c2ae105c50d39cddd1fe7175e78a2ffcf175249bbf25d94c396d7ed9e7d79bd4c427deea71246891936e03b77c304e9d77bebcee85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3b5cc3cdffea66a3505c74cf7e6f6c099bfda3c32e46f589d2217508f791567c0712e26d07db7572cf596d2b04e4cd1975b327bd05fff96664f76757e23e909d63a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h897473be917452d600b32660dcbc87eb45cd7fe5d97c2e698cdf59548b7d9fee6b81b21091e5c99f0d5dc13744090739caa40ebfc0264249ef225864c6eb2f0fce7a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190b9d7c2840760174dfb0c9084216e97a3071f3b9c2226a340a05d840cda43fd9bc90a12a7581391171336e3cf6107c617926a65adc93f02b895c95afa1174c3b5e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12e89f1cc09a4bea7d389878c9c72f032f393f010295de628e080d0442c7128efbf7ddfa0c0a59975ab7f7e5cf868cea570e2b507c791da78f305075b9e5ff8180385;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc2400017f0624a55c53337f28682298779f3d4fbe50358c81ce3a679d35caaeb19b2c4d7e7b7210caf089a3d0070e07915b0f4662e089ba07009e53f8be66747d0ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ac817a5c2c8fcc1c0e3a92c0bc8fa3e349edd6a7c58f1e62cd4f34c679608c9f6d94c5a6149ac20995edc9067685dbe91460c3d118da50e82a4e3a9d3903cb25be56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h409f9bfed4154a09cb7d09efe40b01c277ee6e1283000901a417dbd405b520b23ae0a85616770fcd3fae74c17191c5743519041cd8dc4863ace3fce64bb845319ddf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd46f05c679dadb464a4c27e9c7f68daf4c3afd7790055c5c29d21971780048c51477261404c49830d028ee27ef64e4fd7bbfc499a35fe990c7faa648be7dac03dff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f16b05e378ca3edcc90345399bef64ed8e990f56088754b6aa2cafd87245935b55cf2bfd0d5679ac17fb5070e187d5bdf4063f6a84eb2ead22d603478953f263c1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc05ef2a1884718cf8564988b74a036f55cc2647efb9b2f3f8b6762ee8081001c949123020701b66f79f41975930ce4ee9707d9f52039ffafd2722c65556d34852b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1548eef91c2dbf906b07537ab42508f4ed8a6565ff4ca430aa026674d85391c014e6e7fc574fe54e409b1ac2d96a9f8d53711ee94ccdff3a226db12460caa64eca001;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149c709eb056c58cee583c63d263f9950ab17d646731cc72db7bd46f85f66dea6bee92a0624e1ac2377c6c81635dbf611fe9b39effda28c43a524cc04902009182583;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2754ce7187159d7fb36da6c0282ef746322b223fffeda28e86ba19f2a690c75c477f3c089e425dd6e55bacf4dafcd5a74ed6f17c6db86333b5f2ea1e15a859da1d27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194b9592590cda1b75651eb455efd008d5fa5fb6f4e024081c11e7cd554f9d82d11e765481332fdc4846bbe2cddd2db19acd9fb8c2d461b3502a8821660aaaed351f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12eecaec48d592e88672b424d8e8d72871562a551cfd948afd4c3f003740be6782822b6c56bd082fdea42354b91ab05bd3557100ff18c0c8d186936e4fdd18bbc4b09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb8c4ccc98c44949f341a1c2a2ab50a33e1bf7703b64a5a6dd0c42161e4fa4c7d20b934bc8e88598d14b931928c3b44beca0bd4aa27fc9c2de9bba10608d927119fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf7d4fb22b43a0cfb185e7de8bd0ab5c90e4884678c4fb7c272635460de9d5a4598f62d41ebbe798be2757dfa6984341af35c2ceeecbbd93c7f95bf367d212896c2b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h996daa24a6585fa13ad39d62fb4630982cc7000dd73acddb0d8a09a199cdf4b76faa4b504e2c9a70c262f51ec2aefd7c36f06b0d7fbde3915231a51d4c8e0e971a55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hada14f00c9a2a852a72cbde7491a22e056c162939d0739ee023e6bf1a282f689f468a3f040400013a8e4a0cba144bf5ede2c9f87b176ff4fc2226741505bfb6c8a5b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86e326905f11ebc7aafc3a9c67c9e1731f612a7c0b824d8d76efe54e96f9e0fc3a6f4e34d898e2595daa28ddf5fa29310d611a357da46a848065fae854a267d29e5b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1fee9cbec8d801f8c882110b043128594e09eed0e674907b20d2d1ec64d54b673d537f45960b40bdf2edf40c4467238236aea46ca2937980b1c8feb07c9802f9e75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e486494b2e1e1432e6d7d6a3d2f0f3285205a8681a6b9d625f2f7a93c52b0c1af626e7cafe9b47e2dc009f8737a23296666fec2fc944d1eb2d12409e5625057c0cf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f2f07e8fe023a87b2758cf1582759843b7b3057708ff0fe83e9598e049edfcf8c4a3d412440d47a2215092f1a831b0f6c2a8931e00ca6bf40bad1d8df0ee319b0e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb145f22b0614718bebaef6ba28e89bb31eb7bc5f442f6baaf3a319d7c8ce1c8a52d67359ba84778c00b83bec7e8969f4217599314579bd256c9c0dbf47d85a544cd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6aefbbdcf0b4b1cb97ccb946f240aad537a75807200c2d59048d82b71e16c9571b4db10ee4ca7207dc922579600b40c416ae4174a5e4d43bef6417c214058e1759f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b97234cebfc1af309ab38f1abd16115e84969e6afcf39c8c5784f91d02cb86bbd42cc7372e6beea55609ba79701913438652e19834630d8ca58b07116cfe27cce8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cef0543419e645492b86755b0820dc5786cf5cb1b1b99d80f611ab5bfbc28aebed385d6214b3b061ed7ae53721118e6466d35e5f5a191ab59bf34ec40579824b7083;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f6be3fa0880dc8e4ef3d08f201cbc0e17545a939d030ecacc9278e1e1cd925431bfbffe6e83ace53b731b1d7ba2d91979e2bc4f78e160a207a797669e75cc7993c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187694f9ffa0076e256552c3f35efde6367a72689ad7f876a59697ad217e889d7a5c4d52ca5f63b54a2809c39b29ad6f53eeb15b0b98a0b77eea9f456bf687b2b44a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h152247f2b99ec76447473af0af64a994a0565d2b3c87e5f163e750fc8053c61c4aab49938f357b0f9322f181da2c7b97856989911cd65b01061849ff951e1e80f232e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e9170c7d4b589cdf1f8bc288a91e64cc82930426f28498066f93ef5cf2e5a7938cb0c33de9bc5dd18f334db02803d78b1820e81b59b9b4506611d66243e6787587b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69604021de772459280b84005b638b8cbc8de38fefe3e7d490a08f16db8f1d99435c296616039240af9557ebfb45f7b9d7caf7cf5b30289c5be1f1f48b7aaf4772ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a018f4a12865ed5991d7d6f335de0d07b6e1deb7e7aebf308ad8ee8ffc9ac4b514bb0309234c5c14a47918b755bb550bb7bdd77bddae6e81bbbbf8f2d19f37b4846e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a4e8e1459e52c6f3334fa8a35afb22fe004a9f506ca2db8e4ca4a41080933c82cb29867a8fc6bcb99a960b1dca0acb1d591490b3ac25aa5e9d81c2937f3bcc04ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc8cbd7f8509bd349433588751108e9f7e4ea2e68f2910c92f553d800180b9d55ed6a412933975746bd5b536d345aadd60038892ae0b5e162dff4abfa2f79635c6610;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6da4333e9f45929738f92b7320bd6da9ae6dd19b2d6ceed358835287fd9191c2214167d8cc85628ac087d7bb5ae5d1b4ed2370c8f9c73190b8665bca65a7010b1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17ff14c705a9e0b46b59581328c24970b95a3703e75ae37ebaf618be8766a64c2b63268f8f33fdb06fc8c8399321877f367ca7be958f91d69d6b82415ea3f0cea0515;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d272de24c0333fc273be52016321732be6de68bbc4ae6d3741ed6c9a7766f39e8b3a11bf19ffe46b28070ca8d4d0883c8fa64c22666d6b6955b73cf7c10bea1df335;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6b7b2aa8fa947a519c392cb3719d1f42b54b3b0bef86791c819cab97d5ac5424b66f96ed836847d2262d708a26b47d875fb11dbac2b3a04476c6e02f4a0052011ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1683d17565a84c330edb4a322287666473dc62969b7769a3787016538ec255af20c1322c2065e420e8c1d7c5cb014cf6c121785cc5b287971b52bc3eccfe09bf00f8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3f7b3ebd3f6aa69d11b2362a92d70b704a59a6cf6734b71cfb561f4ee2c8dabefafa667f3426f23a7786f66ec17def602d89eaaac14f3291486608df189d93bd73b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1655390616dbe5c105b922fa83c29bfccb1e05f10f7b46becf2e1cacd5caa73e4bd347cc5d3cabb5d95df8472da691047b0d16a8d4c08654d3b2148a0775dc52b6d62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186b4a9a5cc4fbfb2818b8e6ebe732ccaadfb3b0003e2607ccbcf0ea2622308582d87eb206a70e580e1d349e3810cb85af1f3052b088bc712b165291abb8f1a2d265b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6f08ad772e5ca1c263e469c82765053de5dd3f5ad3405479ca6b5ad366fe03f2e313dbd783d7279001e2389500dc352be63730886492a20fff2c6b8b67798e755fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1efd8120e4557cf9464c1865e80b3886e8392987a078ebed041eee0be01818c6f51c1592f02e83abcf75ec56ff3cff808d345882ac75d21b76de4ef8d2c6ab57112c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h154f12d3e1230ea4614581253b7614c08789bf1e7d9cd18584c3b044f1559ecbe37e97b5b17551e4ffe10bd3b4cbd8cd6a3b126acfa174dc1325cde8c26e311722dd2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha0f001e2a5a8ebd0781874473650e237e164325a3d9bbb602f9fc599beb3dbdbe81c2760629534fc78ee782dda5a2d734546c28c92d4d37a466b14408439aa2c4286;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h199d65faf2708f3f17d857ff6fc4fd9517b13d1878b552d4ddbe4cd909936744b0eb144425a37a85bd6055c006db21324cc7033e6618e79b84020b3cef186414a4275;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1906df402828687b755e55fcf2a9fbbb0bf02a3ea8bf08077a855594839caf06d2567794c9fd7bd635a214de3779acc5be2d9919fc6f47e8ce2338336f13e70be06af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bdcafc8130b9bd977001bd54aaab4553b2cbed7c15897378cfdcfec81d47f4a111d388985207600cc2a82899d5a224e62dae1fe03d62c92c956612a14ff1b8c3e130;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1809a5e3de9754aa43a29f7ab91e0eb1b67d1a564da503c9080c4b92467ba530951e6b5bde1d64dc014ae67edd6ea77d89c21d7857c73cbf53d923e635d3fe3558ec1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ddf1b74fca66299da0e97ddc5e684b398e5a612eb7d69778e2dc51e035b8ebfc68077697b22afa578e7cb7dbc092c975e8549e3e98a37e6cf68beb6afe2f6d681716;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4de8dcb60d041ec65d1916262c6f5f7d1705ff6d6203af4797a29af4016a6c9942090b5d16280377a2245b076704f7ada68b4dd21ea499b18d2633716f3cdad73a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a604a4fb7c353e2fa59a4f99a1e2939a95730ac99c269ba0c39d8ba6469d9ab0ab5524c4d0657d730dca1d5112e96f4c1f10679099693a2926df169b6803a77e134;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1194826b80200a2297299cf28cfc12787e909dee10d2b8fefd5e88d9f09f60705daa0f5f9602a33a1d7b56b39fc1819fe87f5f50e788b1d7b4d11a6e1c61495a8a6eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc4b6bdf1a42d113ba83d6fbb347bc04c819663ba232afd94f4e16564a4819badc4f222de0baa7c2d5b6fa20aa904ef80d29031d87e6354139b0c6f7163c52d43fce7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc094ebd365827cb99916d6337ccb2dd65faf5d4d6fdfaf7946dd96048525461fe2e25cc43404227f94ba58e37190cdc1f96abbf56083331c5d7287d32cf3094e270b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha473e3a34cc4b637f65c29c00a91041e329960798128bf6e529ad9780e95c7cecd10ca781b7638a6668634a28379e6e19c2c4432f1e5af728ffd8cf041acc48cf0ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c143b2ee39fb166fb7af07faf3672b6b601bc38b4ef32789882c048cb5cb155db9ae9420d0f3a492157504cf33d0879d11cf71049448a033d37ceecd71c4e54942b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1757e82d2abdedc0dd4f313df4ffa9d206b88c0b7c08ae5f75385701c76087d74929e0cc530099e446ea61005fedb3cecfafaedf5d06454722ccee95ff8259666a644;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1188d4877a167ecbce86d8405b30b586448c0484d4c7c63659de68d77727f3a16af9cdc82ad72415a5d384cd6590396b74a09e7882b3ab461700796a3e868bc19580a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1678fb8d4e3e5d18624f10181a65e84c89b092ed7a1561274da7f6ebb3aa4c4b8a359640e3f0f4071576b99e083b3e32af8488325f58e8f9eb619ba934b65d4c4899;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120985947f5126f762fcd7e4a1845effebe4938f3fe34be301de41b777492c8616df4e7170eb06d76622f40391f9215be90a418c02464b47445956d4470ea3ace8dda;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h40b9e47b8c81e6255137b2a8efc09b8860d47a3d2c999beb232626d1d77b1578d90ed9a3074ddc349517c82ea5eac753001f9ae89a85dad913e8aa9cb487b0c905f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9334f33ddb6bab47a746b5ced4d8bf5965af42469ebbd15c148d1940a4cbf75970ebbb0c76c485e3e58edb99cad2c84e1b4603ef8c7a384f30f5c890f9ec60d249bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13586cdbdcec9c459b13ad90f9eff6e31e11db2d70e94f3f99f69068cfa87425f45b94d0e0a70284ad27822f760285acb63ffdb20f4d671eec127786f9557fb622876;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e836f54aeca9dab1d05db7461fea12aa64fd7f568ece77a602a807fe2a9dab60d95c751e14b7f36d46d485bd7c3e0ab0e666adffb9933481ae89414f3a149d069f4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h125acd5077534007680708bb8fc8aa5dd864954c90e95a2e531f8b58059bbf3be59b415e26b5b18b3aba430aed4aaa2fba696410e32d085d6f64921e051403b68e01a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a9851ccca966e2fb263428a18de6a3e34b108542068c16f87fd26b52f75630b36dced96c9aa061995ce0aebf1f6ccbd134cbe2f88845e803852ed82d3c041037d15b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc4a42b8352e74fc508272b8b3d478b4c122d38c81fc64eaa0ace0c5345611e9caad4de3368f54ac3b11ca380ba267796b2f13dee3e33ebb0b17fb9a76660f31afa86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175edc249cdb1cb12d5a246d61df591f132b8ccbbc2f89f9cf8e7c7917711bb17acb4d9a95a124d765cff1848486806f7557f24c895df9ebff32e372976687597d97b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186aa01966b6f5d848fcae695b83099e337a3cd34752b4ef3081f9c1dba28cb39f892c2ff9d2f45fe4a1a3f6e968d837f0183552f66095dd0af33a341c24b37367929;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15060c4c49d57eeaed85dcfaeed793bb19e6619b1bddde945b69646a8b604a8005292c5c7455a899e09657f7beab7469bbd39c2fef871769b02372557f4aac968361f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e47fa5bf8ce813095d69d467311d40528aea14c9ba17e7f3958e9018443b2ceb703264a7df491e14d49b39610f10b0b7bcf0f89746a5be1899723d538370946409ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1583ea16aeaa593c1e8a5087f65ecf78b84990b3c1b6ae631aebb110dcb3bbd1d7a1f0c962fe53e6e62bfb5882f8d67d2666e4737c2d078265db5a0d27a744d7f502e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h102bb3be9e1b9902446ecb91dce76cd500296c95092e7ce380986ea59fd3dd6e3bd7a3320e51551d2ae62f1e0bacd28423e0222a43a04fcc5c791669f14207f45feaf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aae883ef745b25be2dec62feef89d2edef5153214df1c8384b7e5b4397086922967827da63dbf225eef786f091b00d8d5a55fabec14306c25cf6181841474bc15d4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h189ca5415fa8510e99f1f2ca5e98585f600872feabdfd3e2ee277800989f8c37294326f0447e00a40103a073e5955e7bbf614d7f60d81548a183e6dcbd6cead022221;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h169ed115f48a7090692dfc7ee0324b0017c9f0ce1bea647619346cbc32e1a869f54e7a9c567ec6ee7582199a73c2bbf239354cd1bce50b1e31e0185595ba4ccb145f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61f449f181e6e9e9c1391ea09bd7cbe8f4274eca92dcd3b15aad93f10281cf6adca1f61a7b8848e6a6c39799c4dc1a3fbe12a257cedc9723ec74615cccb568278b83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h168aecd9e9a1285cf57d51ad07a02b62a5602d7e7755619410acb2b2fd3dce3b76ebeb525ca52964946826117754aa37600bc19a12e7c9efec5770ed333854a3c1e67;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d4f3eec7373851b47df4438e9b3accb15f289ff2d7699abc2d0c364e577970b1cbbbe059454719df4c8e87367b043dd3342dceb8f8fcef113c8bcaac92cf44f5759;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e100d640c7cdbfcb51caa54e06bf5c40b161d71e3a735a24d2defef8837e86d09fa8bc0ac156f6fd5fec56689262f919b1a70f63a31f79185f28fa0fa07f9ad44ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heab8e05afe14117531df7b76012042716c0a8990c2971677ae647d31ddeb537de551c544543f5a3074e3eb489f17431455a1092b9b593aa0ba72e0c49db350a4f683;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ac7d3fa5263e77dd09f89abcf9e8c4332f14de133a7ecf80b2fd0cd5063d634cb45d97d55539d979392241ad778680abd229906a4cace2d26f699f352b57a905d595;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171240294a19b2213e17c449ed975faa8b990a145db45f0ca5bd69a1a2b69c68468bfdcaa61430caafdde8f7e2241743f515f70c763ff622a5e812b7d60c9f064e7cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e49bea5aae7a7c9318b3e781177c3dd972d17a8a5550ac23f188bdf6589a63ee96ecccfeca96823f65db4248f600b5369b3e281d50b388a2469b5aaa8a21095c3bc6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ee41bea4e19b1ac98ebdb32c29fba262fa96cb04a2d641b576ddc1865a24f8791038f249bf3ecc206991996aaab105c3a191363204ae51649bfac5dc7910b35568be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd866976ab8c97043accd75aea4cc005f551282e637ed4049026321ed80ee6c9590daa7ca5a050bd2f2c9586c9bbb378db518b0f55f35fcea1626d0ba86690b38d95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ec6eaaf83cbd1adc456dafec3f37a4a72aa5913edb69d1a84a5d2047c171f3b2311c0bac07072d33d706532a115998b0ca56dad480c7311988fb0bd9bcd380a0e8c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2b52c97194883eb846ec2045f14bccc43d80f462d5d456355823c25009f85e17b806f3c9ae7d216973b0d6f6b23d866a3b08aa98b7b56c68a212783b3df2d53cab1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1674b24f55223c97d5418f261c519c8e273d5b9112b1f38bcbc0000a83106b20410272e3e942489dd7eb3e70abba348adee184fb7eb0e6d08c9867d54f2694307a71e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e54c9c031be676735f9a5a147657805b2427b004a4f11a725ca29b044646c189d0147a7744a980ee1b258bf71bfd3dff8481f806bb869004ee0417b0b6e187e55b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h21d8a1d705be012f3d2034f3c8d633e53ef6e8c9ce669c15f25b5d3e54d3fd4deafda8887e7d233fb7fcaa883767ee46f8305caac33296c08331e7505a4296b140e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c8e36c804155028e8f5dbf20af099b7d27cdfd3d09502467c8704f32409b67e3ed9848ea3b0e86a0a5c7e41ef3cd68653cfb04d90113461bbfcaffd27d2c6f2befd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h481515d742119e1b73f1ad8db7184d552376de19efed109d648d37ca28832078bdff4af4fad310c96964a0a1ff1a8f6158b0ba9af9bc69b53873a9ee141b175140ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dfcf2cd0684a711bd376ddd079f0dedf21a185ef8d8b91a746669988ddfa28d02f0f27b71fc2ba711146c6063ef25d2716f4d567a5233382a64c69f3cb4c51348665;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d5fe43c0dbc36fc2ea8b450995e1692ea8a2bbb56f1435e8251347f687b4cb249d7bd582ed5a3893cf40cc3ec840674fd73ae99ee53bbb8c1fc26a6b6341c5fdbb6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1103f2431f0270f60cb85d911a07ae4430ddcdbdaac9a938809a45cdaead40fc637a3cbc097f4e50e01c9ec64aac81340153b3648c5105a1dde9d5e40fbc3a19f3f89;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf12db4a701cf918ce63f0d64d9b96cc659f4c3b465e4f9d32f98278828ef19711194439d759e7803498007b3ab4a4a9c1247dd4b0c7d787adee8c655f28d8d40a07a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9c53b0bc91dab710dc3225d5c72c871c0df3b6c89b4a183394c0e590fa162848db3fd72a56bfa1101d7c2d1a2f3cf4e31e0c1d3cfdcb4e9f1ca4c25bafbd0d9fb89;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15f518f89d55a33aa7e42d70659d514b690d07f8e8388c384d50b03cbd1e238fa4d33c80826c76cdd1763a4635bd42c33d3b98729f637d6053005bc8ec0a3628d211e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ff3006898bd3ab876152928e1879fc6a24f8c343896ef0a72bbc3aba52f2d3cbbac9cd4ad262c9e41854b9189e5ce8b999a2964e234e3c7b1080ffbd256cea15055;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d67d3d0884720d6035b21f7ad0f528a903f4dbd4574f88ddecb503c1e5eabc3927cda34d258e1308e6d77179ec1fe622e9e53d63bd09330d4a7fe00740f2cd80af38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186102f0b3d011c17b3724363ace2e73fa256febc659c01a0ace49bff2eb1ccf2a86fe6e093fe40de01e1a7b40337785b17bda808fc9087dd52b32e4ad99a342aa600;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86ebbdf327f09cae4af599b345682e6d2f99770d1aae268e6368776cfe98af17b6b28187f7547dea3d1b8bbe87a251387c7082f1964357ed50c474a60bcfbbb55fbc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3cad1acc2bb13bc46c672f78745a1358f12d514f3180a993734f2a1162570a2b971b2153fecc0b1d292458f2621cb1cb06ba8cf7744a88dca0e027392d27c3fea05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90a6b661f376bf128b2eb9683946ad8c2faed39f288f73912b16219692f2bd8104da798f10525fcdf6f988ccafb58df29977f9e11e6feb2da41efb70748decfd8720;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h126c1d7a224e9461d7a12e5b846420a513d7ddbc5eecf8b1d24fa5c7df4476c0a9b91d236fba7850c72a50f327d5213b366ad00247680a7244aff963b05119936eb09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b95c10786c3fe6afa3733d8d16dc03d748eedf051be262e734d1109eb26e3009aad48bd0a2b8a35143a5a700491f289de730ed551384261876a151ab85cc14d3f3d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3833df335f39bb392848237e351fdeef2b7213acfd8de856c857f247dd58fc09bb77997e588719b4322b8cc29fbaf8b32026149a38244e89db0412c6db0e20370bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd448755455ba20cb1da586a9167d293f02509dfaef5f91949b4c7970510d36eb6dca4b0eff09a775f9c7181be2c61e727fd484a4fd74c855b30460a045acda1ef9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2386e79b29edf9e15c6208a70289c4be15f0c037e8f1356f7f2e96d22ceec4318ea027d480e12f944850904479e7f23fc49a4fd3057409b8cf33b88e902db263f5b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7934840415507e719f01aaf9e920ebda0b74cb43cd559834bf076e8b289e473bed8b50a2946220af0d50bd5163eb4f7f27c0fdcd981e579d419bd93ff53726b5db4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc5d951343e838903549ec29434caf004900d1da5902c32f3cc7a69a8189fe383bac2f2299a83f5e9f1d64a2022dfdbaa30abe6fc04a8c407a406e739db6020651485;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60c25559a749927db6a9251e1e820edd9ae5cdce0c4f41cc1501ad74c0594c9b36273a0870bc41ae8850d9e859ae8e39c80a119830602fb6dc0a8291ff3f7d2c5435;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h106fca2c19c81256a4e9c74117591507d7f5dd471e0e4e9a3679e7cbe97c2af2e4f8da9edd98f04796306add1e1e4d51784abe0c079c2d5ebd84ff66fce294f181d76;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h155602512a6c6850098f3bac5a90a594938c7d07e72c3bf366b920376e29c621adf595111f6518d5ac58183a41bea44c20f4bdc2ec7a00234e1abb9f4fee414164b87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h22754ac0758e3b19f6c84969f02d35126075e17365fab7cf8d8204553886e8489f5d1dc9bb959228ccbb821ef8ddd7764adcb97183f86f0ba6431473bf4ee2ebc108;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149118e047e3a3050c7e617e7e62ebe4246849042a2908db1a2e9879888fee9ac0cfdc94eb05ddafd69d4c71dca83bf37733c501c5fd9ebf4f882ccd6bbf09460a7b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a2d64163e1b225caf072e657e3a1e36ee9e3433dd32c56f45844ac2a43fd19845b47592b82734415252d876128d256a2c8cfec774f0d901246316c984b677c1ec84;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h100f92862d41de9d2e72f3652d0255f266277760e8d602e54546597b716d5e095e87eb6da285193255d4c6d6b0b05a9fda1d666e8ac4d72024c747d9b6ff3640d36a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e456b420a6e08daa099cf779fb778b25bb010f6896c587b7a55853e4defa525b4c5b5b6bd381b78832e024b31704d153f2948afd8e74c5923d6d57a962a2389e225;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a2bd39b1d85fd2b7bc17a6cd76a2ff528e79d984301a7fbf8434ed1f1f358bf424941e21685f13e23efb77ad557b3d968a398fe1e40167b0a67055789ecaddcaf0b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1999e856ecb99deda11d9349cd14a4a560d139ae17625d898372d08d3a88ff5a034f75e5b86280be3a91aa9645ba62752e3c4a7420c4d8702560bc74fd04d5ffa9dac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10152426dcfcce21aab395eac5f1e716b93a12f1e60c489208f13fdb54ade60f83e0f4f56a3cac505d1000accd60fcb8bb8513dc3e88e863a00cab9fc31678df52342;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1794bd42ab111f4d44dfd7c4ffe7267d5722aa42ea3cb118518f2a7be643ebfcb475ef0b38ff6a92d671aa805d1c9e84c57304fbbf8191eea50b932f88ecee7af95fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ae2dc1a5c970fb32f001e939027f4edd1e299efdd1d1641c324163bf1c8efe563774ba7f2cc2642e38e41f8f9f5e5cd3f79e935490b29253f5b23391d064940b5bbf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1646a58631fdc36728a753677d3cc75ec206796760e21d2ba614bead4616234fc9dc7f3f342b0d7584c53dd1314f266736c2aaf12b08ef2809f3f673c52590a45de34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24765f5772d8c5739d4a5126abac32ffef99cd7d08570beede4389c29d0e9574e8a5bf404b78ac023e02070a059ac1689e4ff8295765d5961f3743906aa93ae2d6da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h727a02965afcad324968f82154142d74b3a5ce3f0ebe4e2f80c47da2df88ae600b09a99679fccd479ee0f95c7e1ad2c71e4ca66c77ce36ff024898510ba3dfd0cc1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b56e58bf9808a2aafec3842a28f2b76a59b12b8ca0b9951f3bf78635e475d9b225f74dd39363d2ec5cd00b8b76df8a3cf57dfe8a99535311d21c53cfae739a56dfdb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c3566f021352b07ac499b79ca90c988221d48f4c134343e9aa93543c4223e9780d9405428a62b66f338974ea24a175f81bf096e18b6066b32f8f7d79edf444c9c22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfddbd1cab531c9dd68e755ef16e8fe7a68ab2f0b57a33522bb2ec5d137273c34cfe2557314dfc7dc682f5e734e0a09a7828ec8e78cb8d825b3f9e588ac347c962198;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd6fd7bde997b6e2e7f5c97994b3ac048b3b5934f5a22135462831fa170989293b19323f9cb299c4c49aa0e9b5db0a3a3c66487958654f4a0cd3796acdbaf14df45df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h20485d8c01b85f530b8f3a8c18531819662bc915a2c892b592ec81a8b224573c2fda63a1e6ea23ffa8dc432838448d84f3e9ecba685900491121d05559ac16620510;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6b4e05b489e2a30c64d5790028f8752dc26d45a21ce069b9a550f19b3d07eaa42fb8d3c896615ce78b68960f6cbc0946d89f6061ecc76171fca9b68f3ccbb9646594;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd8e3a84a4853e01897ad7a9d19d350c90c004ba21eeffaf0cb24e3979ef5ab691abfbc3fe9cdeb1fa2821da75e36990fc6c1fb04842e90d50caf1e803cdc1b94bb14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3fdbf4a46533198e4c06959015ec274796652194909cb9ba53d74ee69a9f53d23d6d4db1a1ea9815f11241ffc38128abe1791154d3d7950f55cc508d88c7a82ba606;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18cd19dd8d786c96d07cf96f64598dfd9b3e83ce31208bf144164a76a3ec1f067734b52623c82d1fbb6a10a7a644c738d77170062bcc6d4cc7888c9e7766d017d26f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6a20b68d48bedfc6fa3acd94a4f5c8d43eb688ece1eb7d263059cfc33fd8f56b1e9c70325fa304ae3a1db16777e42ece9f868f72d9d02fb68d4ed5e7bb0d9154362;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c00e9d0de1d8337f01d3342146237a18002a10826cb1a99c33ee6706f50faa5a438384b0a6b5c746a164a90ae894f572f89a92dcb8a9cefc55589b5282ef58f23d91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129b16a8541bfc178f129f5dc3784ba686b387e0f67565b164230dbe85840ecfa759cff15333b8df6a540cc081f7542203574faf92d36c07f3269c4361d1a89c4ac5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h125a72b6daf46b1e7a83a185fa834c74129e349ca30aa51c0a403a448f43ae9fbf5a665ba1294ffae1702fe3f6acbbbb25131afb4490bd03601d50bb9f8846525268f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd14f116391079944145242d53f1b38e7f8a175bc78fb0600025ea287132132d574921d6d2983c1df95be3f18f9796fc2c6fe11f85a0d83d91642419f7e771162157;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15ffdeeb6fbed77939ada106f380ec60af316db4bb712c33d1e3a785340557f3a0aef0091cbc8e3d200fddacc3b5ef244d34b60e395a0d18213ae212ae956aea9db7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf74d1fe8b43b43014f8bd599f5bc4389f337cf9d06edabc899b7d7ea22f10cdda5a0c45c7fd1d8ec18927f2fd4e1da34b5cfc0787da1809c347ee0b312142a7c6a2d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17ccccbca5602c9f4944bb52070eae601722e36b0ea4fb5d4208791f66ba533a2b984f9dd49b752e3524f221c5d85218649255bfa401de5f297b05c05599d5c4f892f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdfc25b9dd60729500a5826937da242f9cc5837d97909a1ccc45dbe847d9123b0cea2b1e28d6424faa057bf8a534fac7c80aa39b18e5953a29e82ce6740b91ea7f5a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h41e8ba707d2245fa512a42e698db8d8dbcf5265b96a7c293596cf3d83db7e2f37e5734c33f8f0652f9adcea9202ab04f45b4a7a1e45e815b333d4bb18d6e6c6d2594;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12aaaf6785c59a3e6726d347f1599326ac6fba68ffa45aa2545d7730a75df1d9e9bb25e4808cea7b6a679e385b8637c0abbdc953b2f420eb1e3a937e8478a57da9822;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h116d129b34f21f9fe5fdc370b6056557e1a99e0a8b489cde3494fadce72652e9eb697002110e2dbd4dcc50c4fe55e5069c5f069c28089c30be4a1894ddb30801d1a2b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h124537001da76e850b59e23ef4548232c9e88c3951141a30f61a7ab50639aac1aea6ea6e8851773ddced48f50b20faf15a62d8ebc2443b418d59697b4ecf08792ec3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h153b1d47516a4a341a83b862f785dfa93d786b435f018ac70c69044a0e6e01ef5fbca9c87805c9c79dd59a12180af708ce848d46a785d41a1c8868f9b91fae1abfc59;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2dc5771204159dd14ea98f2582d9a4f5fbed70812f5dd3313045c2dfaca177384fea42e8abadb8cf38d8d601c8e6cbc64704d5559b650cb9d920d8629c6ca3736dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0d9e21d92b20eafcec35c80df9d5d7f9d9150c8213c18d16a0ec13e5de7d28650d4fc7656ef69fcf4f71a474b24ddf6297bfb2da9ccec7302f7e4befd22e73e9bfc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hacf32fb64198f09fca980cb1ec3c0b81960d0a95b87efdee8b52225acd07ebd8f1fbbc251a969ce45238e408ee51afa793f48ffe33a7a189266807c26f64f038164f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9c0af71f7fe424a813b4104a084a44aea537e9dad36dbb9fc4753cd99f7878a161f78298e384e67b7093cd49caeb6c0f1308bb604a97136f55ae4223142fe112374;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2169a0ace8c8e22dfc80cbf4e7beafbaf07f5add3d245b04be495db4a1a4d128cf12c9bee0b8d7b6b77e0a3bba40123ff5c3655d5849faefa99085d90cca55d35a8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c0fd605f899dd1eaa8b8a291397787d78b4e9da9efaddaaef5e7f7658509bf627719ae29bd87121fa0d1fa22b7d4172ae7049056a8863def388ffdf0f719ef38b96c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff670c366f242c1f92a2781a81eb80a42eeb846a1d737eb1bddf83c3df03441cc4c2f415b11a7c46ffc6850a5e7fee32460363d56f5740808ac9756e57a927565921;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c160abfcbf61e1f03792a58531afbe53afdd93b0bb7afd25ab373cf72701b6364f485bd058efef7aeb791234d42967bdfcaa795d6e4d34c1e196c6476e9c8186f148;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17fbe3f79ee15c17ff36940f42168d773245b3d23a0f4b1ce9227d687c0d5c52c7b63258a5c54fbdbf935c04517b4dd38f3d1f15c4535095269680e3ab8c8035a08d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd0bebd22bf234663bd75017306d586c87812a71acd75aa3813d65185981b30ef329c56fb09dc0c305d4443bbb2f3a8e17d86e3ce4b59fa0c48b96e74f5943181ead9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad816b27f24101ce1e23fbad131243c516c56344cdaa111fa97f578960599469d34cdafef34c383f344fcd2448ae4c2645c76eae739411ee34e42f938bdd6fe2c9ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h124536725525b962db3f79fcfb0ddf078507fb31976ed7e72ce4abded7667f6a832e7b5a37db0a1552218713c403310ec0b220fe2647acb10ccff2b8d117dae71b6f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ef0dc4621c44b91401b48c3b6c3aeae0dddb05e83a759edb52191b87d49aa3af50155f8ac50f158e2791e224f0590c55a6f9b35870ccc201ee5bb03e6503ce70ac2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e5b281d085a52453d31afe346dc5a6bd5e199aa4fcbb8acdb9833e8ee6d5e2d48b12004650f57075bf93b727d537230a2edb314717908b3b9eefc0f5218eba5b64c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h584755700902797e1c381e5b8ef894f874333fa6eade66eab597dab5f9bcb815bcf324f2307fa36af6038fc2b4a596a3f881d8d79618bf745cd4c68aa6b713b54705;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1060491c2daa88d32131870c924c2305aa02719dc2099e36ef3a4c2a09b2c54fa2b73359eb75663696f52a6e0dafe6c923aff8204007e8ffcfd4cba4e2f496a0657cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h692e0606f54894bf2ea3419db6b28ebebd720007fee5ed90f231bd96dc0886fea405ecb5fee767a7690a3917a61d62846e88374f96809446fec286c88421feae1454;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h925745c1c9413122db1c1b9ac10c32d0a01901de9f65644639002740fffa062c66c877746e98d6dcd198bd9f85be1d4dc96a5b1287d89bbb0dc43c658648aadfd162;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd82109cc2324c3f9019659b7c9dae87bc33ed240f7cabfd3afe483db67734cde8bb749dfbca121ac93b49b681598664d77195ad51bb4732704de10a37dc82fd635c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha22dabb151d4f619b4da482d13cd625eb4d84bd8c1814c3fca918ee193615a76fe3e91bda686337889dddc6507430c7f5667972a0d6cc8f806cdead8f31666888cd0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b10603e4b637ce2cbacd9030ff2a44931d9ffbdec7cad8e8c9c605cd56dd41212e77db324415697b420f3a5d41af06552c14c1f42d8669bf64bbb3ff29717cf04678;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4817b3fc3e22434558efa0568d8d9745fe2f4573f89e4b0a859e90cee25d73c6179f4dcd5b8bd68b690cf25316980621258be2bbbd4b6833d5dce880afb4970136bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h184b6f1a02d000861e0635c6f09e413ad6deca6acb0cc3b097ed65d29ba93eea6747e39733f48b7ad861eb611c21c0815083f2602c1b46d9b1d9b315ac7657c878f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h25bf518b77e648c937f8cc3ea6b0d9905a70e4cc2f7291dc36baa961b4ee1530af0bd0e729ac07075bc3ef30bfb498585a03139b651bdb1d8e583ce6e6b17b506c6c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h474ddabc6b39e125ad7038ac1f7927132e83a3a66f5356f8e12445c8547710a0372047f3c1a0061dde0c8a43867cdce5313bd5386e347123e6b9699609e21e65fcad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b563077390e0a7339c036a13009ef90f373444abeef6cb9d523beba5c5bd007089814ac93b79b1232d46588f13df60b54cdd9357250dca7b0601c6708e5c2f530006;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb34dbf8ee04ba896180f3db88d8f8b7872958b5ccb6579ac43a398cda83013453f87893f8faf1bb2a36c9afdc8fe4ec1b02c580d6ea2e3a5e77087389e597d42d657;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d634d5436e806a89ca0ed00b32fb4f5780ebf845f160a2f866640509dd703a81097cee81b22e1c830bd36e6d4d32ec6669c2ab683fb67daf7ea13a332e5ace6b1d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14c8fb15faac1d2b2f5a3390bc182b5ed3478fa43571fff3f5d1c3e6dcbdabaaf5902c7608e1d7181ff4115fc22344fe034d6657e644cb4b29ec5feb20487d27dbfd9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfd2edcb401b365a6c22530a4f2a761d197175e5679f230414e5310ff82c0c269ca4cbeb30b604f5b270fd0d710101c369a19b7b58ec822ea57ff8395f22a7a931047;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2acac3dfff8e4e280b058eeea340329b30929465664b605521374863a25572fcbdd0f85bf4e18c8adb253672da2584a786f6418ab683b47df73bc6b5e4d4337a125;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb0fddd464f17ba2bd67b03f55ea3f718774117b3a70b4032e8be296c483091033552717ca561ef2e51ef1a065d03bddb59bc5fbac7d9411ee63e21a19721aff188e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h918655dbf07c7c3a2a549eeeba5475b09d242ee3c615d1ae5fbeb72327c4647a0d24ba9a963df4c7b2f00929c3d7dbc06d7a58ffdc27d8304620dfc0471818cca647;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h123e7321ca685ee7dfb842e5c262c9ab6de0c1d981ab3b6f85b97cbbc161cdd8de1a83e44334e90c2bea4b44b4c82e1a707e7c5f32507133f28fc0afb50af38caf7ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6b1ff8c54a0aa3547841c9232bab76ba7777eaed5f03c1609dd2406b08a204ec190cda28bb6a5a2e3a72a4642985c665e2a5764522b8e88ca99fd76f256562614a4b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1995f86cd4d0453e11c3697cc34a9042721526cfbd86aeee27aa78702b9fdbe876bc7746feecf23f084eea320e5bf21829575e6864faa26a7d53262de5925d44280e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd8ad1da5bacd1b48bd37dfb6c2505b167e3584177538c05dccb5c35c5d670789e0d199a257c3aa21bc991f51c91daac48fc5037413cee4dab504e5b478f8a7a48de2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h25461362ca6f30cd476f81c1786821ba62ee3077f90f0ac9a9a2548d5a35e90664bbf129aa255c45864aea4d69662b7f202bef92299c5691c16c11184c5bafa17238;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed12323bdab35b96767e334f0bc453e2ed549472b1249aab90ff35ef4773a8967fda609b0c90cef8e41076c28a0d9d6498881945c478074d83cc71074a1671925042;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c03306f46c396dae94e3e10d13304a0d67c1d36bd4712969d3a4115c350aeb8eb7a57b9aaf434fccd15dd128a465dce51101f5947701f61d63290f4506937c905ce5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3cce18ca4019c422c130c59d63e5804400c8e3bc09527f9c2d96cb7c63173c2995c744479ccf2b880100d8df3a15bfbed5a063b9b2a18cec7ebf2e7f1c4074d4ba9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd37bfee8878e5bdf089150553e85a1a8bb0c9802f229c5532df15c98b44d2c1cbe683857399cfcefffe968941264c1637cd329864b1de39e3c6289eb3b1380f24d76;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfab9ba0b67f0aaaa03e37228e044e7cc8eb3e46602853db665e2ff8f297b63c676a6376e4b516aec58f3113d4b96a6e20596212cbbca1aa243dca36487fc50b9c1b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h31e515281c940553fbdaf0b19e321f67de818f48c0bd3182d462d1a9b19e1f04af69330fb86a5a1a0ee9ec65a190bc91f397f31a37bb1cf197089802c5d466638b1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd032f9dd6e8d6d6d11c2602f6bfcddaae56153f60eed24eb8c76fab03976157716bbdb0cc40e74680db42f10adf235298ae74201596a691283835614fbfacbca471;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d2268f4f0d21387973d0526cbfd3936fc3104658a7c45dd001a2c38695dcb2ffc2ccf46cfd8c8b49281c916b6101088fdbb1d39b2fb9a4abef39a0eae652ce76cac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h153ca9cf6b9dee0cf9459e7d2d9005da024239256078a177f63709232417b2d05bcd78fa95e469ae7d6e32b17a8a9fb327c088f8b63e06a54f8dea6500f84e3e65a9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h117748c2ab7ec8a94b0998514e6dcec68ccef2e639ad7871f61ccf71668ffab157e2d3dd9d9263143fa5bffbd6b2639708ad6f339f150bb2882291d6a57bd419904d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12e736956847810dd7577e403171b0c0d45148f45f733ceaa087a45101437827d927c5c607281a836bda5ab464786d310b9585978e403df6442147bc7c34a7c583fb9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd24050e5039cb4bff91996046ccdfea33038c941ea1b49c74c1a6705086ac3cebf5142b35501d6aaa19bf82998b83ef0c3f9e7384d2eee66ef3fdf0aa5eab76b0fc6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d5e5967dc6be5e25c96dc2e560af9de9f446232192e706381ec46991ace95593caf25bca2f3d696c3fecf33485dec74c2c36cb069b52ed31049c636a6a3450d4291;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17804b3659942547f4ad0921adca33112a9657bac76e209e56ea93fa2ef13eb06431acf138ed7176efd65edd1beeeea6be2099287061efec4dedd13b3c583faf85e47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he53d66a1e9a255464ff457ec280dc16826e1109c084eb79378e18220649fb8da7a877a6fddfc534424244fdddebd9d63bf7aaf3b8e166c1348ffead179559ca8f8ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f69c65eeb08cc1c74d1c4d9551aa1c913875a6057cb1652b0d5e2ae685ea0dd060aefa5266bd91e6feac43b1127f0407fd9b79e0ae19fef147214ec0a5237ba97f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16cad46fdf75a66b7ac427e257ff3f193247bea60c8dc8e276ef5427a5290fc364ee1850d232b9d3bc9fa8623ab187db2d7587a147bd71f171f996af163ef012afc9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19194c9b3e3917938adcc8d2ea65b427714834cbbaa7392c1880dedaeae7b7c8051709b1a9f139dbff9f9f8e0ae78882af97d27d964c454c0a02c7e5091d213f9653;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69d639ddc52f7320fe23233007f8434de168591c177904f6ae2de356999c5d34a522c354a2bf49c20bfb00c4628a4b97f7fdf003d0f75bff31c137368fafbac6b549;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c5eb98c52cd8b7103f439595595e5224c44a8b57c1fd24866c8f4d9d885b071fe7ced0eb3e32bef914661e895b395016003855a84ecdd13334101f8a786722f2eaf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3fd7fa02e1e1909e49cb2dd7f90257ebbda9636d1feb1f1f215641b22795362b1a2eae2fe0831b356d605598f1f065607107c18af3cda3f62a8ddcee3903fcee42f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a800415bf2292cfe3597221a7508a3e3dfe99f98b8741a8acb631fc57d51eb5a14fe4880d2b545c6a1fa3d8e802f1c915975696ac31dbeae6465586e87d0a12b212b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c726b4dfc9ed5a5277eb23af11e507f0ebc0a979a7ee8c8da1fe9a07ff7c62cf2865c3565dcfa4b0d7e208fa6426994c4deb43c46e6a00204989a42826f09ac748b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd2f58e070eda70361f4760f38487e55636202cd4055d8e5b34f33f69e902909535e2d6516a38f1200a147834d477dfd70236a60fe7056b2cab6b128a1be6f7af73a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d0ea9141709b9673be2bdfa2683d2bdf1efb2575e8427c1e06d64614ba4428ba53dc667820e1ab79797198ee05951ae7ec6d5b64fa5698f9054f9e9c92946c3d25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce475f7f580c0df2ec36758b4acae5fea18b9bfea16ccf1340cf3eb8de679b9b5048a05da052796f2e04a578d280eb9190e9a2305b8846323fe37c334d80d77056a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f26eae4846774aab6c5f290d17418dcf427b54a15ef5b807f9ab86d189ad5ebd5771e46a32c6bf83ad377ed7985fe2a6e8df25ca1e64660327c3bcbc64d35510865;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h156fa2e1ca76b940dbbf4f62127d36ee2f1c3ef698f82634cfeb7cde445aea2f44c05e6d509d7daa30a0bff6e3b1394620f8e64cc81ddaa83f2368a1ad0f858edf368;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc871800cb9f577c5d76d5c2218ada42c0263e9ac63b7eb4c9c3f166da870ef60a95718d6c2f263ddf20a53b7cf36ed6188795b4e6ee7450d112c9123269f6c81cdff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9e40732b540e1943f0220e02178d5d36d6d4bd7c91e766279cbe232f4423ac9a860bb1003027ada15030b081e36c17dc93420c8bcfbedd9560733d91ff6b0b8b7f2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f17e36e25ca04d8a5996080db1ef393e4b416978b68df364cd22e3b9df2636dfe666d2984a3e5bf370fe900ecfc4de109dd5943767f0b1370e21e293f9bb888fd7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10aac2e783d1a7fe26ec073ac789c640579e540722082b6bbc18017d297561a59f5d034c425369d8c85e9dfe459ba88aa783051250d7b3523a580e1423426c80bd56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15458e8698bb9c69824d40e79a08b052780314a5182edc2274c6b7ceaf6f50dac08200799d127c5792a8c536f1607131d2c63de6f2eb56d6509aed620636295cc2228;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a8cba828da0cb034ea0fa9c324dc98e3264093fb16be3473bfa76dcd104c571e0167349206a7db854d229a92f820c0b0c3f9748c6d64ae6238a51c6cb43d8d9804d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ccf798a0ce2ddc9cc80968c80a98e05ae9f393247643aaac5e11e0ab0c33e3854be50887441c54c4ba28f348663b13db838b1a071e9faa6cd66f74faae2539b487c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h445dd5a9fe89a8846f59972a476531a7e47be68ef696c8656fabcaebdd0d3c838585b96a72616be8d6f6e4ec68348aba408aa1a9eb22fbec45e11c9e28ff0cdf0d50;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74820b4e8cecc8be75cf0f588ef7a1ba16ed8f923d4f3ca5966401a427a8ae5cbd87b6d4cdd624f2ee18dad730d129e7d02124bc2ff1fa6167b864b882d9a58e5f72;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc3a534a3bbeaae85039bafa91ba8144eaf74eb75b090181d21fa27e705ad07518cd4db5034aa078e5e350a55d9714611b94999aae6d81dfdcc0a8208034b45ed538f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ac5a6e84b7c66f4a388d0387daa77718fcdc4f180271125fcd9f24d4bf832706843f4dc7d8462101342b564db582e658722abb1352503f11e9050e4bfa7abe1dad3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1073bada351578230cf349eec105529c3187da5cbe82f7b51f6a7eefb2cdbfc023674ddd23b0fd35c3e931bb8d49fc8930bd8e7542c8d9215f5e1783c7591268604d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h493f01fd96b7baa85604d7a152a587760aa27f3f8024bbf967b82da42f8beeb5009f31cba863cd36aa2994684c0cc65f811f8a107e00eee882ee8edba74dcb34cdec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c6908e6d0b64fffe1e4298829450cdb9260b79a7090915527bf61fb256d873364b36599ba0ddc7e61ab337dfee99690e852e0a3e1ef9c6dd4ced1317a5c4673a737;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc6e03fc63dd041fb02f66dff44583829791e114df48eada5b07c2e13f0f1cbe9e28617068c3b582bccf0fa7c08a80e02bd4f5cb824585e72ec74207a46ec598ee20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5efdadd3c7a35a1caea8b8ccbbd6ab361901bedcc66fdad86fe965d8a69be275df4465b1d8d015a1ddc4052f21eba0c6ec7c09fc35e91354b533e2e1210fd41d9617;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9c71a14fe976c50ee96fa9a122f84a123f1fa675c8ab454490489c52a29526d54ca5e28e5cc01cdbfad3b20f7112a7cfeeb22bbe72fa741e61d45a42defced75f16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he1b6dfb8bc810385ee24d8db52bf186ee5c0b10c10ea4e1e08c9650838839f02279a5a3f6ad7ca72c3165756b07e76fded57d501f7b1693e50a0ffcc1bd3fe7ca0e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2bd996f5e4dda91fb1cbe54d548919cefba81972e923c4bc181d80aac3085ee17792d49db33436f95ade13ccfe128aaae5e1e9b99b9ffbb8d846d4faad64c926ca42;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf3d6f7b971d660b6de771d1d3a1ca02f09f48601e81659da84466beaf1e70b3e80b267ffe62cf7319c3c840dafa4ffd3a4c37b88ea2deff4eaedbcb48753113d077;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf1bd9532cb6f1f385fb641867cc6c1d45e307584e87d18f5b720d0b8792d2b52f6eeb50803fda7b1ddcca54e168f808e45e5e51c96458ddaca6da60331f13e28a5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53dd7ecc8d0a9e12e6889d90f4573a5a25e422fb588ef19997315bc36382780e674758310bb9e67b5f82c51fa03dd691bd6779eb734733286fa21104b27068574945;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e6eec4b22b7f8a1b0177dfc90f3e54dbea545bb18af562a86f3135afad7edc587c561901a17535e8cfe3c89e65aeea83e28332cde7d0b9bfa6f64334dd5222fa98d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h81dbda5ac3a142cd0560544f26a774f66937f540a66a8f474eaae0282429e9da8fa24f261769124f03bbbbde45e2ea88611ccc4c347711513127330c1aa2b8a27428;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfd0e8a42510ecfa8150c9116aae36bf388edd9edc89cdf0642550a5dc3cd2c7658a828000c888ad3f5feaeed0760bac15581ef988a3b1c8727d02af52220e62b2d79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ee094cf99f1fd59953179f0dd9ae58a71ccee7f83d8e27bcb1e8f22a87ab3777512ad7c0e0da3c942aff1f64c2bd19906668b0fa4809e13a13075e737454aaaac38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3b2f0fceeed378ee3c826f137a5367e31af6b341bf3cfa883db5bfc7b7e6aa6c671b2e1e00983be5c545a5db8f1c6362e8fefefd7733d5e210ff935cd389fd9fc080;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e3b2cf9ba1148928e5274a62978a66d2dfd2fd8d91ef6d791c102b8c37ecba08620544ceb514710712118ee674e8c6ebf9bbe6c8ff76a700017cca0b776822424862;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c8bf925f418a0880e2f4467f4199545732ad7cc41231fb42591ee476a6d5e09965a4d08c880b0173f38c30d693e7f09e1f295b14be67353ce64e7447ea0a9e62e35b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h944d462716d14ccfce8d4c9a6e65535e65beafb04625a1e91e8a00aafc2a4666313d5742141ef459da202951d87adeecdb3dc79c40601a7f8d43a11c59f9b114e57f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd016010c2a36402b387c648f5e740786d0ccbb0e2820def4085a96fc88a91402504274a773c31bfffad810381bd6e8bbcf7caf189676c6378849a70d680f52de801a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bb35499a42781107260c0d34dffe0046a3fe00921dc27b3a6fc1cbc425587999a7264e60f1e07ce5bca38d1cd0fcacf7f181fe937d3f209f010676a63474302d5173;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h835edbfe14f28afa1c63f0e7267dd20b9d6814de9e0b5683894a3e58f764235e9a74823e971ef26e5b3ae4d05f761aa2fd5296dce067ca2a24fc12ab9461ea02c887;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3305f34e52ba918316ac2c358e596710d68f8dc4e1a8852b0c09278b5451ad0174ceef358dbd2122461cae9c76f465b925e853e4f2cf34ba633cb28d7bbdeffee40b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f642a11df21ad4e6295ba4cc306c809eafb43015f34d18181cabc85d0c7637a572ce9581b9f12af9bdc40d86f134379638b17647521a245ecff6b3a55d5a5e25b5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89917b109a81605577f84777a96ed1cc659e4592beade0bb6de67334d05ae949302f1e5e74db89e60162f194e7ee8bb238b2adc107eaad9e2305ef4d2b557b316298;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4728d320755369b3da4e82c3644c44f68a66236087af74da444dd412b2e3b6b29c0984b40888e2dc09ca38015a4ce62b88d9743af377f7c79da34c5ac6caacaf2e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h151a38396e38268c012cce67376e6dd2eaaef1b7904d82a1305c80b06eeb30b976d5c9a229c1406a90d4c83056e64e5065b01a614a32352b56f74ca6b3004e849325d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ed73ca5032e59abb75dd12c7b35368397063a4858d63d82c21b4479064d7446c0ffc843a5259d95627e4fe9a0abe18ae018a59f9e42106bfbd224792c8505a4c6664;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f62e4a3f59df219ba201757d684cd9e07856d6376bd9aa6883e4cc96eeb24046fdd9827797e6fbb465c4cc78799d6b8dc026573f3ad8a721818a8437bf589217626;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h291a6591e565b10523054a770a30b872e95c96edf029a8816a4cffa6b86be2339fbb679e84a4ce0cbd8a74e834cae9e101a21b7269be88d95404c348012ece6a8795;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he00e47fff91c0b5e60c041cd26d71cf49ad52cf4d3212e8ef8246bccb89eea9f3a7668ef01bd41b92bab6d78fa79c39dddcdb67f2601d07cd11c909d3cbbfb9ae686;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e77635cf4e4348c356c61315008ba22a72740115ed50a795971e535975d0f8d40d4ddc280177b09837d2acd252b3f27462d3b0d675b796ae0f3a28143090b776eb7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7bb842ed48e1433860220ac9064bb6567e27b8a8824af0d4c323548725de5c60619d34dd81dc97d7ebe0620ffe3983e5b948ecf44117f48777e47554e4580ff1f299;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1739937a0ba02227f5739c3db5d5df32a23bc15819741caaeea441deda097c24e8ca11e62961656b39780c0820390b2e4e4c891255ea57bb3c59362ced031447e8320;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e113861cdd44a8fee9951e698fd2bfa30ac4ff63941d3fcacc3bc886dd67aaa83842c7e8abac9d1f06a99af69c986ae20646371e57ddf8ccb6e00e70b5d170236e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha45a494025b090d573879677fcaefe6d73d008d064a2929bd158bd3a286e297702bb0196f56a08e75b8096d4686fdbe1442e2d8bc81bf28775af1a0a265c3ec00e82;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc8f249c7237ace3665f616b93f33c72170a48fd83d38984f97df97979d5e410b842bd13a5dcf0f161218130387047d66079861b2732cff2ec12938fe0616db4adaec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b54fa272c537db3157bca6a327a17495ea9aa2896be24ec24fcfe07658844e32261c87b7b99346641451af4825dcf1deb560733c4f4bd6c2e7685306afaa2cf6aba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38bef2e575a7c86452e0e95655ae6b67ad5a0dd991e3bddb5cbca58b1ece98d6974776f11ed9f96e55e209a09afea4a2ec8c7251251eaa9f89ca3e184241cec373ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b7a8aa28dc539ef5ba4f4129cd82b9c4ffd3fbaadfcec0bfe2933684fa6528f2afedbfa29c3f3b98d4a79bc68c4648ab914ed5419038032d1ddfec9464d973b1538;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9f17c45c6a5c1c4e110f9ee33d253b3bf0e298ee40e621ab9b91a0ab5f2edcd47817aa2eeebec5b855463c06ca0eaf23aefa204abc65999085d59926bbfaace8769;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h87c26ce6fac5409699a7af5ecb90555c7583e1f1559ba9fdf6a879ae5749d0c47fa843c74f9ca101fb10faff9485db47af295114adbb6f86b8c7580219ebad8ee469;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15dea6e8965ed792150598f3c67bc2d102503730d533a4e27be370b8ec06d606da1141b2b6446840a682601c08d1ccf8fd28f1445400027bee6bc23d73ebce265f431;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9297bb4ecb85338bfe53fd068577ee2ed45a12cef5f5662eb8337842334a1bc1ceba63b415a71e237380a5209dec1b1c87ce30beb7c2542cb1b5539527afefd8087;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h81ec1f62a54afe4b5f5b2b5042f39b894bc08f0656b975f6f70067246a6feb6e9eb43bc37b7dc75fb10d67cc2ade3eb55b1a71c8d755ea2cecb5cc0c946a9ec9484c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b939a2adf03e52e599cc0ec9bd6b3d6774e97a70edb7465a21d87d17ca558d090464a3718e5529398c5caf914d1a43499465de5d5e7899cdd6282026e4a1c620b0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f7b1822c064d389bf9b28069e98a62ddeba01dea84366dec5570bb544bf386cf4327bd481edf2942be681a5fdc744e14af5865d220b451d7efb3e767b429dd906c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16b0fcfda284e9000ca930b7ffcc11c7946a3c443986f71eba2e7638a4e47a0fab448a59b6cc0efb0b91666ac749f9b49b93f4c0cee4f49c6b6184b7cac87e7560f8f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4bd365613aded422de4c29cfe1496cff6ca28e47bb60fe2ceeb3e38fbb27277fa6c8b59ac1bef07a48d8311fb56f734a0299689844d82bcdf1acc2fcfe68e7de877e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c2eb878446a150068f4425e89221d27084d4e7af243cf606e0e2a7412f400726090a52f1d212c62258c67b4908a973e93e95649ef7b229b82f50fee6e9b3c0dec08;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2a27740bfe1be8f46958c4ed1cb416a3a1421b00282009643f499449190b72d9924de49bd43a556127e063d6965743a6e39eda54ec843fef8245b112ac0ff903b609;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f6292602babbc07933ab9ad134df77a7fa215a5134ec9ca1600ef335a492bca73a7ba431833cbf7157d86df5a48062bbdb35c79d3b888b0845d3560d61892cb3a46;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4842977f1f88a30967d20580f11bcb1203d58a2d4dcb4ba09a531e16a659adb81334f01e87a11b99a689972eae2d64d8786d121e52996aa9ae4b02cb2d2fc09d1109;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1770cda9a1427e3c42a0e6781c622b9af7203848c421dfae49369a1d7156e7367d9fd55134c38340ce58f61c34f673abc7ca3b7807dbc8f64b8c71367af38a92687c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a00adab9a7bb5b6604f0602ce4b8733fa822bb956c47e87621492ecf25929a2956de4f437f3e40d648e197f407a92194236bfaddbd77cced0460f151a2b00c65e14f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6ce856bca0fb666c5e1ce9d891401f7d938eec8129fe8fa25872c50bfbac860a6137de9cdb48c51675679b8e718114cf2b3f2efd478eb23fe081fb1f0f5a99db64e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ae44c6c4d470aaec291a0d5a4c31738d7b625e40380e40a8fa13e565beac5b2aeeaa570f5d075d5d1f645af119f8c6d0e4c3d89ef9295bb51374ae9f8bddfdee504;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa784967449ad2eb73456d180ca395796b188f9aee502e2bddc46c55861c417b9c43f5f64e2dc5d5857442453f18ff6c54c17707a6b278debc22ec68109fb30ee54;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha76a71842ae059f2a75a36ac36505616849ee8f78be23c57aa4b24ac0ba62363acc91f9664ec9e9eabf896b4d331f207dba4d1a68deae5b253fa225cd743366ad41c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h176c260cb18656b7a8348c10d9480d62e75e9879f1cd14221d70e80e980f8eefbd350fa9a2a2908b8b17385c26b35a2f2ed2da16a335e72c838e08ef5c8e581678335;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h78a5007e37d2546fecb50cdfe7e5f22db34aaf0a0d5eff144e53f16ecc6ec81b1393a484a13a02188a86c5ab4d4ce20bdc3c1e94e3943c60788b7187eaa738a44ff6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9277118040b45ad7e491a4e4086cad0dc5ffafc6dc8232712f4b248778c16ec5e22484be786efbee13a549a1ab04c3f92f6f6c1cde4d9354366de5850ce636e60abb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf91aca8d1d51cfe499f0ae9520191ea4f6cf0047d4ef8cd318a4284ba4e247adbf119d8d224a0e110a2ffbabe505d0bb8093d2643ac8365d5db19fa9374c14812fab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1590d5694653f99a98fcc3858f7dbf25f8663a9b647daff4fc538473a855f1dc26a1d1d418d8bdae81b239b673a1c29f16f97ea76e9cf4b495c709bd5b448e7cfbed4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7738f8e7c012407850c15237ad5a2bc77c4848a3ede4bbfb7f940abe52e192d06b89a329fba85c7faf84db23e58b848feacd79578d8b584a099ca951facd6e02692b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7fd234e3ea7035912d7c8c14ccb3e28f7fb9c3ab7af9a2c2dbf36c26c82f132a1e2ca7297c851caf58f779ad40f62fead07477c1750df2f8c2d5ada8c21047a1ee9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dc528a7e1a7e0c07e27c6cc35bc09d88c4ac3ac8493cc77a81c7e358687205a1d03b3bcf02ba3f3a76c6b1f1ed8f96b9fff71806bd850c97f45d9e9579dd9384b163;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcaedf15868d81c85a10db0c2d51b27a280972000bb2420d43571c0caa05cf7dae0f9562784ba5521a3ea93c3b8a511af3e1d90f583cc891687b16a781828953b9aaa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74555dac48df9e4576b60fa7a754f8db9433bd13b2ebdee589d318ea6c501aff7590d8f6b46fe338f414c0dd6a3f6061c996dc3f17a805e559bc0a9af2cf2103779a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ee8645f7164f32b1abbf9ff09d8c99dd047443514b3e4bdec2df337d1bdb4fb645c24253d1422691c53bdaa91fcc9febf3d8249e0edc99a1e2b480026fbf2b56a66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h124890d2dd11a8e5d462b8a01e389b03de01c4a79f2387c31adc821ba227769b6bf0eb9339af76d925cf460f4ba52723969f4e149fd5ed9bfe66e6ec98c1325cb68d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had8c0675ad0a1b1f56842b948831b5d18d5d7267379ac877ebfdcd819d9091445c3230ee0f32544d3bb548b6f3b60d75f4a0fac0f98224859896ccf1fc3ffd332901;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he11331d4ec09674c359d5e585daf9ae6e47f0c42fb1b5cfad9e4b88264c30f8a235e5c98c8542bc23a27b30485e269709a7d7e49d81ffcc6b6040ab1c3c22ee48085;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4eabb14286f7e9d7b08a1e675086a808c12a19caab07679aa4b90d78f10cd393f92c6be71c9f01f4f732c6f40dcadaa54dd457768777df8b1dd77a3d25a60a2722ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67dd84af96714ead33cc183496d5bebdc8169504e826027c0f98e9672c0c914b8ee829d89282a25e9029b4577cd79357e69bdc5d1b7561687ef28f2163dd6cbd3fd9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d027fc1c4a212a454fac7eb5ec2b6e938f9350e1325cd11111c3de3c0da1203cbc5afef5cde310af82e2e791b217acd2aa9bdcd560206b518a31e9c4138a2ed6043;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf34dfc9a451e8d26954a7190dd89de818414f362ed460226db0ce222a212b0dfe1034c21093e54152df186636f94c9a28c4a6cd183d28f513d933b974c1ae8dc89c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12315f9f5cc624c7549e7783c1518bc2c1db655cf49f42c3077dddc2cb0290e40098f5f069e0553ce7b4e17aa6f8eb9896e59f26181d1fdf955aede9f48ef01b434f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he628d4f3680db47a19ffa359f83fb401a20ac03b8c6a6bcb6cff1d22db7a8a02776ddc5e6c600c53ec5d1bfb6e59c2e5965e961960e10217693c6cc1d3f6cdc99d1a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129660c832d270ac99f978cd5fafab08841361877785f142b58da26bb3ae7b0305718eb1866640a7402ddfaf40c4f3dbbf4f35933a6ee72bd86c59d758cf36f99c942;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a810ac6f133b932ec27f8debf68690771bc3f8f2ea447f899458e4410053c0597899a7d76f37687046d24444aa59eaee058bf99458d9d8b84ffd855a9a4669b44cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e377e3fec3562e21ce60abe885ea757914a7939b1b0b5ee2de81198faaaeb0b313d62bdc50f3dab945d0f23385282ba6240962cbf9b997ee81b0173b102d2922033e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1943eab222247f9cada7b57dcc903b539a0f901e6a3fcbf36da6bcf681272e6e47f00b12af0c05a3455e1ba11097e4a9bcdf040e1866c911590b54e71aef020049f10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1282ff8a81b661e202c61c90f40ffa6c6aa646a49662989b6bebbab047a48c1ce3f1d9f5a791557a6efd144495200b9342cfb63783895333cbe254d847c0c6a3d7e07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcca87d5f59723426b7fd3435fe384a7723b4721dad1a051c350fcf65f4c2253fcfeaa954829e16960060c9441e14e40abf2404fbb5f02aefb659fc49eba7123fb0a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73ea85316fdd6344f93147a487b0071e20ead39f1d727c8d3891e474b1ca2bfb404897c5d1020c1aca051a8a46ee5a5a5930c41628c11adda32ff8f42813ee34816c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121486c9ba2a6616b15d0f854bbdad814601300cdc25b720ec0fc7e862e28fc572984d4a9b377d348c62c6e289cf5022282d0f530b4cff83acf4da6fdcb0901a1660c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b0b14959a30bcc33a8216d47cb12dfa7482349d48365cd9adf6d07ab1636c5f9114bfc6667469b2f17f9c3cd23efb96ae06eee5133b435baddd0093a18c46fb4cb5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hee59dafe1335874d87bab31dcbe132c3eaf3825c525ed1fa7fdf0b06e80dd38d4abe192fd2b4920c148aa281688568a7a6097c29599f1d475c009f7f3d3277d01a2b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e8f2917513d4acadb06d177cfe33ad506e85893bbe11fa5a3c930a10d60aff7e4a7c5127763bf945884b2c00b3959dee1b67a68ec1fe0c567c5238798707ee495692;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h967191779aaf06f81553c935e19be2981082ad9363b98f082a1727331829e7d643b3f2437f33264c71bb0e57fdbf2fc970fca86da1a3d9813a6d4d2af4fe9cef0427;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h35b0793f54c622481d5e7f51be5f8f472a62d78d6c785d981d37bd6e08ce1aeed5dec2f8704b9b8feef584fec45bcffba1d7ebae0d7ffbc451e8492ace05dbed3aa8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ed9c6845009c6ca6bc83b850aae5e6b67223edfc95f745fc67c18ca8b403dd07482b920f48b226a8b52b26fe15f96566ed668d16f5b685c15e6e4b0c15387eed1b3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2066e65197313ed99549d2ca8f21a38d557066864c5a246d41a51a8ee63eb0170fda8948f1db69fdc03f627ff62c50860091143d429ad108ad4ace8f940b3c8211c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd0e634cbc21029e9fa96b4b3e287390e6e49793d24d80dbcae126f4b01d4646b9af4f089e880e571d65eacf4731669f15775d1bb4ef750bf2814916b5eb7bbd1c1d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a71d3adaba17f097fd0cfa949d6767e8d0a1cc7f291e8b1d9d8c63556fd90ce27ce96e80586df0be55e0b7f79919704b3412e63139b8ff9e84c11a74619a03bfe51;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbb6bd86f3a4adfac938738b50927edb822d38e8f9b6bd04d2ce1deea7d0596c8b27999f70a75b67446bc03a8b6ba7d48c2e4c5867fd146ab292edd01f6a1f200080c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d152db2df90606b568f4a687f3b5fc3f6dc81b15d1f8f87279447a1d1371ee56474920d37fe812de91a62bb8697c73cc882b325c1029548040e2adf6c888ca4ecc59;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ebbada5cdb393e4ca6396f56ab62e037aa4b6786df94db106539b259c9354161f831652c0c64de2e9200ffda98d80c45b5af75d3f5333100452ca25a9ac8b2cc395;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9b7606ce471c8764c02b39aba160daf062912f0ef8b793dc773954db702c3759b150e0f0060f99818ed33320282b245e99728377dac67b53c542cee2f940fdf6ac2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf78013fc69cebacb20f07746dfa57f59578e312b2126ef9196dd209f060b85ec2eef5cdd7093e15211658198cc0ec4f455d13d62e8b8c5c4ad1767329cd422f37c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd12657d3bd4b8242805c4c9537d6beaa375c60b76a5211f1d1644d102964dc484701a8834d802366714ecab1215a6f2d6cecbeb84486e62cbf0f2a00cb5d5fdf79fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12ad44bdca1b47574e62d9c26cedf21a2c622d2b0a7c54e19e6d03905fd520ea24f65a7d6fb2a47fecda540ae5fe1a0d184d5583baddd22baabf3648ab2682058a7a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15904677b5d9f639a0126fdf1f66c59bd59287cad51a635063568d137aaf786f84180372aeed129cae3fdedc31b19cf452cabdc11c7c737e17e475f1b5919bf795b96;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1502e01034870891305194454bf2b863c99045d36b065980006058037663a314db975cc79755ff3e24d089a06f5a61dab19c9d199308550dd79290712971b232fab7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h68f70754a565581db1da82491aaeff837eff2540d2542757ce2738e1bea81eec1aaa317c2822bf83344d8848094a450519d6346b77c06a2bbfbbce91620cac4ed92;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc5ab321835a7c8f399763e612ad0734ad0921c6ac0f1ca0e8b980baf17cc061e79a88a56f019ccd1fb10443c95b19de00d7837ac90060cdc554ca34a0f74aa73c35a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a56e6576e6cc46d288c281eb3cd288030bd42309dfa414290691593608b3060b359306a52a4ff38a969bf8c82f9214b1c5f2222708199f0acb83328aa1e2ec6731a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12aafc50f42e4b6f7b76c4775ce9e5f1910b38400367d4f1cf0d44db1f44254387d9640b35a80896f0810058e57fcba88e410d5413b4315b94dd076fef7ef7af89d5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd0929e2d723de36f55bbe17005ca9138b44ddc821455eb296a1b468da02c3c16a2598cbac4f65814c3bf955d195b9d471bcc2486b6e9a470f2d668855704a7af1a7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cb03e27b4aa27947ccfdcf670551fbf47e5af944b4529d656720d549b773a3ff6f6a487e326ec990403f80884c205c0287aa701e515dd17581c744fbb7c34910425c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d3e68f7ad2a366e54179136f9ceea38b29d3c65898e79a934ea45ee3e1bb8d4e6694a4f6527f9a52e786c09dcaa265cf99dfa9de09e0afaf8b386328110f5ed03cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h169e1ad779d2cc179c854e62904acbba68d46d50e967eebb3afdbb53f35c43579e708ef2c66a9f9d408e0eb038451cfc01323a0b0d7b473bfb1a40d670e65ded6c6df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19991564e7cdc54b6e3792c33fb6567977b218405a8460fbdb80f65666dcb4b37978e190537a9fcbc975f579564ae7ad77786b11336ae48f6b2b2ed124ac80e74f176;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1156b007c797ae7282e8d99a84305b609edcb96f609a47d27c44b15c752de2f71cb41d6000fb02aa4c82c5122e8e7601219ae8de5b2b1da90b20e09a9e49c4fe1ca29;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d621bb57df5341fe4cddbfb1727730557ce1d67391b1ece4d1459ad9922a0f7f8c277e5285345e3092ce6219f4badd43189182586d973a8d4f3c769ee383e6f9c7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ae9496a91895247e91bf37ed8f2fe6e3b8e423edbfb93bd37143ed0f5c3eec851aed6eba501f2f0352dd97f34b802301e609820032fbb3798596869151bd8053352;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14b7724583fe10c90c53872c527d8cd1978eed5d1dff7872509cb061274a17a4b1d83f8e142ce5a0c140b98160370a2403c9f8889b4c2adb04d5860ae03893b433a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d0045ca5369ce1b318a50312f4f29a10f00c1722b204cbc3f2eb86d8b17b76c792d08c950604432d95600fea1ae6000c54676d1eff994338df688262ad1e7f082788;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8539cd6a1b29c154380587a5e55161482b59568e5b659876c121676567f63fc2177a9fb34efdb9c43c86655f04ed89791a901e21d9ada58d7f2b0e7ffc9395ddc7e7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea93ac18934f9a21c6f1098693f3a2c8f873ef444b1d66b1b58fa958c56b75011186be7df3b3c56761bf94f4de1d23348ae836cba65763cd21e1fbc2bd2c7dd5068f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h879d0b869dea873108327d3a4169cc8195bd22099a48c80eae023a7aef756aa6d33bafa62cf2d4d51e3e71e9bcddcd2813904a491668686e93160f505490f909dbf0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66d580374bb665e35a468c2fdd336faba0c5ef1d3bd6839bba22fac25b948370817a8eab9ac9672172e100cd04384ee6b35b768a8caf0c37d7f7256f82f1832b8bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1330c1e4e6df608313e6657f42c38e644554be0dfa88f3e80c130da06a08077fae7b09d0d160403437d8ce61f6051024f7f90c473a75848e617ee1f7815b5103716d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc7446bd0770d8f302f584f35196287af9261d2ca0a5dcbd945a83780f83516de289ad8ce5727ca9d422aea7b51d23fbe07919c8403645de34d265805245f850d2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f9efab6546e24e8c61548282cfd493883994f679a7c2489d651227a6a45a5d949d5dd3c6bcbc861eb870e128111b29fbf585071f85fcab1060777d89e908f8aaaa0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7731a8518de9b5fc5891b9c0872651686c0265a79be783b8879b12495802fc57cb08ef3c9f74f97c3d070ed8dcb6bd20e2247838e990dd8c1af05382c128d44a634;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h183a50f1378285f7cb7f2d190be092e2126a3f6e6635de28c02fc7ed3fff6b7b8cf4f11f2688608a5fb5305ae4eeed339c5a49509fa870012934de9904664a8da8b1d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13cb2c496126788448dfe7acf09eb31cdb24e79f17ec04bc83c68b66f4ff3d8058bcb109ee2c7fb28986d9b4a81e0a235c594b2db5c84a6f997323bd20b11ad5172dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h280706da7adf211a61ea041dbd46a5a86d57fcf8f02f29288287697965b94cdcf1cd8fed10d6432a7946abeaff88adcfec38090930b85e369746f4dfbf389c1e7e77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h192bb0c6446cf5e546391b6241a456e041a62114d5b70189ae79398d920c969bcb092dc7abb4b2e841c54d6fe44bbfc3ceb8e286aacb33008708d7d8e8694e43e9209;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h52d7e78e3be7d68b0da74feab45293ab2edd0d2a5449d9dafc014cfadbd9da09fa4d8a66fd29bd8c3eb1d21445ece3fa2835da798b20f9676556880ad83e2cf68a6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heed01d36ee2472e060cebcd3afc795c12c51d236ffdf658ff1c6316d534221a681bc74266b03e3e69ad66ad064540f0cbc3d86707b013753032d991ea644d131fd61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d594f3d4050b97cc59714d72b907409de6c2f5c757e58d515769a498799e4aec2ffc96812e426939f108b4a733c8d81ef16b8291c7de5ed94ff3da51982b22ffdfe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5da42a3fd8bef2afb5709e6795b35154a55f463a18c66f90f25855b00efc13c4b502ff121fc150fb04b2e40dee631fecbb018d2e1aaac5d7751cd86023e91d177004;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h100f10ea5dc7569b5f3bb9ba86ec614c7d51c1e5bb4ff87bb01d041840ef42348d1c12e2b444cd5079762cfa81d40a5eb9c3faf5431162b8f97090e513cfd33259879;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha63439ab4bce5e62aa963f6957a8a313c23f45d629f1a65b690dd660c093a0a3c99a6decc3f047bbae1d5070de5ae63f2e5c69ce60c84f0455dd3eaeaa040f95c924;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ab1c7e83d94920eed3fd029499821a308352de3d2145e992260639e43fe4eac7f0cc0c7b2d3a9caf8312fadf4a658cb868c2174226fe7997c2bd1ffa08ad5e03b9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haf8a1e2881d5441b81ade90f71d2440935332359bba24227d65fc78469b5a4ff3c0506f6d2d44df7b03508b6b19c66b5135e79c1315b0edd826555481fb7585b23c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea74767d018f1a4071f646c8e905b4ef8f6160496cc814ac73b31fa71898f808d42f1d9c5efaf1b3d4cb6ceb95f0cdee31be1daacd4588ca3a70a0762d44ea172b08;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1263080521d8bda444299b4737d852399fd3e2245a566397342da9f107241e37c6583d7e8d90b2af4d09572dd69993717a08b39602a073724948fec041f795406fa5b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e4d44bade5f1edc6e725511aa35836013d2561d877ef72218c5ae8c6f59a0350e73c6582e29f340afe2fc24691c850f546638bdb752c5acc00610a1622e2587df8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h683154b6da2d12c02f4e882c1fa5ca7dd2fdc2a48990c33dc48b0ea9a4f47ce16d42f27ffd8ec08c93cabae9265bc9818e08c4380977fbb912230899608d3d388d69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heeee811adf45a2a4c6701ced5dd2935faad17a40bcf385de88ada82d1694ec293d64b3119f0f78fd13adfe3dc84068ddbc5355dd77924efbb67f0f2f87484fec1bdc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149c224f4d6a4e0defb7b3d52bdce9fd1baaec1b5ca17fae00279e678304b8e9e7ba1af86bbaa5ee365049d76cb3065ed1f970a4e0194846f15ceb25bfa4724e8da10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2f06e4f173e99d3a38082d4f033ed28b8d38727712143138828e89a2124e10a0ba86297de2dcdf8a8bfe58314d4a0e86d94c4881be345604966c8f0927b74135785f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2df346e0afc05e239d718d0b8cbec1087becbd883cd4d66e74256bf7926348afa86e598bacb1b2f29762c79ccb1828ca95252850334c202a18404f1e1cd8b9845e02;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h122fd561fc96d00b8fb36ad83b70b96f1b3e43b4a5909700a1c029339d5b9b73c85b3f8836e195a24920eb6629eaeba7f8e85ffe897a45d13bafd665a0c949b7bec65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4826e4e1d4a66666aa8ca6c51b040f35581c6f8516f475df8b59fa803079bb4d4fc74285698e9755ca0d2c2474e43bc2beb209ef9b8c7ac21d112e57f051a3901ce9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1876a50dfbcafb447bc8c84658c33c6248bc8118e28383d46f4dd2faca616d192fa7072ea34c69db662be0cd7465f2aa8d807859fb5562f3933be894e994398588295;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ae29f1cdb7e1873a5a9c25cbe819e06ea810453db2e3b2f2d852a44330fe4b160b383af0bae6844311789a04813b561f35b9705e27e8e7d508d444ef7a1c575255b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h122ee992e8caa5fa885a1ca8c134cc7123f925d2f60624cf510671c5e4810a7a807f595b1d0702a134aece6ea00a5171b5b558e06ed08efb8b6563babb2e3bc2b30ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heebeee8388b214a04872d1d018aec7ffd89451a4eb1d25455352d91c0bb86445540e60db5cdaf0f1a9f0e20e39f18223b6ab1b0492bd5dc07c6fa5cb595952827fc1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b9e50ac15ff186f625eeb48b4757426558080a230db34431f9d001c4b83ee71dd11a8f1e3219372e0a3c169f0d795e7bb3c67ae06319518b9805b7da6bc587f98a49;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ba38de025670c5ad0a39cf7b9341013736abcc6594ab9f1c48874437c9ae8a7241c76b33ef8ae6a10692a2e19e303ad148d6226a3e71e8be915c8a10e3be4a2025f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4ee628b0cceba20f00e38b6fb08fe3d5138aaf43ac03749fb0b6de0b96937140ac1ae3bfab975990975f594f1a6adccf02343a354053cc384324feda53944a62125b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b33654d0b3bb4986a91d81dde1fccf335e28e0fd9d99c081cc30a7dc42a8200ef044acffc8929b517812c128fd2ea97470f79028f77c69cddc8520e12f3ca44ae04;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb6bd2a3e7878caad0ce267d368cfa356aab30e54ad678e772e5a3bd5ae6363de93e245178eaea4c59e0a2c8470a3e2ce65e3494a95a4620e3d9a7489301ae86c7a38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120b6f62de3ed1ecd8d5aa29dcbb87bf534ab76de4b6469c050defe0541d78b1a3cd892866d1b72fd2fe0f8e1d78435163ea617e9635cf03a34ed4d1db11d89d492a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e60542e9dd8ec2565a6de8384b907a4a20ac8078d3cd097e3abc570d0f3dca2152629836100dc191824636cb5c1bc31069bb9141fc866eca2475ffe4d2498dbc0abe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc013f9887bf8cb0db42f80edcaf235a4fbd834f06823abbd5ef562a4220cf6278558487397f684b2f8ddb1f62ffae1fcff8d0b40cbbcb060de6121081c1d33cdb8d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1053ab7bb6e48fb1dce4ceb97b99768bcbd6a28510fa16ddfb932e21594e90a4f2f289dc019e9a7b7a2589fac6833c9acc0e3054b4ef1cb4fa6ebf638a1eca86992ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e43601066a49890455b352aef511523c56829b01585963ecf993e33bf5cec16304d55addcc00b99786a0480881a26cf46efc399caf6f344370a1364df7112bc7528;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b9a0ecf8f7bcb360f07a423b182da4c1408bfaff4a820f04f54c09efed6a5ce58eaade8993abee381c0ab8248439c1bb3f1de91c7683835bd7751ebabea6823df80f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1637e37e4b6c895e6066c4c32dcaaff8dc6ebf2e34b08e238dae314c787f02a8e2db45d2a752d76582d3c8fb3e8516e604e80fedeafc14332826fc84200da6e6558ab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc8c486ef3a844f4da54a58d71f359396fce07f47a5b1088c56bca7feaa7045cffcaffebaf813fbdc17a591e29d3f5fde2c4fde2d3dd887e61576d1bcadd805e0692b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38b23e3eb3ea1e10ea4dc8a9b50231a3810add1e3070e008b2f51f67e6b4fafd04b887f2efd5941e6ec99cc1712c23440144bed6e376f2e65b9c559be0b5259f0c8f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba9644ebdf2937edfdfbcd0129fc7ed4c4f135620ac8f2ca3cd01d89cf4bd049d428587dacce8cf85a54d4c1fdcd2ac6c58281660044754bd541f42f06495a98871d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc73d963acaccde049fde3f083637a9a05c6816722719d305dc763c1cf2a937c1c4ba31ffd927ab861b89e8cc1ee1f2942349d7e32b91b66dedf464158af3a61d3b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h155b9f1ae1456dba1d3b9a4804b62cb33513f041c56966d5eb4ced8d1f47c6c0cd14c36de63f0cce64d1727ff503bff9a210f085f12b23c307dcbab778c8af448b95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1faeb6a53442537e5e30484644fac8657864873bce43221a05487de158155ffcd6b5137035ae313974c62a6b9f9beda396ed5ce8a316319bff1cd43b76d54103ef2c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18e5a8771585ebcf39ac460664aeb80e72e0258fd186a44301278af739d658b1541b56b1c1200d7bd94eabfe43aec041548b158d68e47a938c413b77f085dd2cfec12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10bd10a5fbcfaccb38bbbe7b3c3e57a69bd467aa4fd49e7ac267c862c597b28f467cbb531bd98ffc26a955f25e3c4cfbacf1e6cc859a6d96d6411e2f6540945c89fd6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf9eaca7b2c7e0c1a287142f3fd574f04aca90819e1ddfdb171172fba994269e864e1d35243c15231e12362c209b880cc0ad59d377295c40ce5d685e62d8beafb2d05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b88d169902011a20c24e302db772704cce373773a92646d8ccb6781f3febb89a2ff3ef4dc5426df40edf7ce083db01ba98eeb1a6dcc15fdd620d315eadc17040586;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9d6beef8c2ee1827b1202b9db787caa13421e75eb42f346d17ff01653e31262a8a89721dcdc2e68dc0d18ac54ad9f087dd39c63fdfba96d66624b5b49a505d14a1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149f32b001fea2481f97449bfee8741f70ae300e23227975ae415e7c462deffda9a2ade3fece28ab78f11ee9479b282adbaca685d551dba3d220e5157694e1627305e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1adbde6e4c1970fc4aeccd5a95793e72b5dd5354ca3286dfc0de088349ec48d746264ab5adb09e2126ddf4bf4eeece20284b4c7a95919f78bf34cc1d2338e8f386f8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hafed347dcecc0290729dc1d40943af5a11e8aaa5ae407ed3e45486c557930668087b12524960854eb64358f0ad8d524373639971e1291a66235612c4ef30718713ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hafdc8ae6bff1520f94f201eda84228470d1b788b35a7b936151ad9c0f1891cbbb392177cc395ec2187cb2fb4e750b219cee5cb50afcc34e3bb597b46b983c701faec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a4053094aa8392093219a53cad34459df08ccacf66cb8217e59ab25dd29b8560c0b235acdb7e4fe56223421e70eb353c6551ecbb809c49938c8dfd5985ee565e8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d9a54c958e922b447ab5706295391ced00274b441438b71bc17ceb57fdc4a03580b01b74121779d2e93b86fd71e054b0bcb66940242d572072b753084604bed9d8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha950801e9d437037619a6c37e6092e7ae2c5315469684d26c830146be0d5ef69a9de6a5a4e9d75cdc8e6fa70073a781d4c9f10d88a0a97d4271c371a7114669c35a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h353cb2c9e4a57367a77578a78249e5d572eb13df6b85d5cd03fadf9c3abd31ed23805f4a6585d209d8bf0711774f87436fa7b0eaa35cf0998228dfc2ef112966583c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ae2d4412fb57863cd658ccda28c82a6233c3e7c62351be63a5f206a72062d080d868dbe9af48d4f5bc6e95db724458d91e6d7774e97043c764d448c90d12ebb3b8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h157a65f6d6b6a0ef5aa525849ad67475e52653698abe6ca2eb95bde0d3802620625c240a69847469c169c65b16aaa7edc876fcd9b4ac4d20da1e13a3b8e0d210e6e3b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7ab0940cc8e40203417987978bd1754c8ba3924c65f6d7c036aee570d2c86c688f270bb10ed001e4a539c9b22bc1d6230e7b3a15c23009d06dac3c07c23b5de3684e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12eedda019bfa136a4c8e50dedfc90fe6d68295bd034ab074366417a259c4acc5395f64a60f73b2fd77c8b92a6865a18b2286fe2865a57c04c2928f445ea2a42a5841;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1897a01e090061df363e53d513c818cf7385c901a24ed9e0f8133846df37e27235750f9cd0e76b97be633ade12c0891f31e45af8f8d638cf2b1649fcd5bcb53f554a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15fa466d92753ba0c12394f8a187af507087555a9202e4376c1956e1ad938928a82962f1a7e16f515001e128ac211e905091ef3734b323cf4928aa2821c7724d7398;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c07416447abfb94587582948b835b49ba129c04bec5b4e7a7b766beb57208c42f852d7bf88c5c9fa0e39e8d2af889ddbfd7188e04d716407636d6f6a5b1ace9cd6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a83eeb7f036a5047d46f5f0432aaf9ae31b749ef77245d0d3649dcb1fb56989e719a664fae3236d0da73414f30d6706dab5fc35afd2ecd2d3b6432847c3fecaf6349;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1830201d6dcdbf98a5c10384076dc17440b64b0b96e32d906cebc7e330517613e168fb374530d5c4fd55296784f9d2ecee932966bd6ba22bcd707712e1ddadc7c470f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17a556276c8136c038a40c04773dca24c3143f461383d38cc71d7e5a2105127ab2f42a29cbf84ba98855cc2d4a694a7ceef81d58ae8275250f2be8e5292737cfc2dbd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea8d8257b2a97afb16d75719027a200eba173264b9a602b0dac9e4c019b58d5b93c16a4c7f68a0c00bf9873ae8bc88f3c7e59d456f4b1d30ae77ce7c8cf38ad26c24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d8e9e27c376d0352f7bd3b28e665c4c455dcffd4a0efa6dfb07af24d277fb4198daca55fcc4f6c62a12ec2c9f0ae6cf33cc5d8eb39b01700f5ecf974c46ec9ba8849;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h77f96af7bd69fa2255989ec08521c8d492b94a8a187ce7f28ae01a874836d18917d3ace63b727887aad45a2c2b4548c1cb6e95e6a0cd1854099d6791ddbb049e3e02;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c8cbf6bcd8bd42b599c64bb7b7352962373134b0d4dcb14e61dc8b9d596d6350365706057ea04894c303dd22d44cb57706cae8628fe9b79a7518bec679de9000a74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h44cec2e10b7d0b23f150b5805b195c142a899ce6394401739371180da71688110e6c7256f6c476e866fc3fab14e207e1cbcd3ce6eaa94722bd1c9d71d096638399b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e78b55fc2bcb642c45546d73d2ca3bde5aaac868e0939352d64c6c100dcb47ca4b5fdf12216c5754ffb66522ed4a015e54dd9a260d75d808669a341f292b80e20f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h128e7225eb8a952897037960b0a920e663f722f7b9bba3a77cf89a1223668eefd8291621a3ca9269c3e80e5d94cb664c23f69d02d1d0bbda74ba5a2f24e0e0ac443ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h404f15d9743b06505eb395d7f548ab0b1972c18216ee9b46c7da7eab6d6b299daf576f4cbc94b9cdf67190e380dbea169ee9c009b0066dac2aeb5acacb445ba188e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e8bce94bc21ca9138307e34e1c9636a34004a6b4d5bd3bfc8dfb663a08a08f24fad41c23d02e57c6b99a1d19d85901be8ad8d4e0be410bc173ce0c49048efe85c050;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dbae87ba11641a392e02ed97d4e1d580d5217d04814aad2951c53d8b704776e9548ed45a3953cb8d30f92365c775f4a1c9dcfed872707e1fdd8fab9310d1769f7ec9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1047e0aba641a6383af72480c7d0a64a584e4a24b9099db0f54d56ed8fed3294feab7110ded4700b535609e2c225299382711bf33f1aa7e9de32fdaab438d6133f3aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17d9aef61252d6c90990638d4d861816bdaf06d0959992aa42fbe3115b95cbf344ef64b22d915a57a34febeb5df0df09101d0eb7fcc31fbd72c642adcccc74d88de47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1362ca8fcc4982d87393ab8eecfa440931f52269902dc7cf7a3e422d537ce295188c2ef46a6d0aecf7fc5d79d3741db911f83581de11ffd97dc9a0e5728dd3e752ec5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h135e97706edafbc1d4b884abf64e426f09e2ac140628808581a7f3f364df07337ec5b692fc370831c3b31fe024913deb84226b73459314e10aec0b5741c3a2bcdcfd0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c83081578a3c827019b8b5d91765e29419823a7faac50aa0f8147ebfa32686ecd95fee995bbe794222eaa8d1d0a7cd1a3b1f9e8847fd8634be33752405bd2c6ef49;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a873c9d248419c35b82a4350bc9e24648c22822ec02580f887ac23dc7e837d854a874fc5b875e7db6ed45bfcdc49c3cc7af4ad9aac5f4e278e54bacc296eb7272786;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67913a516c23664929bc6f629cad508b2406cf492ba52d2438c79f8f14ed84dcb2653fa69320baf45d6c7c8c2bd3925fba504fcd6d48dc319ac090d368238d1df563;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f2e0ca03124e135d82567397bd776435d3917577b309fc9a9357250613fef66e3d927e2dece4e6b669ea8a361cfc4874dbdd315c3373318c86b5d2d2f47187f5a246;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d849648b945b510a071b57561cf2fd139d5c2ebf869602c0509a90db1ae457f20ca199461d6e83632f0ab2e55e2087648fb5e39ff620abd0680353875fd439911a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193c1256f4863bf00e7ac662e1d56fae3f10999832808787bea3483c132d9fe334d39d75f3cd091ba6f8dcf1661c287f295931160066b93f51dba8f93577a4fee6926;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1afcc127ee28ac515c454c272402f82c3ffa21c63aa9c927083c3a6628f98820a4602e5b2d8038ad5dfa55b090c5298c7cf2c52605fd6bba7f355968085aa88b5f915;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1db0e3c859b8aa01c7356bbde68a1b7f753d1dc35d299192b90b5cf05a71fcc2a352c2c0669f42d65e3b16c116da32d33fe16c137857ef9f761a1e6c34799463f77f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6277efcbf4a996eb5f865c4a0e1bb1e179fcb72891ae2de7c6e1084d2b1aee2ea5a25594ba6639e3fa48e4bc0a77c11af9d9c33f6a2a1e202dcfd2b0da27a692c534;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h160a16e8363078177d3be8ebab3f549ef02b52559ffeeefce5b2c8d703151b92c2ed6d46a30f26d81f27d97aedee1b9199db42d16e3a015b874bceccf86ed29e02dec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f56ad94e31ff939132254a2b828f5f4eccf191138e1c1fe469cc13fff61f3d4d4df7ce97213a0509d37f83896dcf3a3f55560a8b2df4f0bc5244f759a8a6093e8790;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c57758471704ff8e11f9a8911347e817b09f0605043bb37681754dbdeecd7e7f466c0eb44973393024357c3cc03bb03aed808f1e43e4f02e92fa12776f46f58d9a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1decfd7a13cfbeb212556a29984a186104e1346b970db5d29acf69d9e63048c935eef1b6397b8a839d487d90d8e4950a579981ea3976aa2a23f644f34b43dc5df9e75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0e83558e62da0eb7f3352a72c8f16fdc154b1ec982fa9e546051a6fa61955e801d64aa84fe21e888687b1f0cf1249ad18ea25556c2427627c10c37a060dfc9b10c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e9214a0c4333d6f66a42f1e4688b49b124983ef4410ada30ad7e0d1009d4a47eede891d5f9cebb7a6b55618807d7bf869ca0d19e918f8824bd1f02a38ca19252c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h152f1879fa08b7a8979eb855f96174740f319702653f65194e6eef3b1ac3b80c2cbf6ba234a53151e4e4774a79f2ca0d11f60702690807bec64a0afba499ba4efb7ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd1dea478b0b5fa5f27e7cdeca75685048ad294f8151e4260b54844c22251280eb4a4bbf2e77b812f0d76716c41f859ce929ddbf9c48f0434d9c373284085c0a1393d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7268e8f1899d0be282c3c23410fe3b57c876f22c0a7cde93fecb3699b98eb53b4f2b486e0c89b60059e0119d6291ca26b2b3e7d4b0c137f33ec0d2bf8b1959acf13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b185fa34fc118b5fadd8b4467a08ff1e48b6498914c8419b1984df638bd0aff98a1a2075f91c65bead6eb686b6cded1fb98163afd9f8b9c7bce41cd6076fd85f776;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13329ec387f59f4c72e99fa5f90d1987849ca634d4b71017c3c1304dc99a623828aab7f12a13f5c41da157ec7a779a6bbe42e0b322239d8de42f920c0289b713ed4e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h778681ae0d9fc4852dd14c7d9d79878ca50fc3719ce3052d21a5449fc5c73ccdb79d6293ebbf757103908df116855786e794b0b1566965117f54c24f7eb87d31dcc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h462451676f19a2a1af9a72540af90d8c5b4a21f52ac2453e14e3372afed13d59cf383d0638baab8d2101f441742d6f73cdbd207662c96b367fed2b591d3bc63ac087;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc3dc8982926ac393048094690e0459aa41920806ccde44f076e9107075d629620c0d93fc73372ede325600360c9b66b2ca6a472664827ea6d34a4902d1864b370df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14e15452efc891296099fe1f9561ff01e47b824dbb687b1a1061d1fa284f9367891f3bf3418533cc4bc1f864ce2231d3ab8537eedb12fd962144f2e1962161a1db975;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1299015ce73988df6fbc97417a007d007b32c5c389935745831e185b70c2c8185538c4227d588f75e46b0f41bff4df20c08261d51c6230a715ed1ffc21f0ec629b94b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1acc9cc32e16db27516a82f15e8a1110987b4d357fc5fc0f388dfeb7bab592687bfd6fbf058d8fafb9f0b723af8b15e05fcb92e7fd20602a279f28f0058430073fbe1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c1eda3f6c9612a8bb0960a8487bc63b4289c01eaf55a3e76720822593eccba2123ebc73394e22f33dbed22e34153dad2ddf4b5fcff5c8bf757eb920e34d793443ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd3e544748278ca9805406cd39efeef9724141c2f671e11b16c160e424a74a0f3c22ea0bccbf62a542a958e352da925ff827c946d9d765f5039263df2887d56ba911;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14daab0880cd6414d01fc6dedb1998e821b5bbd70b843eb2e1ae86a78975f49ea2f5c4a35f55376dbc253ea095f82843f8cf0a3e1856c948839dd1a3a729ddad20d36;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e55e692f88200e89f82ea765c7d097827f05193891a513719e8a3179de40ab892b86d60e0f4c3555bf30b29ad1c4f5612b80ca8f027dee8d76cb9c7ad8b80e35163e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h221af74263732c6073dcb3683382c867f1146ccf599497ef7f323ac0c0fed69e63c8dc27f73d32130a916c42b80c03aa7477d129b76950d72efda3abb847b20307dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6e22d5888b348d91b8bb2f87c26a52e24fbc6a3f69b1cea803fc8abbe97f4dd1de57c2a66028300b4debdc9b9c4e2330ebcf0cefdc3726ead2ed349f7bc0cc9a5a75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1789e47495538dd94388b6562406d5f3e7dfbea2d44afe1ef03caaadccd7f3dc2f7da7e26c09b5b8862dcc0f444375ab174131fedf276f531e544de8ff1acb1c6ceb6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c950dce33b72a272bbb0166d1f581bc922205991ae119461b6304f09924b3b00995a747abc64816348c6cd8baa86129b689fd56b57913c75e7caebb26a63a21cad6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13edc3699cef369543dd8a87d9f6b6cdb6d1235c3ecb5c399896e3f1a672b696d8148b5ec005bcbe1d2e2bb2c85068ec6f97df73b1fc0fcf1fc3eb9158bf302c6a8f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97c62006ca741c4bea17d4bd58c00343f65f2ffe3a9b29e9789c22207ab89126280bea475408dd4c1f75a593f154ef80efac573a7bc867484017ab92f120c3aee7a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97a9ce46c5a7e432c152c7648be09304e4c32d468f9b50ce1c8fd0300e6cd63e83e29f3ee9624793dcc21330e7c3f87ae4a94bae276e4e4d6a241aaf1e698993300a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2083d4ff337612d87596a27832d80576067a7df7d3f16813f0ea2a88985003569a66b4aaa0648de6174bd81636cb3a42af593bc54b01dbe2e5766a004501278685f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h81e328250e1d0704ef52fc42f9561beb73c157fa79619df4db665e91232ec600522917a07c8d65b7b66b0ff24419c8883a33850b586e8539ab2fe8de2fbfdbd0026a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8fd33f9016e65c130de67c7f3c7817dbbcc7b1bf1fedb6f2248ba6f2fc50734f8404caa84811b0a746af4506d406869dae44c878d88740b7c9ecde335545d2d8c35b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbea40e342d75b3c837efd0bc67ccf802a7a732955ef948f2527be19ff3acfe7adece561e183efa3d3da268decaed931c7a84e278bc8b4ec8c15b0dbe58faa31609fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149fcb4612291a9a7100d8eeb639496abed9a3733d73582d4f0eae10df86ca311251d534b80638fc86e7d18ce0cfa2bbebe8d0b5af1d559a5866f74f9cea40d65ad9a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27ec408fa21ee6f0cd6c5ae6ec42f2c2620cff0872a7d35e81fbd7e943c44baca4876dc15cb1bd17e6d21a09d32853894aae77c0152fb8f4363bca74599971da5de2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b9f22f643d7a4c353079a230f975fcc82a4ab835ac3f5006f8a8962ba33fdf346e2da550d360fa86443e0cb71b1b40870ad9053b6a79b9572073705cf24706510dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb1e0d0c3d139a1677df27d42b5161a1ce89dd2ddae99b34afbd10984872dc4285d4404b84256a1e8cb214c80b2c3628e863edc6691c80ca9760928254acad800164;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcb2bedd0b0d994de0de548c614dd005475da1be1024738739736d1fa08f924ee08842c33353779f566030a247dd11b6db9ee6fb464fa81a1a4178e32089fce20158f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1335d5c4afbd055019f2e7a0d4d06ce8fba316b4605cee9fe2599f2e95f6f8c3638944efcb857b79bd70167803fc610883427c422ddc0693573c9ba1305bd00991761;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9af82a1fc72188d2679ed8fa26d64c14b6ca006d377a8a6cb000ee45441ed1a7939b6c3ab9260b42aa8379d6ab66e529e921852bf8e99a6cd81780e7a9d39aecb70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hddfb725d8d4f89b508f50a1da6b83e4c680500510aa2d9686326bc8ebe118e050c39cebc547f1be59eaf03e87d8d5fcd7ac13452f88f97863c5b6a35803d2f4221c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a4f5abe379059413f0dfd33e489ec7aa90a2f5b0f64aa775887c667bdcdc400bc12f2619bcebe297d3422ebf1b9b40aa082b2f50aedc8c0d46fadcccb9af322a4d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd78874e055f4bb45701709ed49a784038307736cf1365424d889d9b08288378e0f3a9c61ad93140cd023de577c76657a41f0ad3e57d224b354ac61fc173cf6b00af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1015b60c3b71c3921edd859680632495fb407f753af9a67f0a2ba4f0a56ab0c61498d3061c39970ecb54bfb716625ae4011d893a7dbc28b62969aa2d9c52fef737314;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2845cff977a1330e17b6515fabda7be4778629e8abbac30f6d49f84fb54c936c918905ef51d84db536c93ff2d907d7b5fc598680417e8a959ffcc002a104634a0f69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c1ad16cc5f2967351a695e5b3b24e4037270ee8ee7a6c3afd9687635d70cc9f68169b87862fcbad37302482476d04345d24d78120a217415f36ce54d2c516e3e35d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1721c9ba9311be0be2eac0207ec9a33747c0873bfe2402725681f1ec2a6f4e3a1b126893e6593e6db113c64bbf1cc5a02e6d508bb28bde80cbfa76ee967576fc43651;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193d2dc71b3339964ad138c1c2f9d5495a08a1f7c572fcef802f4e5e298223f8b4f7da1836f63531b5a83fa7d79e8cbe66cb0b693ca6b4ce157c200a62c31325144a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1983cb43c2e01e55834fb6b99084e3fb012f3377947e52a1a803aa64a2342a4f097741841b37a5ecee74b11623c1170af7ca0f23788823a4ce12786e6fb5226bd2ff8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d8e94e38aa2e832b10855c5c318ab1e40b70fbf3b6b3a5184ffca951cc65cd984779ce8dfc12323e310a081e35b67cd0014a3bc6d7249c0b707975e57f722047136;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb690ed8bafdc766dcf834704e51fd342acb706fd8bd8a06ae440849dd8b17d6617f1cfec4a8cab8e58c9b8f2ae519c8ab55f6716479a45035ad66500962798f13a08;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cfcfe3dc22a664de93ca2482c00bcaffa3d1a78d7c166688d193de579f6fb5216792993c5031731d6d72a9baedafe0d21a5e7bbca318e99a9dc66323358fc410bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce6c26e4b4ac41011b3d79cefd0bdf9aa77445166912d412f3604c45cf661191c76a3f50a6b900fa1ed539899067c2939d3d39d8c9cb125ef34a1fe0543e20a6da94;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h259f27021ac44bf942b11bb606560788b7958a6cf2ce91e2b4d7ce26357e75ca45001e1b35dc53d9d6773d05f59d9d7f00f96ce5be52e828c5a83d0e60f63cd8e110;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1058d6611aef15649dd559527cfb3e26be3c9286fc69b4a9fa9c0a2c4aad81822866b27a7827f27e4658954057b735ce79022444e033de594b39b2777a71f8cdcc8b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2541be51f7ea7cdea8e31af06a91da5cd0dd08e161535662b261eb77d68f40d4e54862936edb67da1aa2fb333e18978cab749126dbacda2ae368132b4ce3210ec15d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0df39ca21ae230eed6f64b56daee1f388d06a5649fc8b447c56a066e5ee1b7f44b7793779a8cb688ea7e58826cef47031bc1be4bc1e5cef5d97d3e5a63469361333;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h822c7ced1f4bd97a4251e9c2be25d9a371c8e40dae83af6b0b9789493583470d3c28f38704da6d877e60a918d1f292aca1acfae0ee4fcb77bd9ed98318962190c020;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha33c6c34eadadf8ad52e3e6fbbdbb0828afbe07b00dfbd39262c05bd732572a172fbe438dfd74f62cae5fbe59af24de045e26d4712f9085c6f416889af8c7159cd49;
        #1
        $finish();
    end
endmodule
