module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70,
        output wire [0:0] dst71);
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    reg [255:0] src16;
    reg [255:0] src17;
    reg [255:0] src18;
    reg [255:0] src19;
    reg [255:0] src20;
    reg [255:0] src21;
    reg [255:0] src22;
    reg [255:0] src23;
    reg [255:0] src24;
    reg [255:0] src25;
    reg [255:0] src26;
    reg [255:0] src27;
    reg [255:0] src28;
    reg [255:0] src29;
    reg [255:0] src30;
    reg [255:0] src31;
    reg [255:0] src32;
    reg [255:0] src33;
    reg [255:0] src34;
    reg [255:0] src35;
    reg [255:0] src36;
    reg [255:0] src37;
    reg [255:0] src38;
    reg [255:0] src39;
    reg [255:0] src40;
    reg [255:0] src41;
    reg [255:0] src42;
    reg [255:0] src43;
    reg [255:0] src44;
    reg [255:0] src45;
    reg [255:0] src46;
    reg [255:0] src47;
    reg [255:0] src48;
    reg [255:0] src49;
    reg [255:0] src50;
    reg [255:0] src51;
    reg [255:0] src52;
    reg [255:0] src53;
    reg [255:0] src54;
    reg [255:0] src55;
    reg [255:0] src56;
    reg [255:0] src57;
    reg [255:0] src58;
    reg [255:0] src59;
    reg [255:0] src60;
    reg [255:0] src61;
    reg [255:0] src62;
    reg [255:0] src63;
    compressor_CLA256_64 compressor_CLA256_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70),
            .dst71(dst71));
    initial begin
        src0 <= 256'h0;
        src1 <= 256'h0;
        src2 <= 256'h0;
        src3 <= 256'h0;
        src4 <= 256'h0;
        src5 <= 256'h0;
        src6 <= 256'h0;
        src7 <= 256'h0;
        src8 <= 256'h0;
        src9 <= 256'h0;
        src10 <= 256'h0;
        src11 <= 256'h0;
        src12 <= 256'h0;
        src13 <= 256'h0;
        src14 <= 256'h0;
        src15 <= 256'h0;
        src16 <= 256'h0;
        src17 <= 256'h0;
        src18 <= 256'h0;
        src19 <= 256'h0;
        src20 <= 256'h0;
        src21 <= 256'h0;
        src22 <= 256'h0;
        src23 <= 256'h0;
        src24 <= 256'h0;
        src25 <= 256'h0;
        src26 <= 256'h0;
        src27 <= 256'h0;
        src28 <= 256'h0;
        src29 <= 256'h0;
        src30 <= 256'h0;
        src31 <= 256'h0;
        src32 <= 256'h0;
        src33 <= 256'h0;
        src34 <= 256'h0;
        src35 <= 256'h0;
        src36 <= 256'h0;
        src37 <= 256'h0;
        src38 <= 256'h0;
        src39 <= 256'h0;
        src40 <= 256'h0;
        src41 <= 256'h0;
        src42 <= 256'h0;
        src43 <= 256'h0;
        src44 <= 256'h0;
        src45 <= 256'h0;
        src46 <= 256'h0;
        src47 <= 256'h0;
        src48 <= 256'h0;
        src49 <= 256'h0;
        src50 <= 256'h0;
        src51 <= 256'h0;
        src52 <= 256'h0;
        src53 <= 256'h0;
        src54 <= 256'h0;
        src55 <= 256'h0;
        src56 <= 256'h0;
        src57 <= 256'h0;
        src58 <= 256'h0;
        src59 <= 256'h0;
        src60 <= 256'h0;
        src61 <= 256'h0;
        src62 <= 256'h0;
        src63 <= 256'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA256_64(
    input [255:0]src0,
    input [255:0]src1,
    input [255:0]src2,
    input [255:0]src3,
    input [255:0]src4,
    input [255:0]src5,
    input [255:0]src6,
    input [255:0]src7,
    input [255:0]src8,
    input [255:0]src9,
    input [255:0]src10,
    input [255:0]src11,
    input [255:0]src12,
    input [255:0]src13,
    input [255:0]src14,
    input [255:0]src15,
    input [255:0]src16,
    input [255:0]src17,
    input [255:0]src18,
    input [255:0]src19,
    input [255:0]src20,
    input [255:0]src21,
    input [255:0]src22,
    input [255:0]src23,
    input [255:0]src24,
    input [255:0]src25,
    input [255:0]src26,
    input [255:0]src27,
    input [255:0]src28,
    input [255:0]src29,
    input [255:0]src30,
    input [255:0]src31,
    input [255:0]src32,
    input [255:0]src33,
    input [255:0]src34,
    input [255:0]src35,
    input [255:0]src36,
    input [255:0]src37,
    input [255:0]src38,
    input [255:0]src39,
    input [255:0]src40,
    input [255:0]src41,
    input [255:0]src42,
    input [255:0]src43,
    input [255:0]src44,
    input [255:0]src45,
    input [255:0]src46,
    input [255:0]src47,
    input [255:0]src48,
    input [255:0]src49,
    input [255:0]src50,
    input [255:0]src51,
    input [255:0]src52,
    input [255:0]src53,
    input [255:0]src54,
    input [255:0]src55,
    input [255:0]src56,
    input [255:0]src57,
    input [255:0]src58,
    input [255:0]src59,
    input [255:0]src60,
    input [255:0]src61,
    input [255:0]src62,
    input [255:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70,
    output dst71);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [0:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [0:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [0:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [0:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [1:0] comp_out69;
    wire [1:0] comp_out70;
    wire [0:0] comp_out71;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70),
        .dst71(comp_out71)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out71[0], comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out70[1], comp_out69[1], comp_out68[1], comp_out67[1], comp_out66[1], 1'h0, comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], 1'h0, comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], 1'h0, comp_out33[1], comp_out32[1], 1'h0, comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], 1'h0}),
        .dst({dst71, dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [255:0] src0,
      input wire [255:0] src1,
      input wire [255:0] src2,
      input wire [255:0] src3,
      input wire [255:0] src4,
      input wire [255:0] src5,
      input wire [255:0] src6,
      input wire [255:0] src7,
      input wire [255:0] src8,
      input wire [255:0] src9,
      input wire [255:0] src10,
      input wire [255:0] src11,
      input wire [255:0] src12,
      input wire [255:0] src13,
      input wire [255:0] src14,
      input wire [255:0] src15,
      input wire [255:0] src16,
      input wire [255:0] src17,
      input wire [255:0] src18,
      input wire [255:0] src19,
      input wire [255:0] src20,
      input wire [255:0] src21,
      input wire [255:0] src22,
      input wire [255:0] src23,
      input wire [255:0] src24,
      input wire [255:0] src25,
      input wire [255:0] src26,
      input wire [255:0] src27,
      input wire [255:0] src28,
      input wire [255:0] src29,
      input wire [255:0] src30,
      input wire [255:0] src31,
      input wire [255:0] src32,
      input wire [255:0] src33,
      input wire [255:0] src34,
      input wire [255:0] src35,
      input wire [255:0] src36,
      input wire [255:0] src37,
      input wire [255:0] src38,
      input wire [255:0] src39,
      input wire [255:0] src40,
      input wire [255:0] src41,
      input wire [255:0] src42,
      input wire [255:0] src43,
      input wire [255:0] src44,
      input wire [255:0] src45,
      input wire [255:0] src46,
      input wire [255:0] src47,
      input wire [255:0] src48,
      input wire [255:0] src49,
      input wire [255:0] src50,
      input wire [255:0] src51,
      input wire [255:0] src52,
      input wire [255:0] src53,
      input wire [255:0] src54,
      input wire [255:0] src55,
      input wire [255:0] src56,
      input wire [255:0] src57,
      input wire [255:0] src58,
      input wire [255:0] src59,
      input wire [255:0] src60,
      input wire [255:0] src61,
      input wire [255:0] src62,
      input wire [255:0] src63,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [0:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [0:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [0:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [0:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [1:0] dst69,
      output wire [1:0] dst70,
      output wire [0:0] dst71);

   wire [255:0] stage0_0;
   wire [255:0] stage0_1;
   wire [255:0] stage0_2;
   wire [255:0] stage0_3;
   wire [255:0] stage0_4;
   wire [255:0] stage0_5;
   wire [255:0] stage0_6;
   wire [255:0] stage0_7;
   wire [255:0] stage0_8;
   wire [255:0] stage0_9;
   wire [255:0] stage0_10;
   wire [255:0] stage0_11;
   wire [255:0] stage0_12;
   wire [255:0] stage0_13;
   wire [255:0] stage0_14;
   wire [255:0] stage0_15;
   wire [255:0] stage0_16;
   wire [255:0] stage0_17;
   wire [255:0] stage0_18;
   wire [255:0] stage0_19;
   wire [255:0] stage0_20;
   wire [255:0] stage0_21;
   wire [255:0] stage0_22;
   wire [255:0] stage0_23;
   wire [255:0] stage0_24;
   wire [255:0] stage0_25;
   wire [255:0] stage0_26;
   wire [255:0] stage0_27;
   wire [255:0] stage0_28;
   wire [255:0] stage0_29;
   wire [255:0] stage0_30;
   wire [255:0] stage0_31;
   wire [255:0] stage0_32;
   wire [255:0] stage0_33;
   wire [255:0] stage0_34;
   wire [255:0] stage0_35;
   wire [255:0] stage0_36;
   wire [255:0] stage0_37;
   wire [255:0] stage0_38;
   wire [255:0] stage0_39;
   wire [255:0] stage0_40;
   wire [255:0] stage0_41;
   wire [255:0] stage0_42;
   wire [255:0] stage0_43;
   wire [255:0] stage0_44;
   wire [255:0] stage0_45;
   wire [255:0] stage0_46;
   wire [255:0] stage0_47;
   wire [255:0] stage0_48;
   wire [255:0] stage0_49;
   wire [255:0] stage0_50;
   wire [255:0] stage0_51;
   wire [255:0] stage0_52;
   wire [255:0] stage0_53;
   wire [255:0] stage0_54;
   wire [255:0] stage0_55;
   wire [255:0] stage0_56;
   wire [255:0] stage0_57;
   wire [255:0] stage0_58;
   wire [255:0] stage0_59;
   wire [255:0] stage0_60;
   wire [255:0] stage0_61;
   wire [255:0] stage0_62;
   wire [255:0] stage0_63;
   wire [90:0] stage1_0;
   wire [82:0] stage1_1;
   wire [130:0] stage1_2;
   wire [106:0] stage1_3;
   wire [121:0] stage1_4;
   wire [95:0] stage1_5;
   wire [115:0] stage1_6;
   wire [109:0] stage1_7;
   wire [131:0] stage1_8;
   wire [119:0] stage1_9;
   wire [155:0] stage1_10;
   wire [153:0] stage1_11;
   wire [132:0] stage1_12;
   wire [96:0] stage1_13;
   wire [84:0] stage1_14;
   wire [131:0] stage1_15;
   wire [119:0] stage1_16;
   wire [110:0] stage1_17;
   wire [99:0] stage1_18;
   wire [125:0] stage1_19;
   wire [129:0] stage1_20;
   wire [107:0] stage1_21;
   wire [91:0] stage1_22;
   wire [128:0] stage1_23;
   wire [139:0] stage1_24;
   wire [109:0] stage1_25;
   wire [140:0] stage1_26;
   wire [118:0] stage1_27;
   wire [126:0] stage1_28;
   wire [109:0] stage1_29;
   wire [90:0] stage1_30;
   wire [114:0] stage1_31;
   wire [114:0] stage1_32;
   wire [110:0] stage1_33;
   wire [103:0] stage1_34;
   wire [118:0] stage1_35;
   wire [144:0] stage1_36;
   wire [104:0] stage1_37;
   wire [136:0] stage1_38;
   wire [124:0] stage1_39;
   wire [91:0] stage1_40;
   wire [142:0] stage1_41;
   wire [171:0] stage1_42;
   wire [78:0] stage1_43;
   wire [145:0] stage1_44;
   wire [158:0] stage1_45;
   wire [100:0] stage1_46;
   wire [129:0] stage1_47;
   wire [107:0] stage1_48;
   wire [151:0] stage1_49;
   wire [98:0] stage1_50;
   wire [105:0] stage1_51;
   wire [139:0] stage1_52;
   wire [107:0] stage1_53;
   wire [159:0] stage1_54;
   wire [89:0] stage1_55;
   wire [177:0] stage1_56;
   wire [104:0] stage1_57;
   wire [85:0] stage1_58;
   wire [147:0] stage1_59;
   wire [141:0] stage1_60;
   wire [108:0] stage1_61;
   wire [200:0] stage1_62;
   wire [68:0] stage1_63;
   wire [63:0] stage1_64;
   wire [41:0] stage1_65;
   wire [29:0] stage2_0;
   wire [36:0] stage2_1;
   wire [36:0] stage2_2;
   wire [53:0] stage2_3;
   wire [44:0] stage2_4;
   wire [45:0] stage2_5;
   wire [51:0] stage2_6;
   wire [42:0] stage2_7;
   wire [42:0] stage2_8;
   wire [59:0] stage2_9;
   wire [69:0] stage2_10;
   wire [48:0] stage2_11;
   wire [53:0] stage2_12;
   wire [63:0] stage2_13;
   wire [44:0] stage2_14;
   wire [73:0] stage2_15;
   wire [54:0] stage2_16;
   wire [56:0] stage2_17;
   wire [65:0] stage2_18;
   wire [36:0] stage2_19;
   wire [79:0] stage2_20;
   wire [48:0] stage2_21;
   wire [40:0] stage2_22;
   wire [60:0] stage2_23;
   wire [81:0] stage2_24;
   wire [50:0] stage2_25;
   wire [51:0] stage2_26;
   wire [71:0] stage2_27;
   wire [72:0] stage2_28;
   wire [45:0] stage2_29;
   wire [58:0] stage2_30;
   wire [53:0] stage2_31;
   wire [46:0] stage2_32;
   wire [51:0] stage2_33;
   wire [36:0] stage2_34;
   wire [58:0] stage2_35;
   wire [62:0] stage2_36;
   wire [54:0] stage2_37;
   wire [46:0] stage2_38;
   wire [80:0] stage2_39;
   wire [44:0] stage2_40;
   wire [74:0] stage2_41;
   wire [62:0] stage2_42;
   wire [61:0] stage2_43;
   wire [51:0] stage2_44;
   wire [78:0] stage2_45;
   wire [62:0] stage2_46;
   wire [70:0] stage2_47;
   wire [41:0] stage2_48;
   wire [114:0] stage2_49;
   wire [67:0] stage2_50;
   wire [78:0] stage2_51;
   wire [50:0] stage2_52;
   wire [77:0] stage2_53;
   wire [74:0] stage2_54;
   wire [34:0] stage2_55;
   wire [72:0] stage2_56;
   wire [82:0] stage2_57;
   wire [47:0] stage2_58;
   wire [47:0] stage2_59;
   wire [62:0] stage2_60;
   wire [56:0] stage2_61;
   wire [52:0] stage2_62;
   wire [74:0] stage2_63;
   wire [44:0] stage2_64;
   wire [17:0] stage2_65;
   wire [16:0] stage2_66;
   wire [6:0] stage2_67;
   wire [13:0] stage3_0;
   wire [10:0] stage3_1;
   wire [17:0] stage3_2;
   wire [18:0] stage3_3;
   wire [20:0] stage3_4;
   wire [34:0] stage3_5;
   wire [16:0] stage3_6;
   wire [27:0] stage3_7;
   wire [17:0] stage3_8;
   wire [15:0] stage3_9;
   wire [32:0] stage3_10;
   wire [30:0] stage3_11;
   wire [24:0] stage3_12;
   wire [23:0] stage3_13;
   wire [26:0] stage3_14;
   wire [40:0] stage3_15;
   wire [19:0] stage3_16;
   wire [29:0] stage3_17;
   wire [27:0] stage3_18;
   wire [27:0] stage3_19;
   wire [23:0] stage3_20;
   wire [23:0] stage3_21;
   wire [28:0] stage3_22;
   wire [15:0] stage3_23;
   wire [30:0] stage3_24;
   wire [33:0] stage3_25;
   wire [23:0] stage3_26;
   wire [21:0] stage3_27;
   wire [28:0] stage3_28;
   wire [34:0] stage3_29;
   wire [25:0] stage3_30;
   wire [31:0] stage3_31;
   wire [27:0] stage3_32;
   wire [26:0] stage3_33;
   wire [26:0] stage3_34;
   wire [32:0] stage3_35;
   wire [19:0] stage3_36;
   wire [18:0] stage3_37;
   wire [22:0] stage3_38;
   wire [30:0] stage3_39;
   wire [29:0] stage3_40;
   wire [23:0] stage3_41;
   wire [29:0] stage3_42;
   wire [38:0] stage3_43;
   wire [21:0] stage3_44;
   wire [38:0] stage3_45;
   wire [39:0] stage3_46;
   wire [32:0] stage3_47;
   wire [23:0] stage3_48;
   wire [67:0] stage3_49;
   wire [29:0] stage3_50;
   wire [47:0] stage3_51;
   wire [39:0] stage3_52;
   wire [27:0] stage3_53;
   wire [27:0] stage3_54;
   wire [29:0] stage3_55;
   wire [25:0] stage3_56;
   wire [32:0] stage3_57;
   wire [28:0] stage3_58;
   wire [32:0] stage3_59;
   wire [34:0] stage3_60;
   wire [23:0] stage3_61;
   wire [27:0] stage3_62;
   wire [27:0] stage3_63;
   wire [17:0] stage3_64;
   wire [27:0] stage3_65;
   wire [27:0] stage3_66;
   wire [1:0] stage3_67;
   wire [0:0] stage3_68;
   wire [0:0] stage3_69;
   wire [13:0] stage4_0;
   wire [4:0] stage4_1;
   wire [6:0] stage4_2;
   wire [18:0] stage4_3;
   wire [9:0] stage4_4;
   wire [19:0] stage4_5;
   wire [9:0] stage4_6;
   wire [9:0] stage4_7;
   wire [21:0] stage4_8;
   wire [7:0] stage4_9;
   wire [13:0] stage4_10;
   wire [11:0] stage4_11;
   wire [17:0] stage4_12;
   wire [13:0] stage4_13;
   wire [11:0] stage4_14;
   wire [11:0] stage4_15;
   wire [12:0] stage4_16;
   wire [14:0] stage4_17;
   wire [10:0] stage4_18;
   wire [13:0] stage4_19;
   wire [10:0] stage4_20;
   wire [8:0] stage4_21;
   wire [14:0] stage4_22;
   wire [8:0] stage4_23;
   wire [11:0] stage4_24;
   wire [13:0] stage4_25;
   wire [12:0] stage4_26;
   wire [6:0] stage4_27;
   wire [11:0] stage4_28;
   wire [16:0] stage4_29;
   wire [11:0] stage4_30;
   wire [9:0] stage4_31;
   wire [17:0] stage4_32;
   wire [16:0] stage4_33;
   wire [10:0] stage4_34;
   wire [16:0] stage4_35;
   wire [12:0] stage4_36;
   wire [11:0] stage4_37;
   wire [6:0] stage4_38;
   wire [8:0] stage4_39;
   wire [12:0] stage4_40;
   wire [11:0] stage4_41;
   wire [14:0] stage4_42;
   wire [19:0] stage4_43;
   wire [13:0] stage4_44;
   wire [11:0] stage4_45;
   wire [14:0] stage4_46;
   wire [14:0] stage4_47;
   wire [14:0] stage4_48;
   wire [35:0] stage4_49;
   wire [16:0] stage4_50;
   wire [19:0] stage4_51;
   wire [13:0] stage4_52;
   wire [14:0] stage4_53;
   wire [17:0] stage4_54;
   wire [12:0] stage4_55;
   wire [11:0] stage4_56;
   wire [11:0] stage4_57;
   wire [19:0] stage4_58;
   wire [11:0] stage4_59;
   wire [13:0] stage4_60;
   wire [11:0] stage4_61;
   wire [11:0] stage4_62;
   wire [12:0] stage4_63;
   wire [11:0] stage4_64;
   wire [7:0] stage4_65;
   wire [23:0] stage4_66;
   wire [8:0] stage4_67;
   wire [2:0] stage4_68;
   wire [0:0] stage4_69;
   wire [4:0] stage5_0;
   wire [3:0] stage5_1;
   wire [1:0] stage5_2;
   wire [6:0] stage5_3;
   wire [9:0] stage5_4;
   wire [7:0] stage5_5;
   wire [5:0] stage5_6;
   wire [6:0] stage5_7;
   wire [4:0] stage5_8;
   wire [9:0] stage5_9;
   wire [5:0] stage5_10;
   wire [9:0] stage5_11;
   wire [5:0] stage5_12;
   wire [5:0] stage5_13;
   wire [4:0] stage5_14;
   wire [5:0] stage5_15;
   wire [5:0] stage5_16;
   wire [7:0] stage5_17;
   wire [5:0] stage5_18;
   wire [10:0] stage5_19;
   wire [2:0] stage5_20;
   wire [11:0] stage5_21;
   wire [4:0] stage5_22;
   wire [2:0] stage5_23;
   wire [6:0] stage5_24;
   wire [5:0] stage5_25;
   wire [5:0] stage5_26;
   wire [5:0] stage5_27;
   wire [3:0] stage5_28;
   wire [7:0] stage5_29;
   wire [5:0] stage5_30;
   wire [6:0] stage5_31;
   wire [3:0] stage5_32;
   wire [6:0] stage5_33;
   wire [6:0] stage5_34;
   wire [4:0] stage5_35;
   wire [6:0] stage5_36;
   wire [11:0] stage5_37;
   wire [3:0] stage5_38;
   wire [2:0] stage5_39;
   wire [5:0] stage5_40;
   wire [4:0] stage5_41;
   wire [6:0] stage5_42;
   wire [9:0] stage5_43;
   wire [6:0] stage5_44;
   wire [4:0] stage5_45;
   wire [6:0] stage5_46;
   wire [6:0] stage5_47;
   wire [6:0] stage5_48;
   wire [7:0] stage5_49;
   wire [8:0] stage5_50;
   wire [9:0] stage5_51;
   wire [7:0] stage5_52;
   wire [14:0] stage5_53;
   wire [5:0] stage5_54;
   wire [5:0] stage5_55;
   wire [5:0] stage5_56;
   wire [6:0] stage5_57;
   wire [4:0] stage5_58;
   wire [6:0] stage5_59;
   wire [8:0] stage5_60;
   wire [3:0] stage5_61;
   wire [3:0] stage5_62;
   wire [5:0] stage5_63;
   wire [5:0] stage5_64;
   wire [4:0] stage5_65;
   wire [10:0] stage5_66;
   wire [6:0] stage5_67;
   wire [4:0] stage5_68;
   wire [2:0] stage5_69;
   wire [4:0] stage6_0;
   wire [3:0] stage6_1;
   wire [0:0] stage6_2;
   wire [1:0] stage6_3;
   wire [4:0] stage6_4;
   wire [3:0] stage6_5;
   wire [1:0] stage6_6;
   wire [2:0] stage6_7;
   wire [2:0] stage6_8;
   wire [8:0] stage6_9;
   wire [1:0] stage6_10;
   wire [5:0] stage6_11;
   wire [2:0] stage6_12;
   wire [1:0] stage6_13;
   wire [6:0] stage6_14;
   wire [2:0] stage6_15;
   wire [1:0] stage6_16;
   wire [2:0] stage6_17;
   wire [3:0] stage6_18;
   wire [3:0] stage6_19;
   wire [3:0] stage6_20;
   wire [1:0] stage6_21;
   wire [2:0] stage6_22;
   wire [4:0] stage6_23;
   wire [1:0] stage6_24;
   wire [6:0] stage6_25;
   wire [1:0] stage6_26;
   wire [2:0] stage6_27;
   wire [1:0] stage6_28;
   wire [2:0] stage6_29;
   wire [2:0] stage6_30;
   wire [2:0] stage6_31;
   wire [2:0] stage6_32;
   wire [3:0] stage6_33;
   wire [2:0] stage6_34;
   wire [3:0] stage6_35;
   wire [3:0] stage6_36;
   wire [7:0] stage6_37;
   wire [1:0] stage6_38;
   wire [2:0] stage6_39;
   wire [1:0] stage6_40;
   wire [1:0] stage6_41;
   wire [2:0] stage6_42;
   wire [5:0] stage6_43;
   wire [2:0] stage6_44;
   wire [3:0] stage6_45;
   wire [1:0] stage6_46;
   wire [5:0] stage6_47;
   wire [3:0] stage6_48;
   wire [2:0] stage6_49;
   wire [3:0] stage6_50;
   wire [4:0] stage6_51;
   wire [2:0] stage6_52;
   wire [3:0] stage6_53;
   wire [3:0] stage6_54;
   wire [3:0] stage6_55;
   wire [5:0] stage6_56;
   wire [2:0] stage6_57;
   wire [1:0] stage6_58;
   wire [5:0] stage6_59;
   wire [4:0] stage6_60;
   wire [4:0] stage6_61;
   wire [4:0] stage6_62;
   wire [0:0] stage6_63;
   wire [1:0] stage6_64;
   wire [1:0] stage6_65;
   wire [2:0] stage6_66;
   wire [4:0] stage6_67;
   wire [2:0] stage6_68;
   wire [1:0] stage6_69;
   wire [1:0] stage6_70;
   wire [0:0] stage6_71;
   wire [0:0] stage7_0;
   wire [1:0] stage7_1;
   wire [0:0] stage7_2;
   wire [1:0] stage7_3;
   wire [1:0] stage7_4;
   wire [1:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [1:0] stage7_19;
   wire [1:0] stage7_20;
   wire [1:0] stage7_21;
   wire [1:0] stage7_22;
   wire [1:0] stage7_23;
   wire [1:0] stage7_24;
   wire [1:0] stage7_25;
   wire [1:0] stage7_26;
   wire [1:0] stage7_27;
   wire [1:0] stage7_28;
   wire [1:0] stage7_29;
   wire [1:0] stage7_30;
   wire [0:0] stage7_31;
   wire [1:0] stage7_32;
   wire [1:0] stage7_33;
   wire [0:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [1:0] stage7_37;
   wire [1:0] stage7_38;
   wire [1:0] stage7_39;
   wire [1:0] stage7_40;
   wire [1:0] stage7_41;
   wire [1:0] stage7_42;
   wire [1:0] stage7_43;
   wire [1:0] stage7_44;
   wire [1:0] stage7_45;
   wire [1:0] stage7_46;
   wire [0:0] stage7_47;
   wire [1:0] stage7_48;
   wire [1:0] stage7_49;
   wire [1:0] stage7_50;
   wire [1:0] stage7_51;
   wire [1:0] stage7_52;
   wire [1:0] stage7_53;
   wire [1:0] stage7_54;
   wire [1:0] stage7_55;
   wire [1:0] stage7_56;
   wire [1:0] stage7_57;
   wire [1:0] stage7_58;
   wire [1:0] stage7_59;
   wire [1:0] stage7_60;
   wire [1:0] stage7_61;
   wire [1:0] stage7_62;
   wire [1:0] stage7_63;
   wire [1:0] stage7_64;
   wire [0:0] stage7_65;
   wire [1:0] stage7_66;
   wire [1:0] stage7_67;
   wire [1:0] stage7_68;
   wire [1:0] stage7_69;
   wire [1:0] stage7_70;
   wire [0:0] stage7_71;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;
   assign dst21 = stage7_21;
   assign dst22 = stage7_22;
   assign dst23 = stage7_23;
   assign dst24 = stage7_24;
   assign dst25 = stage7_25;
   assign dst26 = stage7_26;
   assign dst27 = stage7_27;
   assign dst28 = stage7_28;
   assign dst29 = stage7_29;
   assign dst30 = stage7_30;
   assign dst31 = stage7_31;
   assign dst32 = stage7_32;
   assign dst33 = stage7_33;
   assign dst34 = stage7_34;
   assign dst35 = stage7_35;
   assign dst36 = stage7_36;
   assign dst37 = stage7_37;
   assign dst38 = stage7_38;
   assign dst39 = stage7_39;
   assign dst40 = stage7_40;
   assign dst41 = stage7_41;
   assign dst42 = stage7_42;
   assign dst43 = stage7_43;
   assign dst44 = stage7_44;
   assign dst45 = stage7_45;
   assign dst46 = stage7_46;
   assign dst47 = stage7_47;
   assign dst48 = stage7_48;
   assign dst49 = stage7_49;
   assign dst50 = stage7_50;
   assign dst51 = stage7_51;
   assign dst52 = stage7_52;
   assign dst53 = stage7_53;
   assign dst54 = stage7_54;
   assign dst55 = stage7_55;
   assign dst56 = stage7_56;
   assign dst57 = stage7_57;
   assign dst58 = stage7_58;
   assign dst59 = stage7_59;
   assign dst60 = stage7_60;
   assign dst61 = stage7_61;
   assign dst62 = stage7_62;
   assign dst63 = stage7_63;
   assign dst64 = stage7_64;
   assign dst65 = stage7_65;
   assign dst66 = stage7_66;
   assign dst67 = stage7_67;
   assign dst68 = stage7_68;
   assign dst69 = stage7_69;
   assign dst70 = stage7_70;
   assign dst71 = stage7_71;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[10]},
      {stage0_3[20]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[11]},
      {stage0_3[21]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[56], stage0_0[57], stage0_0[58]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[12]},
      {stage0_3[22]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[59], stage0_0[60], stage0_0[61]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[13]},
      {stage0_3[23]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[62], stage0_0[63], stage0_0[64]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[14]},
      {stage0_3[24]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[65], stage0_0[66], stage0_0[67]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[15]},
      {stage0_3[25]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[68], stage0_0[69], stage0_0[70]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[16]},
      {stage0_3[26]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[71], stage0_0[72], stage0_0[73]},
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_2[17]},
      {stage0_3[27]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[74], stage0_0[75], stage0_0[76]},
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_2[18]},
      {stage0_3[28]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[77], stage0_0[78], stage0_0[79]},
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_2[19]},
      {stage0_3[29]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[80], stage0_0[81], stage0_0[82]},
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_2[20]},
      {stage0_3[30]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[83], stage0_0[84], stage0_0[85]},
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_2[21]},
      {stage0_3[31]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[86], stage0_0[87], stage0_0[88]},
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_2[22]},
      {stage0_3[32]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[89], stage0_0[90], stage0_0[91]},
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_2[23]},
      {stage0_3[33]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[92], stage0_0[93], stage0_0[94]},
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_2[24]},
      {stage0_3[34]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[95], stage0_0[96], stage0_0[97]},
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_2[25]},
      {stage0_3[35]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[98], stage0_0[99], stage0_0[100]},
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_2[26]},
      {stage0_3[36]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[101], stage0_0[102], stage0_0[103]},
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_2[27]},
      {stage0_3[37]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[104], stage0_0[105], stage0_0[106]},
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_2[28]},
      {stage0_3[38]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[107], stage0_0[108], stage0_0[109]},
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_2[29]},
      {stage0_3[39]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139]},
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59]},
      {stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145]},
      {stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65]},
      {stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[146], stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151]},
      {stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71]},
      {stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[152], stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157]},
      {stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77]},
      {stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[158], stage0_0[159], stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163]},
      {stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83]},
      {stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[164], stage0_0[165], stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169]},
      {stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89]},
      {stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[170], stage0_0[171], stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175]},
      {stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95]},
      {stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[176], stage0_0[177], stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181]},
      {stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101]},
      {stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[182], stage0_0[183], stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187]},
      {stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107]},
      {stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[188], stage0_0[189], stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193]},
      {stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113]},
      {stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[194], stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199]},
      {stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119]},
      {stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205]},
      {stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211]},
      {stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131]},
      {stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45]},
      {stage1_5[0],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage1_5[1],stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57]},
      {stage1_5[2],stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage1_5[3],stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69]},
      {stage1_5[4],stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc606_5 gpc52 (
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75]},
      {stage1_5[5],stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52]}
   );
   gpc606_5 gpc53 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81]},
      {stage1_5[6],stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53]}
   );
   gpc606_5 gpc54 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87]},
      {stage1_5[7],stage1_4[54],stage1_3[54],stage1_2[54],stage1_1[54]}
   );
   gpc606_5 gpc55 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93]},
      {stage1_5[8],stage1_4[55],stage1_3[55],stage1_2[55],stage1_1[55]}
   );
   gpc606_5 gpc56 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage1_5[9],stage1_4[56],stage1_3[56],stage1_2[56],stage1_1[56]}
   );
   gpc606_5 gpc57 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105]},
      {stage1_5[10],stage1_4[57],stage1_3[57],stage1_2[57],stage1_1[57]}
   );
   gpc606_5 gpc58 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage1_5[11],stage1_4[58],stage1_3[58],stage1_2[58],stage1_1[58]}
   );
   gpc606_5 gpc59 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117]},
      {stage1_5[12],stage1_4[59],stage1_3[59],stage1_2[59],stage1_1[59]}
   );
   gpc606_5 gpc60 (
      {stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233]},
      {stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage1_5[13],stage1_4[60],stage1_3[60],stage1_2[60],stage1_1[60]}
   );
   gpc606_5 gpc61 (
      {stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[14],stage1_4[61],stage1_3[61],stage1_2[61]}
   );
   gpc606_5 gpc62 (
      {stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[15],stage1_4[62],stage1_3[62],stage1_2[62]}
   );
   gpc615_5 gpc63 (
      {stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148]},
      {stage0_3[124]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[16],stage1_4[63],stage1_3[63],stage1_2[63]}
   );
   gpc615_5 gpc64 (
      {stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153]},
      {stage0_3[125]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[17],stage1_4[64],stage1_3[64],stage1_2[64]}
   );
   gpc615_5 gpc65 (
      {stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage0_3[126]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[18],stage1_4[65],stage1_3[65],stage1_2[65]}
   );
   gpc615_5 gpc66 (
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163]},
      {stage0_3[127]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[19],stage1_4[66],stage1_3[66],stage1_2[66]}
   );
   gpc615_5 gpc67 (
      {stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168]},
      {stage0_3[128]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[20],stage1_4[67],stage1_3[67],stage1_2[67]}
   );
   gpc615_5 gpc68 (
      {stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173]},
      {stage0_3[129]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[21],stage1_4[68],stage1_3[68],stage1_2[68]}
   );
   gpc615_5 gpc69 (
      {stage0_2[174], stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178]},
      {stage0_3[130]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[22],stage1_4[69],stage1_3[69],stage1_2[69]}
   );
   gpc615_5 gpc70 (
      {stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182], stage0_2[183]},
      {stage0_3[131]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[23],stage1_4[70],stage1_3[70],stage1_2[70]}
   );
   gpc615_5 gpc71 (
      {stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage0_3[132]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[24],stage1_4[71],stage1_3[71],stage1_2[71]}
   );
   gpc615_5 gpc72 (
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193]},
      {stage0_3[133]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[25],stage1_4[72],stage1_3[72],stage1_2[72]}
   );
   gpc615_5 gpc73 (
      {stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198]},
      {stage0_3[134]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[26],stage1_4[73],stage1_3[73],stage1_2[73]}
   );
   gpc615_5 gpc74 (
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage0_4[78]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[13],stage1_5[27],stage1_4[74],stage1_3[74]}
   );
   gpc615_5 gpc75 (
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144]},
      {stage0_4[79]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[14],stage1_5[28],stage1_4[75],stage1_3[75]}
   );
   gpc615_5 gpc76 (
      {stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149]},
      {stage0_4[80]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[15],stage1_5[29],stage1_4[76],stage1_3[76]}
   );
   gpc615_5 gpc77 (
      {stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154]},
      {stage0_4[81]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[16],stage1_5[30],stage1_4[77],stage1_3[77]}
   );
   gpc615_5 gpc78 (
      {stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159]},
      {stage0_4[82]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[17],stage1_5[31],stage1_4[78],stage1_3[78]}
   );
   gpc615_5 gpc79 (
      {stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164]},
      {stage0_4[83]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[18],stage1_5[32],stage1_4[79],stage1_3[79]}
   );
   gpc615_5 gpc80 (
      {stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169]},
      {stage0_4[84]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[19],stage1_5[33],stage1_4[80],stage1_3[80]}
   );
   gpc615_5 gpc81 (
      {stage0_3[170], stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174]},
      {stage0_4[85]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[20],stage1_5[34],stage1_4[81],stage1_3[81]}
   );
   gpc615_5 gpc82 (
      {stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178], stage0_3[179]},
      {stage0_4[86]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[21],stage1_5[35],stage1_4[82],stage1_3[82]}
   );
   gpc615_5 gpc83 (
      {stage0_3[180], stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184]},
      {stage0_4[87]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[22],stage1_5[36],stage1_4[83],stage1_3[83]}
   );
   gpc615_5 gpc84 (
      {stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188], stage0_3[189]},
      {stage0_4[88]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[23],stage1_5[37],stage1_4[84],stage1_3[84]}
   );
   gpc615_5 gpc85 (
      {stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194]},
      {stage0_4[89]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[24],stage1_5[38],stage1_4[85],stage1_3[85]}
   );
   gpc615_5 gpc86 (
      {stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199]},
      {stage0_4[90]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[25],stage1_5[39],stage1_4[86],stage1_3[86]}
   );
   gpc615_5 gpc87 (
      {stage0_3[200], stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204]},
      {stage0_4[91]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[26],stage1_5[40],stage1_4[87],stage1_3[87]}
   );
   gpc615_5 gpc88 (
      {stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208], stage0_3[209]},
      {stage0_4[92]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[27],stage1_5[41],stage1_4[88],stage1_3[88]}
   );
   gpc615_5 gpc89 (
      {stage0_3[210], stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214]},
      {stage0_4[93]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[28],stage1_5[42],stage1_4[89],stage1_3[89]}
   );
   gpc615_5 gpc90 (
      {stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218], stage0_3[219]},
      {stage0_4[94]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[29],stage1_5[43],stage1_4[90],stage1_3[90]}
   );
   gpc615_5 gpc91 (
      {stage0_3[220], stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224]},
      {stage0_4[95]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[30],stage1_5[44],stage1_4[91],stage1_3[91]}
   );
   gpc615_5 gpc92 (
      {stage0_3[225], stage0_3[226], stage0_3[227], stage0_3[228], stage0_3[229]},
      {stage0_4[96]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[31],stage1_5[45],stage1_4[92],stage1_3[92]}
   );
   gpc615_5 gpc93 (
      {stage0_3[230], stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234]},
      {stage0_4[97]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[32],stage1_5[46],stage1_4[93],stage1_3[93]}
   );
   gpc615_5 gpc94 (
      {stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238], stage0_3[239]},
      {stage0_4[98]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[33],stage1_5[47],stage1_4[94],stage1_3[94]}
   );
   gpc615_5 gpc95 (
      {stage0_3[240], stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244]},
      {stage0_4[99]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[34],stage1_5[48],stage1_4[95],stage1_3[95]}
   );
   gpc606_5 gpc96 (
      {stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[22],stage1_6[35],stage1_5[49],stage1_4[96]}
   );
   gpc606_5 gpc97 (
      {stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[23],stage1_6[36],stage1_5[50],stage1_4[97]}
   );
   gpc606_5 gpc98 (
      {stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[24],stage1_6[37],stage1_5[51],stage1_4[98]}
   );
   gpc606_5 gpc99 (
      {stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[25],stage1_6[38],stage1_5[52],stage1_4[99]}
   );
   gpc606_5 gpc100 (
      {stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[26],stage1_6[39],stage1_5[53],stage1_4[100]}
   );
   gpc606_5 gpc101 (
      {stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[27],stage1_6[40],stage1_5[54],stage1_4[101]}
   );
   gpc606_5 gpc102 (
      {stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[28],stage1_6[41],stage1_5[55],stage1_4[102]}
   );
   gpc606_5 gpc103 (
      {stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[29],stage1_6[42],stage1_5[56],stage1_4[103]}
   );
   gpc606_5 gpc104 (
      {stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[30],stage1_6[43],stage1_5[57],stage1_4[104]}
   );
   gpc606_5 gpc105 (
      {stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[31],stage1_6[44],stage1_5[58],stage1_4[105]}
   );
   gpc606_5 gpc106 (
      {stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[32],stage1_6[45],stage1_5[59],stage1_4[106]}
   );
   gpc606_5 gpc107 (
      {stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[33],stage1_6[46],stage1_5[60],stage1_4[107]}
   );
   gpc606_5 gpc108 (
      {stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[34],stage1_6[47],stage1_5[61],stage1_4[108]}
   );
   gpc606_5 gpc109 (
      {stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[35],stage1_6[48],stage1_5[62],stage1_4[109]}
   );
   gpc606_5 gpc110 (
      {stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188], stage0_4[189]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[36],stage1_6[49],stage1_5[63],stage1_4[110]}
   );
   gpc606_5 gpc111 (
      {stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193], stage0_4[194], stage0_4[195]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[37],stage1_6[50],stage1_5[64],stage1_4[111]}
   );
   gpc606_5 gpc112 (
      {stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199], stage0_4[200], stage0_4[201]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[38],stage1_6[51],stage1_5[65],stage1_4[112]}
   );
   gpc606_5 gpc113 (
      {stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[39],stage1_6[52],stage1_5[66],stage1_4[113]}
   );
   gpc606_5 gpc114 (
      {stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[40],stage1_6[53],stage1_5[67],stage1_4[114]}
   );
   gpc606_5 gpc115 (
      {stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218], stage0_4[219]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[41],stage1_6[54],stage1_5[68],stage1_4[115]}
   );
   gpc606_5 gpc116 (
      {stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224], stage0_4[225]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[42],stage1_6[55],stage1_5[69],stage1_4[116]}
   );
   gpc606_5 gpc117 (
      {stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230], stage0_4[231]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[43],stage1_6[56],stage1_5[70],stage1_4[117]}
   );
   gpc606_5 gpc118 (
      {stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[44],stage1_6[57],stage1_5[71],stage1_4[118]}
   );
   gpc606_5 gpc119 (
      {stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[45],stage1_6[58],stage1_5[72],stage1_4[119]}
   );
   gpc606_5 gpc120 (
      {stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248], stage0_4[249]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[46],stage1_6[59],stage1_5[73],stage1_4[120]}
   );
   gpc606_5 gpc121 (
      {stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254], stage0_4[255]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[47],stage1_6[60],stage1_5[74],stage1_4[121]}
   );
   gpc606_5 gpc122 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[26],stage1_7[48],stage1_6[61],stage1_5[75]}
   );
   gpc606_5 gpc123 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[27],stage1_7[49],stage1_6[62],stage1_5[76]}
   );
   gpc606_5 gpc124 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[28],stage1_7[50],stage1_6[63],stage1_5[77]}
   );
   gpc606_5 gpc125 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[29],stage1_7[51],stage1_6[64],stage1_5[78]}
   );
   gpc606_5 gpc126 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[30],stage1_7[52],stage1_6[65],stage1_5[79]}
   );
   gpc606_5 gpc127 (
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[31],stage1_7[53],stage1_6[66],stage1_5[80]}
   );
   gpc606_5 gpc128 (
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[32],stage1_7[54],stage1_6[67],stage1_5[81]}
   );
   gpc606_5 gpc129 (
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[33],stage1_7[55],stage1_6[68],stage1_5[82]}
   );
   gpc606_5 gpc130 (
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[34],stage1_7[56],stage1_6[69],stage1_5[83]}
   );
   gpc606_5 gpc131 (
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[35],stage1_7[57],stage1_6[70],stage1_5[84]}
   );
   gpc606_5 gpc132 (
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[36],stage1_7[58],stage1_6[71],stage1_5[85]}
   );
   gpc606_5 gpc133 (
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[37],stage1_7[59],stage1_6[72],stage1_5[86]}
   );
   gpc606_5 gpc134 (
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[38],stage1_7[60],stage1_6[73],stage1_5[87]}
   );
   gpc606_5 gpc135 (
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[39],stage1_7[61],stage1_6[74],stage1_5[88]}
   );
   gpc606_5 gpc136 (
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[40],stage1_7[62],stage1_6[75],stage1_5[89]}
   );
   gpc606_5 gpc137 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[41],stage1_7[63],stage1_6[76],stage1_5[90]}
   );
   gpc606_5 gpc138 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[42],stage1_7[64],stage1_6[77],stage1_5[91]}
   );
   gpc606_5 gpc139 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[43],stage1_7[65],stage1_6[78],stage1_5[92]}
   );
   gpc606_5 gpc140 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[44],stage1_7[66],stage1_6[79],stage1_5[93]}
   );
   gpc606_5 gpc141 (
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[45],stage1_7[67],stage1_6[80],stage1_5[94]}
   );
   gpc606_5 gpc142 (
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], 1'b0, 1'b0},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[46],stage1_7[68],stage1_6[81],stage1_5[95]}
   );
   gpc1415_5 gpc143 (
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160]},
      {stage0_7[126]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3]},
      {stage0_9[0]},
      {stage1_10[0],stage1_9[21],stage1_8[47],stage1_7[69],stage1_6[82]}
   );
   gpc606_5 gpc144 (
      {stage0_6[161], stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166]},
      {stage0_8[4], stage0_8[5], stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9]},
      {stage1_10[1],stage1_9[22],stage1_8[48],stage1_7[70],stage1_6[83]}
   );
   gpc606_5 gpc145 (
      {stage0_6[167], stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172]},
      {stage0_8[10], stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage1_10[2],stage1_9[23],stage1_8[49],stage1_7[71],stage1_6[84]}
   );
   gpc606_5 gpc146 (
      {stage0_6[173], stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178]},
      {stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21]},
      {stage1_10[3],stage1_9[24],stage1_8[50],stage1_7[72],stage1_6[85]}
   );
   gpc606_5 gpc147 (
      {stage0_6[179], stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184]},
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage1_10[4],stage1_9[25],stage1_8[51],stage1_7[73],stage1_6[86]}
   );
   gpc606_5 gpc148 (
      {stage0_6[185], stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190]},
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage1_10[5],stage1_9[26],stage1_8[52],stage1_7[74],stage1_6[87]}
   );
   gpc606_5 gpc149 (
      {stage0_6[191], stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196]},
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39]},
      {stage1_10[6],stage1_9[27],stage1_8[53],stage1_7[75],stage1_6[88]}
   );
   gpc606_5 gpc150 (
      {stage0_6[197], stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202]},
      {stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45]},
      {stage1_10[7],stage1_9[28],stage1_8[54],stage1_7[76],stage1_6[89]}
   );
   gpc606_5 gpc151 (
      {stage0_6[203], stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208]},
      {stage0_8[46], stage0_8[47], stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51]},
      {stage1_10[8],stage1_9[29],stage1_8[55],stage1_7[77],stage1_6[90]}
   );
   gpc606_5 gpc152 (
      {stage0_6[209], stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214]},
      {stage0_8[52], stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57]},
      {stage1_10[9],stage1_9[30],stage1_8[56],stage1_7[78],stage1_6[91]}
   );
   gpc606_5 gpc153 (
      {stage0_6[215], stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220]},
      {stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63]},
      {stage1_10[10],stage1_9[31],stage1_8[57],stage1_7[79],stage1_6[92]}
   );
   gpc615_5 gpc154 (
      {stage0_6[221], stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225]},
      {stage0_7[127]},
      {stage0_8[64], stage0_8[65], stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69]},
      {stage1_10[11],stage1_9[32],stage1_8[58],stage1_7[80],stage1_6[93]}
   );
   gpc615_5 gpc155 (
      {stage0_6[226], stage0_6[227], stage0_6[228], stage0_6[229], stage0_6[230]},
      {stage0_7[128]},
      {stage0_8[70], stage0_8[71], stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75]},
      {stage1_10[12],stage1_9[33],stage1_8[59],stage1_7[81],stage1_6[94]}
   );
   gpc615_5 gpc156 (
      {stage0_6[231], stage0_6[232], stage0_6[233], stage0_6[234], stage0_6[235]},
      {stage0_7[129]},
      {stage0_8[76], stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81]},
      {stage1_10[13],stage1_9[34],stage1_8[60],stage1_7[82],stage1_6[95]}
   );
   gpc606_5 gpc157 (
      {stage0_7[130], stage0_7[131], stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135]},
      {stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6]},
      {stage1_11[0],stage1_10[14],stage1_9[35],stage1_8[61],stage1_7[83]}
   );
   gpc606_5 gpc158 (
      {stage0_7[136], stage0_7[137], stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141]},
      {stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12]},
      {stage1_11[1],stage1_10[15],stage1_9[36],stage1_8[62],stage1_7[84]}
   );
   gpc606_5 gpc159 (
      {stage0_7[142], stage0_7[143], stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147]},
      {stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18]},
      {stage1_11[2],stage1_10[16],stage1_9[37],stage1_8[63],stage1_7[85]}
   );
   gpc606_5 gpc160 (
      {stage0_7[148], stage0_7[149], stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153]},
      {stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24]},
      {stage1_11[3],stage1_10[17],stage1_9[38],stage1_8[64],stage1_7[86]}
   );
   gpc606_5 gpc161 (
      {stage0_7[154], stage0_7[155], stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159]},
      {stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30]},
      {stage1_11[4],stage1_10[18],stage1_9[39],stage1_8[65],stage1_7[87]}
   );
   gpc606_5 gpc162 (
      {stage0_7[160], stage0_7[161], stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165]},
      {stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36]},
      {stage1_11[5],stage1_10[19],stage1_9[40],stage1_8[66],stage1_7[88]}
   );
   gpc606_5 gpc163 (
      {stage0_7[166], stage0_7[167], stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171]},
      {stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42]},
      {stage1_11[6],stage1_10[20],stage1_9[41],stage1_8[67],stage1_7[89]}
   );
   gpc606_5 gpc164 (
      {stage0_7[172], stage0_7[173], stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177]},
      {stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48]},
      {stage1_11[7],stage1_10[21],stage1_9[42],stage1_8[68],stage1_7[90]}
   );
   gpc606_5 gpc165 (
      {stage0_7[178], stage0_7[179], stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183]},
      {stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53], stage0_9[54]},
      {stage1_11[8],stage1_10[22],stage1_9[43],stage1_8[69],stage1_7[91]}
   );
   gpc606_5 gpc166 (
      {stage0_7[184], stage0_7[185], stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189]},
      {stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59], stage0_9[60]},
      {stage1_11[9],stage1_10[23],stage1_9[44],stage1_8[70],stage1_7[92]}
   );
   gpc606_5 gpc167 (
      {stage0_7[190], stage0_7[191], stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195]},
      {stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65], stage0_9[66]},
      {stage1_11[10],stage1_10[24],stage1_9[45],stage1_8[71],stage1_7[93]}
   );
   gpc615_5 gpc168 (
      {stage0_7[196], stage0_7[197], stage0_7[198], stage0_7[199], stage0_7[200]},
      {stage0_8[82]},
      {stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71], stage0_9[72]},
      {stage1_11[11],stage1_10[25],stage1_9[46],stage1_8[72],stage1_7[94]}
   );
   gpc615_5 gpc169 (
      {stage0_7[201], stage0_7[202], stage0_7[203], stage0_7[204], stage0_7[205]},
      {stage0_8[83]},
      {stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77], stage0_9[78]},
      {stage1_11[12],stage1_10[26],stage1_9[47],stage1_8[73],stage1_7[95]}
   );
   gpc615_5 gpc170 (
      {stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209], stage0_7[210]},
      {stage0_8[84]},
      {stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84]},
      {stage1_11[13],stage1_10[27],stage1_9[48],stage1_8[74],stage1_7[96]}
   );
   gpc615_5 gpc171 (
      {stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage0_8[85]},
      {stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90]},
      {stage1_11[14],stage1_10[28],stage1_9[49],stage1_8[75],stage1_7[97]}
   );
   gpc615_5 gpc172 (
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220]},
      {stage0_8[86]},
      {stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96]},
      {stage1_11[15],stage1_10[29],stage1_9[50],stage1_8[76],stage1_7[98]}
   );
   gpc615_5 gpc173 (
      {stage0_7[221], stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225]},
      {stage0_8[87]},
      {stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102]},
      {stage1_11[16],stage1_10[30],stage1_9[51],stage1_8[77],stage1_7[99]}
   );
   gpc615_5 gpc174 (
      {stage0_7[226], stage0_7[227], stage0_7[228], stage0_7[229], stage0_7[230]},
      {stage0_8[88]},
      {stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107], stage0_9[108]},
      {stage1_11[17],stage1_10[31],stage1_9[52],stage1_8[78],stage1_7[100]}
   );
   gpc615_5 gpc175 (
      {stage0_7[231], stage0_7[232], stage0_7[233], stage0_7[234], stage0_7[235]},
      {stage0_8[89]},
      {stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114]},
      {stage1_11[18],stage1_10[32],stage1_9[53],stage1_8[79],stage1_7[101]}
   );
   gpc615_5 gpc176 (
      {stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239], stage0_7[240]},
      {stage0_8[90]},
      {stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120]},
      {stage1_11[19],stage1_10[33],stage1_9[54],stage1_8[80],stage1_7[102]}
   );
   gpc615_5 gpc177 (
      {stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage0_8[91]},
      {stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126]},
      {stage1_11[20],stage1_10[34],stage1_9[55],stage1_8[81],stage1_7[103]}
   );
   gpc615_5 gpc178 (
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250]},
      {stage0_8[92]},
      {stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131], stage0_9[132]},
      {stage1_11[21],stage1_10[35],stage1_9[56],stage1_8[82],stage1_7[104]}
   );
   gpc606_5 gpc179 (
      {stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97], stage0_8[98]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[22],stage1_10[36],stage1_9[57],stage1_8[83]}
   );
   gpc606_5 gpc180 (
      {stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103], stage0_8[104]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[23],stage1_10[37],stage1_9[58],stage1_8[84]}
   );
   gpc606_5 gpc181 (
      {stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[24],stage1_10[38],stage1_9[59],stage1_8[85]}
   );
   gpc606_5 gpc182 (
      {stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[25],stage1_10[39],stage1_9[60],stage1_8[86]}
   );
   gpc606_5 gpc183 (
      {stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[26],stage1_10[40],stage1_9[61],stage1_8[87]}
   );
   gpc606_5 gpc184 (
      {stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127], stage0_8[128]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[27],stage1_10[41],stage1_9[62],stage1_8[88]}
   );
   gpc606_5 gpc185 (
      {stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132], stage0_8[133], stage0_8[134]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[28],stage1_10[42],stage1_9[63],stage1_8[89]}
   );
   gpc606_5 gpc186 (
      {stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[29],stage1_10[43],stage1_9[64],stage1_8[90]}
   );
   gpc606_5 gpc187 (
      {stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[30],stage1_10[44],stage1_9[65],stage1_8[91]}
   );
   gpc606_5 gpc188 (
      {stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150], stage0_8[151], stage0_8[152]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[31],stage1_10[45],stage1_9[66],stage1_8[92]}
   );
   gpc615_5 gpc189 (
      {stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156], stage0_8[157]},
      {stage0_9[133]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[32],stage1_10[46],stage1_9[67],stage1_8[93]}
   );
   gpc615_5 gpc190 (
      {stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162]},
      {stage0_9[134]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[33],stage1_10[47],stage1_9[68],stage1_8[94]}
   );
   gpc615_5 gpc191 (
      {stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage0_9[135]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[34],stage1_10[48],stage1_9[69],stage1_8[95]}
   );
   gpc615_5 gpc192 (
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172]},
      {stage0_9[136]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[35],stage1_10[49],stage1_9[70],stage1_8[96]}
   );
   gpc615_5 gpc193 (
      {stage0_8[173], stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177]},
      {stage0_9[137]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[36],stage1_10[50],stage1_9[71],stage1_8[97]}
   );
   gpc615_5 gpc194 (
      {stage0_8[178], stage0_8[179], stage0_8[180], stage0_8[181], stage0_8[182]},
      {stage0_9[138]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[37],stage1_10[51],stage1_9[72],stage1_8[98]}
   );
   gpc615_5 gpc195 (
      {stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186], stage0_8[187]},
      {stage0_9[139]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[38],stage1_10[52],stage1_9[73],stage1_8[99]}
   );
   gpc615_5 gpc196 (
      {stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192]},
      {stage0_9[140]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[39],stage1_10[53],stage1_9[74],stage1_8[100]}
   );
   gpc615_5 gpc197 (
      {stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage0_9[141]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[40],stage1_10[54],stage1_9[75],stage1_8[101]}
   );
   gpc615_5 gpc198 (
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202]},
      {stage0_9[142]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[41],stage1_10[55],stage1_9[76],stage1_8[102]}
   );
   gpc615_5 gpc199 (
      {stage0_8[203], stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207]},
      {stage0_9[143]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[42],stage1_10[56],stage1_9[77],stage1_8[103]}
   );
   gpc615_5 gpc200 (
      {stage0_8[208], stage0_8[209], stage0_8[210], stage0_8[211], stage0_8[212]},
      {stage0_9[144]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[43],stage1_10[57],stage1_9[78],stage1_8[104]}
   );
   gpc615_5 gpc201 (
      {stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216], stage0_8[217]},
      {stage0_9[145]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[44],stage1_10[58],stage1_9[79],stage1_8[105]}
   );
   gpc615_5 gpc202 (
      {stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222]},
      {stage0_9[146]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[45],stage1_10[59],stage1_9[80],stage1_8[106]}
   );
   gpc615_5 gpc203 (
      {stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227]},
      {stage0_9[147]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[46],stage1_10[60],stage1_9[81],stage1_8[107]}
   );
   gpc615_5 gpc204 (
      {stage0_8[228], stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232]},
      {stage0_9[148]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[47],stage1_10[61],stage1_9[82],stage1_8[108]}
   );
   gpc606_5 gpc205 (
      {stage0_9[149], stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[26],stage1_11[48],stage1_10[62],stage1_9[83]}
   );
   gpc606_5 gpc206 (
      {stage0_9[155], stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[27],stage1_11[49],stage1_10[63],stage1_9[84]}
   );
   gpc606_5 gpc207 (
      {stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[28],stage1_11[50],stage1_10[64],stage1_9[85]}
   );
   gpc606_5 gpc208 (
      {stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[29],stage1_11[51],stage1_10[65],stage1_9[86]}
   );
   gpc606_5 gpc209 (
      {stage0_9[173], stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[30],stage1_11[52],stage1_10[66],stage1_9[87]}
   );
   gpc606_5 gpc210 (
      {stage0_9[179], stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[31],stage1_11[53],stage1_10[67],stage1_9[88]}
   );
   gpc615_5 gpc211 (
      {stage0_9[185], stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189]},
      {stage0_10[156]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[32],stage1_11[54],stage1_10[68],stage1_9[89]}
   );
   gpc615_5 gpc212 (
      {stage0_9[190], stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194]},
      {stage0_10[157]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[33],stage1_11[55],stage1_10[69],stage1_9[90]}
   );
   gpc615_5 gpc213 (
      {stage0_9[195], stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199]},
      {stage0_10[158]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[34],stage1_11[56],stage1_10[70],stage1_9[91]}
   );
   gpc615_5 gpc214 (
      {stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204]},
      {stage0_10[159]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[35],stage1_11[57],stage1_10[71],stage1_9[92]}
   );
   gpc615_5 gpc215 (
      {stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_10[160]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[36],stage1_11[58],stage1_10[72],stage1_9[93]}
   );
   gpc615_5 gpc216 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214]},
      {stage0_10[161]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[37],stage1_11[59],stage1_10[73],stage1_9[94]}
   );
   gpc615_5 gpc217 (
      {stage0_9[215], stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219]},
      {stage0_10[162]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[38],stage1_11[60],stage1_10[74],stage1_9[95]}
   );
   gpc615_5 gpc218 (
      {stage0_9[220], stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224]},
      {stage0_10[163]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[39],stage1_11[61],stage1_10[75],stage1_9[96]}
   );
   gpc615_5 gpc219 (
      {stage0_9[225], stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229]},
      {stage0_10[164]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[40],stage1_11[62],stage1_10[76],stage1_9[97]}
   );
   gpc615_5 gpc220 (
      {stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234]},
      {stage0_10[165]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[41],stage1_11[63],stage1_10[77],stage1_9[98]}
   );
   gpc615_5 gpc221 (
      {stage0_10[166], stage0_10[167], stage0_10[168], stage0_10[169], stage0_10[170]},
      {stage0_11[96]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[16],stage1_12[42],stage1_11[64],stage1_10[78]}
   );
   gpc615_5 gpc222 (
      {stage0_10[171], stage0_10[172], stage0_10[173], stage0_10[174], stage0_10[175]},
      {stage0_11[97]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[17],stage1_12[43],stage1_11[65],stage1_10[79]}
   );
   gpc615_5 gpc223 (
      {stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179], stage0_10[180]},
      {stage0_11[98]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[18],stage1_12[44],stage1_11[66],stage1_10[80]}
   );
   gpc606_5 gpc224 (
      {stage0_11[99], stage0_11[100], stage0_11[101], stage0_11[102], stage0_11[103], stage0_11[104]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[3],stage1_13[19],stage1_12[45],stage1_11[67]}
   );
   gpc606_5 gpc225 (
      {stage0_11[105], stage0_11[106], stage0_11[107], stage0_11[108], stage0_11[109], stage0_11[110]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[4],stage1_13[20],stage1_12[46],stage1_11[68]}
   );
   gpc606_5 gpc226 (
      {stage0_11[111], stage0_11[112], stage0_11[113], stage0_11[114], stage0_11[115], stage0_11[116]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[5],stage1_13[21],stage1_12[47],stage1_11[69]}
   );
   gpc606_5 gpc227 (
      {stage0_11[117], stage0_11[118], stage0_11[119], stage0_11[120], stage0_11[121], stage0_11[122]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[6],stage1_13[22],stage1_12[48],stage1_11[70]}
   );
   gpc606_5 gpc228 (
      {stage0_11[123], stage0_11[124], stage0_11[125], stage0_11[126], stage0_11[127], stage0_11[128]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[7],stage1_13[23],stage1_12[49],stage1_11[71]}
   );
   gpc606_5 gpc229 (
      {stage0_11[129], stage0_11[130], stage0_11[131], stage0_11[132], stage0_11[133], stage0_11[134]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[8],stage1_13[24],stage1_12[50],stage1_11[72]}
   );
   gpc606_5 gpc230 (
      {stage0_11[135], stage0_11[136], stage0_11[137], stage0_11[138], stage0_11[139], stage0_11[140]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[9],stage1_13[25],stage1_12[51],stage1_11[73]}
   );
   gpc606_5 gpc231 (
      {stage0_11[141], stage0_11[142], stage0_11[143], stage0_11[144], stage0_11[145], stage0_11[146]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[10],stage1_13[26],stage1_12[52],stage1_11[74]}
   );
   gpc606_5 gpc232 (
      {stage0_11[147], stage0_11[148], stage0_11[149], stage0_11[150], stage0_11[151], stage0_11[152]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[11],stage1_13[27],stage1_12[53],stage1_11[75]}
   );
   gpc606_5 gpc233 (
      {stage0_11[153], stage0_11[154], stage0_11[155], stage0_11[156], stage0_11[157], stage0_11[158]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[12],stage1_13[28],stage1_12[54],stage1_11[76]}
   );
   gpc606_5 gpc234 (
      {stage0_11[159], stage0_11[160], stage0_11[161], stage0_11[162], stage0_11[163], stage0_11[164]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[13],stage1_13[29],stage1_12[55],stage1_11[77]}
   );
   gpc606_5 gpc235 (
      {stage0_11[165], stage0_11[166], stage0_11[167], stage0_11[168], stage0_11[169], stage0_11[170]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[14],stage1_13[30],stage1_12[56],stage1_11[78]}
   );
   gpc606_5 gpc236 (
      {stage0_11[171], stage0_11[172], stage0_11[173], stage0_11[174], stage0_11[175], stage0_11[176]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[15],stage1_13[31],stage1_12[57],stage1_11[79]}
   );
   gpc606_5 gpc237 (
      {stage0_11[177], stage0_11[178], stage0_11[179], stage0_11[180], stage0_11[181], stage0_11[182]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[16],stage1_13[32],stage1_12[58],stage1_11[80]}
   );
   gpc606_5 gpc238 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[14],stage1_14[17],stage1_13[33],stage1_12[59]}
   );
   gpc606_5 gpc239 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[15],stage1_14[18],stage1_13[34],stage1_12[60]}
   );
   gpc606_5 gpc240 (
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[16],stage1_14[19],stage1_13[35],stage1_12[61]}
   );
   gpc606_5 gpc241 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[17],stage1_14[20],stage1_13[36],stage1_12[62]}
   );
   gpc606_5 gpc242 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[18],stage1_14[21],stage1_13[37],stage1_12[63]}
   );
   gpc606_5 gpc243 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[19],stage1_14[22],stage1_13[38],stage1_12[64]}
   );
   gpc606_5 gpc244 (
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[20],stage1_14[23],stage1_13[39],stage1_12[65]}
   );
   gpc606_5 gpc245 (
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[21],stage1_14[24],stage1_13[40],stage1_12[66]}
   );
   gpc606_5 gpc246 (
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[22],stage1_14[25],stage1_13[41],stage1_12[67]}
   );
   gpc606_5 gpc247 (
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[23],stage1_14[26],stage1_13[42],stage1_12[68]}
   );
   gpc606_5 gpc248 (
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[24],stage1_14[27],stage1_13[43],stage1_12[69]}
   );
   gpc606_5 gpc249 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[25],stage1_14[28],stage1_13[44],stage1_12[70]}
   );
   gpc615_5 gpc250 (
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94]},
      {stage0_13[84]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[26],stage1_14[29],stage1_13[45],stage1_12[71]}
   );
   gpc615_5 gpc251 (
      {stage0_12[95], stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99]},
      {stage0_13[85]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[27],stage1_14[30],stage1_13[46],stage1_12[72]}
   );
   gpc615_5 gpc252 (
      {stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103], stage0_12[104]},
      {stage0_13[86]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[28],stage1_14[31],stage1_13[47],stage1_12[73]}
   );
   gpc615_5 gpc253 (
      {stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109]},
      {stage0_13[87]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[29],stage1_14[32],stage1_13[48],stage1_12[74]}
   );
   gpc615_5 gpc254 (
      {stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114]},
      {stage0_13[88]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[30],stage1_14[33],stage1_13[49],stage1_12[75]}
   );
   gpc615_5 gpc255 (
      {stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage0_13[89]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[31],stage1_14[34],stage1_13[50],stage1_12[76]}
   );
   gpc615_5 gpc256 (
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124]},
      {stage0_13[90]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[32],stage1_14[35],stage1_13[51],stage1_12[77]}
   );
   gpc615_5 gpc257 (
      {stage0_12[125], stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129]},
      {stage0_13[91]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[33],stage1_14[36],stage1_13[52],stage1_12[78]}
   );
   gpc615_5 gpc258 (
      {stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133], stage0_12[134]},
      {stage0_13[92]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[34],stage1_14[37],stage1_13[53],stage1_12[79]}
   );
   gpc615_5 gpc259 (
      {stage0_12[135], stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139]},
      {stage0_13[93]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[35],stage1_14[38],stage1_13[54],stage1_12[80]}
   );
   gpc615_5 gpc260 (
      {stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143], stage0_12[144]},
      {stage0_13[94]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[36],stage1_14[39],stage1_13[55],stage1_12[81]}
   );
   gpc615_5 gpc261 (
      {stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage0_13[95]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[37],stage1_14[40],stage1_13[56],stage1_12[82]}
   );
   gpc615_5 gpc262 (
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154]},
      {stage0_13[96]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[38],stage1_14[41],stage1_13[57],stage1_12[83]}
   );
   gpc615_5 gpc263 (
      {stage0_12[155], stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159]},
      {stage0_13[97]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[39],stage1_14[42],stage1_13[58],stage1_12[84]}
   );
   gpc615_5 gpc264 (
      {stage0_12[160], stage0_12[161], stage0_12[162], stage0_12[163], stage0_12[164]},
      {stage0_13[98]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[40],stage1_14[43],stage1_13[59],stage1_12[85]}
   );
   gpc615_5 gpc265 (
      {stage0_12[165], stage0_12[166], stage0_12[167], stage0_12[168], stage0_12[169]},
      {stage0_13[99]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[41],stage1_14[44],stage1_13[60],stage1_12[86]}
   );
   gpc615_5 gpc266 (
      {stage0_12[170], stage0_12[171], stage0_12[172], stage0_12[173], stage0_12[174]},
      {stage0_13[100]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[42],stage1_14[45],stage1_13[61],stage1_12[87]}
   );
   gpc615_5 gpc267 (
      {stage0_12[175], stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179]},
      {stage0_13[101]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[43],stage1_14[46],stage1_13[62],stage1_12[88]}
   );
   gpc615_5 gpc268 (
      {stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183], stage0_12[184]},
      {stage0_13[102]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[44],stage1_14[47],stage1_13[63],stage1_12[89]}
   );
   gpc615_5 gpc269 (
      {stage0_12[185], stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189]},
      {stage0_13[103]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[45],stage1_14[48],stage1_13[64],stage1_12[90]}
   );
   gpc615_5 gpc270 (
      {stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193], stage0_12[194]},
      {stage0_13[104]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[46],stage1_14[49],stage1_13[65],stage1_12[91]}
   );
   gpc615_5 gpc271 (
      {stage0_12[195], stage0_12[196], stage0_12[197], stage0_12[198], stage0_12[199]},
      {stage0_13[105]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[47],stage1_14[50],stage1_13[66],stage1_12[92]}
   );
   gpc615_5 gpc272 (
      {stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203], stage0_12[204]},
      {stage0_13[106]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[48],stage1_14[51],stage1_13[67],stage1_12[93]}
   );
   gpc615_5 gpc273 (
      {stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209]},
      {stage0_13[107]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[49],stage1_14[52],stage1_13[68],stage1_12[94]}
   );
   gpc615_5 gpc274 (
      {stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213], stage0_12[214]},
      {stage0_13[108]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[50],stage1_14[53],stage1_13[69],stage1_12[95]}
   );
   gpc615_5 gpc275 (
      {stage0_12[215], stage0_12[216], stage0_12[217], stage0_12[218], stage0_12[219]},
      {stage0_13[109]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[51],stage1_14[54],stage1_13[70],stage1_12[96]}
   );
   gpc606_5 gpc276 (
      {stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113], stage0_13[114], stage0_13[115]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[38],stage1_15[52],stage1_14[55],stage1_13[71]}
   );
   gpc606_5 gpc277 (
      {stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119], stage0_13[120], stage0_13[121]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[39],stage1_15[53],stage1_14[56],stage1_13[72]}
   );
   gpc606_5 gpc278 (
      {stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125], stage0_13[126], stage0_13[127]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[40],stage1_15[54],stage1_14[57],stage1_13[73]}
   );
   gpc606_5 gpc279 (
      {stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131], stage0_13[132], stage0_13[133]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[41],stage1_15[55],stage1_14[58],stage1_13[74]}
   );
   gpc606_5 gpc280 (
      {stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137], stage0_13[138], stage0_13[139]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[42],stage1_15[56],stage1_14[59],stage1_13[75]}
   );
   gpc606_5 gpc281 (
      {stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143], stage0_13[144], stage0_13[145]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[43],stage1_15[57],stage1_14[60],stage1_13[76]}
   );
   gpc606_5 gpc282 (
      {stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149], stage0_13[150], stage0_13[151]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[44],stage1_15[58],stage1_14[61],stage1_13[77]}
   );
   gpc606_5 gpc283 (
      {stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155], stage0_13[156], stage0_13[157]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[45],stage1_15[59],stage1_14[62],stage1_13[78]}
   );
   gpc606_5 gpc284 (
      {stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161], stage0_13[162], stage0_13[163]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[46],stage1_15[60],stage1_14[63],stage1_13[79]}
   );
   gpc606_5 gpc285 (
      {stage0_13[164], stage0_13[165], stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[47],stage1_15[61],stage1_14[64],stage1_13[80]}
   );
   gpc606_5 gpc286 (
      {stage0_13[170], stage0_13[171], stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[48],stage1_15[62],stage1_14[65],stage1_13[81]}
   );
   gpc606_5 gpc287 (
      {stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[49],stage1_15[63],stage1_14[66],stage1_13[82]}
   );
   gpc606_5 gpc288 (
      {stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185], stage0_13[186], stage0_13[187]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[50],stage1_15[64],stage1_14[67],stage1_13[83]}
   );
   gpc606_5 gpc289 (
      {stage0_13[188], stage0_13[189], stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[51],stage1_15[65],stage1_14[68],stage1_13[84]}
   );
   gpc606_5 gpc290 (
      {stage0_13[194], stage0_13[195], stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[52],stage1_15[66],stage1_14[69],stage1_13[85]}
   );
   gpc606_5 gpc291 (
      {stage0_13[200], stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[53],stage1_15[67],stage1_14[70],stage1_13[86]}
   );
   gpc606_5 gpc292 (
      {stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210], stage0_13[211]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[54],stage1_15[68],stage1_14[71],stage1_13[87]}
   );
   gpc606_5 gpc293 (
      {stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215], stage0_13[216], stage0_13[217]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[55],stage1_15[69],stage1_14[72],stage1_13[88]}
   );
   gpc606_5 gpc294 (
      {stage0_13[218], stage0_13[219], stage0_13[220], stage0_13[221], stage0_13[222], stage0_13[223]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[56],stage1_15[70],stage1_14[73],stage1_13[89]}
   );
   gpc606_5 gpc295 (
      {stage0_13[224], stage0_13[225], stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[57],stage1_15[71],stage1_14[74],stage1_13[90]}
   );
   gpc606_5 gpc296 (
      {stage0_13[230], stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[58],stage1_15[72],stage1_14[75],stage1_13[91]}
   );
   gpc606_5 gpc297 (
      {stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240], stage0_13[241]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[59],stage1_15[73],stage1_14[76],stage1_13[92]}
   );
   gpc606_5 gpc298 (
      {stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245], stage0_13[246], stage0_13[247]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[60],stage1_15[74],stage1_14[77],stage1_13[93]}
   );
   gpc606_5 gpc299 (
      {stage0_13[248], stage0_13[249], stage0_13[250], stage0_13[251], stage0_13[252], stage0_13[253]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[61],stage1_15[75],stage1_14[78],stage1_13[94]}
   );
   gpc615_5 gpc300 (
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232]},
      {stage0_15[144]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[24],stage1_16[62],stage1_15[76],stage1_14[79]}
   );
   gpc615_5 gpc301 (
      {stage0_14[233], stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237]},
      {stage0_15[145]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[25],stage1_16[63],stage1_15[77],stage1_14[80]}
   );
   gpc615_5 gpc302 (
      {stage0_14[238], stage0_14[239], stage0_14[240], stage0_14[241], stage0_14[242]},
      {stage0_15[146]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[26],stage1_16[64],stage1_15[78],stage1_14[81]}
   );
   gpc615_5 gpc303 (
      {stage0_14[243], stage0_14[244], stage0_14[245], stage0_14[246], stage0_14[247]},
      {stage0_15[147]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[27],stage1_16[65],stage1_15[79],stage1_14[82]}
   );
   gpc615_5 gpc304 (
      {stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251], stage0_14[252]},
      {stage0_15[148]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[28],stage1_16[66],stage1_15[80],stage1_14[83]}
   );
   gpc615_5 gpc305 (
      {stage0_14[253], stage0_14[254], stage0_14[255], 1'b0, 1'b0},
      {stage0_15[149]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[29],stage1_16[67],stage1_15[81],stage1_14[84]}
   );
   gpc615_5 gpc306 (
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154]},
      {stage0_16[36]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[6],stage1_17[30],stage1_16[68],stage1_15[82]}
   );
   gpc615_5 gpc307 (
      {stage0_15[155], stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159]},
      {stage0_16[37]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[7],stage1_17[31],stage1_16[69],stage1_15[83]}
   );
   gpc615_5 gpc308 (
      {stage0_15[160], stage0_15[161], stage0_15[162], stage0_15[163], stage0_15[164]},
      {stage0_16[38]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[8],stage1_17[32],stage1_16[70],stage1_15[84]}
   );
   gpc615_5 gpc309 (
      {stage0_15[165], stage0_15[166], stage0_15[167], stage0_15[168], stage0_15[169]},
      {stage0_16[39]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[9],stage1_17[33],stage1_16[71],stage1_15[85]}
   );
   gpc615_5 gpc310 (
      {stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173], stage0_15[174]},
      {stage0_16[40]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[10],stage1_17[34],stage1_16[72],stage1_15[86]}
   );
   gpc615_5 gpc311 (
      {stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage0_16[41]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[11],stage1_17[35],stage1_16[73],stage1_15[87]}
   );
   gpc615_5 gpc312 (
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184]},
      {stage0_16[42]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[12],stage1_17[36],stage1_16[74],stage1_15[88]}
   );
   gpc615_5 gpc313 (
      {stage0_15[185], stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189]},
      {stage0_16[43]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[13],stage1_17[37],stage1_16[75],stage1_15[89]}
   );
   gpc615_5 gpc314 (
      {stage0_15[190], stage0_15[191], stage0_15[192], stage0_15[193], stage0_15[194]},
      {stage0_16[44]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[14],stage1_17[38],stage1_16[76],stage1_15[90]}
   );
   gpc615_5 gpc315 (
      {stage0_15[195], stage0_15[196], stage0_15[197], stage0_15[198], stage0_15[199]},
      {stage0_16[45]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[15],stage1_17[39],stage1_16[77],stage1_15[91]}
   );
   gpc615_5 gpc316 (
      {stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203], stage0_15[204]},
      {stage0_16[46]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[16],stage1_17[40],stage1_16[78],stage1_15[92]}
   );
   gpc615_5 gpc317 (
      {stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage0_16[47]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[17],stage1_17[41],stage1_16[79],stage1_15[93]}
   );
   gpc615_5 gpc318 (
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214]},
      {stage0_16[48]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[18],stage1_17[42],stage1_16[80],stage1_15[94]}
   );
   gpc615_5 gpc319 (
      {stage0_15[215], stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219]},
      {stage0_16[49]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[19],stage1_17[43],stage1_16[81],stage1_15[95]}
   );
   gpc606_5 gpc320 (
      {stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53], stage0_16[54], stage0_16[55]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[14],stage1_18[20],stage1_17[44],stage1_16[82]}
   );
   gpc606_5 gpc321 (
      {stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59], stage0_16[60], stage0_16[61]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[15],stage1_18[21],stage1_17[45],stage1_16[83]}
   );
   gpc606_5 gpc322 (
      {stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65], stage0_16[66], stage0_16[67]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[16],stage1_18[22],stage1_17[46],stage1_16[84]}
   );
   gpc606_5 gpc323 (
      {stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71], stage0_16[72], stage0_16[73]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[17],stage1_18[23],stage1_17[47],stage1_16[85]}
   );
   gpc606_5 gpc324 (
      {stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77], stage0_16[78], stage0_16[79]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[18],stage1_18[24],stage1_17[48],stage1_16[86]}
   );
   gpc606_5 gpc325 (
      {stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83], stage0_16[84], stage0_16[85]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[19],stage1_18[25],stage1_17[49],stage1_16[87]}
   );
   gpc606_5 gpc326 (
      {stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90], stage0_16[91]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[20],stage1_18[26],stage1_17[50],stage1_16[88]}
   );
   gpc606_5 gpc327 (
      {stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96], stage0_16[97]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[21],stage1_18[27],stage1_17[51],stage1_16[89]}
   );
   gpc606_5 gpc328 (
      {stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102], stage0_16[103]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[22],stage1_18[28],stage1_17[52],stage1_16[90]}
   );
   gpc606_5 gpc329 (
      {stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108], stage0_16[109]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[23],stage1_18[29],stage1_17[53],stage1_16[91]}
   );
   gpc606_5 gpc330 (
      {stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113], stage0_16[114], stage0_16[115]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[24],stage1_18[30],stage1_17[54],stage1_16[92]}
   );
   gpc606_5 gpc331 (
      {stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119], stage0_16[120], stage0_16[121]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[25],stage1_18[31],stage1_17[55],stage1_16[93]}
   );
   gpc606_5 gpc332 (
      {stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126], stage0_16[127]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[26],stage1_18[32],stage1_17[56],stage1_16[94]}
   );
   gpc606_5 gpc333 (
      {stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132], stage0_16[133]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[27],stage1_18[33],stage1_17[57],stage1_16[95]}
   );
   gpc606_5 gpc334 (
      {stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138], stage0_16[139]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[28],stage1_18[34],stage1_17[58],stage1_16[96]}
   );
   gpc606_5 gpc335 (
      {stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144], stage0_16[145]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[29],stage1_18[35],stage1_17[59],stage1_16[97]}
   );
   gpc606_5 gpc336 (
      {stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[30],stage1_18[36],stage1_17[60],stage1_16[98]}
   );
   gpc606_5 gpc337 (
      {stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[31],stage1_18[37],stage1_17[61],stage1_16[99]}
   );
   gpc606_5 gpc338 (
      {stage0_16[158], stage0_16[159], stage0_16[160], stage0_16[161], stage0_16[162], stage0_16[163]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[32],stage1_18[38],stage1_17[62],stage1_16[100]}
   );
   gpc606_5 gpc339 (
      {stage0_16[164], stage0_16[165], stage0_16[166], stage0_16[167], stage0_16[168], stage0_16[169]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[33],stage1_18[39],stage1_17[63],stage1_16[101]}
   );
   gpc615_5 gpc340 (
      {stage0_16[170], stage0_16[171], stage0_16[172], stage0_16[173], stage0_16[174]},
      {stage0_17[84]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[34],stage1_18[40],stage1_17[64],stage1_16[102]}
   );
   gpc615_5 gpc341 (
      {stage0_16[175], stage0_16[176], stage0_16[177], stage0_16[178], stage0_16[179]},
      {stage0_17[85]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[35],stage1_18[41],stage1_17[65],stage1_16[103]}
   );
   gpc615_5 gpc342 (
      {stage0_16[180], stage0_16[181], stage0_16[182], stage0_16[183], stage0_16[184]},
      {stage0_17[86]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[36],stage1_18[42],stage1_17[66],stage1_16[104]}
   );
   gpc615_5 gpc343 (
      {stage0_16[185], stage0_16[186], stage0_16[187], stage0_16[188], stage0_16[189]},
      {stage0_17[87]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[37],stage1_18[43],stage1_17[67],stage1_16[105]}
   );
   gpc615_5 gpc344 (
      {stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193], stage0_16[194]},
      {stage0_17[88]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[38],stage1_18[44],stage1_17[68],stage1_16[106]}
   );
   gpc615_5 gpc345 (
      {stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199]},
      {stage0_17[89]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[39],stage1_18[45],stage1_17[69],stage1_16[107]}
   );
   gpc615_5 gpc346 (
      {stage0_16[200], stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204]},
      {stage0_17[90]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[40],stage1_18[46],stage1_17[70],stage1_16[108]}
   );
   gpc615_5 gpc347 (
      {stage0_16[205], stage0_16[206], stage0_16[207], stage0_16[208], stage0_16[209]},
      {stage0_17[91]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[41],stage1_18[47],stage1_17[71],stage1_16[109]}
   );
   gpc615_5 gpc348 (
      {stage0_16[210], stage0_16[211], stage0_16[212], stage0_16[213], stage0_16[214]},
      {stage0_17[92]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[42],stage1_18[48],stage1_17[72],stage1_16[110]}
   );
   gpc615_5 gpc349 (
      {stage0_16[215], stage0_16[216], stage0_16[217], stage0_16[218], stage0_16[219]},
      {stage0_17[93]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[43],stage1_18[49],stage1_17[73],stage1_16[111]}
   );
   gpc615_5 gpc350 (
      {stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223], stage0_16[224]},
      {stage0_17[94]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[44],stage1_18[50],stage1_17[74],stage1_16[112]}
   );
   gpc615_5 gpc351 (
      {stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229]},
      {stage0_17[95]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[45],stage1_18[51],stage1_17[75],stage1_16[113]}
   );
   gpc615_5 gpc352 (
      {stage0_16[230], stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234]},
      {stage0_17[96]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[46],stage1_18[52],stage1_17[76],stage1_16[114]}
   );
   gpc615_5 gpc353 (
      {stage0_16[235], stage0_16[236], stage0_16[237], stage0_16[238], stage0_16[239]},
      {stage0_17[97]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[47],stage1_18[53],stage1_17[77],stage1_16[115]}
   );
   gpc615_5 gpc354 (
      {stage0_16[240], stage0_16[241], stage0_16[242], stage0_16[243], stage0_16[244]},
      {stage0_17[98]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[48],stage1_18[54],stage1_17[78],stage1_16[116]}
   );
   gpc615_5 gpc355 (
      {stage0_16[245], stage0_16[246], stage0_16[247], stage0_16[248], stage0_16[249]},
      {stage0_17[99]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[49],stage1_18[55],stage1_17[79],stage1_16[117]}
   );
   gpc615_5 gpc356 (
      {stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253], stage0_16[254]},
      {stage0_17[100]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[50],stage1_18[56],stage1_17[80],stage1_16[118]}
   );
   gpc606_5 gpc357 (
      {stage0_17[101], stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[37],stage1_19[51],stage1_18[57],stage1_17[81]}
   );
   gpc606_5 gpc358 (
      {stage0_17[107], stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[38],stage1_19[52],stage1_18[58],stage1_17[82]}
   );
   gpc606_5 gpc359 (
      {stage0_17[113], stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[39],stage1_19[53],stage1_18[59],stage1_17[83]}
   );
   gpc606_5 gpc360 (
      {stage0_17[119], stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[40],stage1_19[54],stage1_18[60],stage1_17[84]}
   );
   gpc606_5 gpc361 (
      {stage0_17[125], stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[41],stage1_19[55],stage1_18[61],stage1_17[85]}
   );
   gpc606_5 gpc362 (
      {stage0_17[131], stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[42],stage1_19[56],stage1_18[62],stage1_17[86]}
   );
   gpc606_5 gpc363 (
      {stage0_17[137], stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[43],stage1_19[57],stage1_18[63],stage1_17[87]}
   );
   gpc606_5 gpc364 (
      {stage0_17[143], stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[44],stage1_19[58],stage1_18[64],stage1_17[88]}
   );
   gpc606_5 gpc365 (
      {stage0_17[149], stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[45],stage1_19[59],stage1_18[65],stage1_17[89]}
   );
   gpc606_5 gpc366 (
      {stage0_17[155], stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[46],stage1_19[60],stage1_18[66],stage1_17[90]}
   );
   gpc606_5 gpc367 (
      {stage0_17[161], stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[47],stage1_19[61],stage1_18[67],stage1_17[91]}
   );
   gpc606_5 gpc368 (
      {stage0_17[167], stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[48],stage1_19[62],stage1_18[68],stage1_17[92]}
   );
   gpc606_5 gpc369 (
      {stage0_17[173], stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[49],stage1_19[63],stage1_18[69],stage1_17[93]}
   );
   gpc606_5 gpc370 (
      {stage0_17[179], stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[50],stage1_19[64],stage1_18[70],stage1_17[94]}
   );
   gpc606_5 gpc371 (
      {stage0_17[185], stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[51],stage1_19[65],stage1_18[71],stage1_17[95]}
   );
   gpc606_5 gpc372 (
      {stage0_17[191], stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[52],stage1_19[66],stage1_18[72],stage1_17[96]}
   );
   gpc606_5 gpc373 (
      {stage0_17[197], stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[53],stage1_19[67],stage1_18[73],stage1_17[97]}
   );
   gpc606_5 gpc374 (
      {stage0_17[203], stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[54],stage1_19[68],stage1_18[74],stage1_17[98]}
   );
   gpc606_5 gpc375 (
      {stage0_17[209], stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[55],stage1_19[69],stage1_18[75],stage1_17[99]}
   );
   gpc606_5 gpc376 (
      {stage0_17[215], stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[56],stage1_19[70],stage1_18[76],stage1_17[100]}
   );
   gpc606_5 gpc377 (
      {stage0_17[221], stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[57],stage1_19[71],stage1_18[77],stage1_17[101]}
   );
   gpc606_5 gpc378 (
      {stage0_17[227], stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[58],stage1_19[72],stage1_18[78],stage1_17[102]}
   );
   gpc606_5 gpc379 (
      {stage0_17[233], stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[59],stage1_19[73],stage1_18[79],stage1_17[103]}
   );
   gpc606_5 gpc380 (
      {stage0_17[239], stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[60],stage1_19[74],stage1_18[80],stage1_17[104]}
   );
   gpc606_5 gpc381 (
      {stage0_17[245], stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[61],stage1_19[75],stage1_18[81],stage1_17[105]}
   );
   gpc615_5 gpc382 (
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226]},
      {stage0_19[150]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[25],stage1_20[62],stage1_19[76],stage1_18[82]}
   );
   gpc615_5 gpc383 (
      {stage0_18[227], stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231]},
      {stage0_19[151]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[26],stage1_20[63],stage1_19[77],stage1_18[83]}
   );
   gpc615_5 gpc384 (
      {stage0_18[232], stage0_18[233], stage0_18[234], stage0_18[235], stage0_18[236]},
      {stage0_19[152]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[27],stage1_20[64],stage1_19[78],stage1_18[84]}
   );
   gpc615_5 gpc385 (
      {stage0_18[237], stage0_18[238], stage0_18[239], stage0_18[240], stage0_18[241]},
      {stage0_19[153]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[28],stage1_20[65],stage1_19[79],stage1_18[85]}
   );
   gpc615_5 gpc386 (
      {stage0_19[154], stage0_19[155], stage0_19[156], stage0_19[157], stage0_19[158]},
      {stage0_20[24]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[4],stage1_21[29],stage1_20[66],stage1_19[80]}
   );
   gpc615_5 gpc387 (
      {stage0_19[159], stage0_19[160], stage0_19[161], stage0_19[162], stage0_19[163]},
      {stage0_20[25]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[5],stage1_21[30],stage1_20[67],stage1_19[81]}
   );
   gpc615_5 gpc388 (
      {stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167], stage0_19[168]},
      {stage0_20[26]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[6],stage1_21[31],stage1_20[68],stage1_19[82]}
   );
   gpc615_5 gpc389 (
      {stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage0_20[27]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[7],stage1_21[32],stage1_20[69],stage1_19[83]}
   );
   gpc615_5 gpc390 (
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178]},
      {stage0_20[28]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[8],stage1_21[33],stage1_20[70],stage1_19[84]}
   );
   gpc615_5 gpc391 (
      {stage0_19[179], stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183]},
      {stage0_20[29]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[9],stage1_21[34],stage1_20[71],stage1_19[85]}
   );
   gpc615_5 gpc392 (
      {stage0_19[184], stage0_19[185], stage0_19[186], stage0_19[187], stage0_19[188]},
      {stage0_20[30]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[10],stage1_21[35],stage1_20[72],stage1_19[86]}
   );
   gpc615_5 gpc393 (
      {stage0_19[189], stage0_19[190], stage0_19[191], stage0_19[192], stage0_19[193]},
      {stage0_20[31]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[11],stage1_21[36],stage1_20[73],stage1_19[87]}
   );
   gpc615_5 gpc394 (
      {stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197], stage0_19[198]},
      {stage0_20[32]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[12],stage1_21[37],stage1_20[74],stage1_19[88]}
   );
   gpc615_5 gpc395 (
      {stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage0_20[33]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[13],stage1_21[38],stage1_20[75],stage1_19[89]}
   );
   gpc615_5 gpc396 (
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208]},
      {stage0_20[34]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[14],stage1_21[39],stage1_20[76],stage1_19[90]}
   );
   gpc615_5 gpc397 (
      {stage0_19[209], stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213]},
      {stage0_20[35]},
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage1_23[11],stage1_22[15],stage1_21[40],stage1_20[77],stage1_19[91]}
   );
   gpc615_5 gpc398 (
      {stage0_19[214], stage0_19[215], stage0_19[216], stage0_19[217], stage0_19[218]},
      {stage0_20[36]},
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage1_23[12],stage1_22[16],stage1_21[41],stage1_20[78],stage1_19[92]}
   );
   gpc615_5 gpc399 (
      {stage0_19[219], stage0_19[220], stage0_19[221], stage0_19[222], stage0_19[223]},
      {stage0_20[37]},
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage1_23[13],stage1_22[17],stage1_21[42],stage1_20[79],stage1_19[93]}
   );
   gpc1343_5 gpc400 (
      {stage0_20[38], stage0_20[39], stage0_20[40]},
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87]},
      {stage0_22[0], stage0_22[1], stage0_22[2]},
      {stage0_23[0]},
      {stage1_24[0],stage1_23[14],stage1_22[18],stage1_21[43],stage1_20[80]}
   );
   gpc1343_5 gpc401 (
      {stage0_20[41], stage0_20[42], stage0_20[43]},
      {stage0_21[88], stage0_21[89], stage0_21[90], stage0_21[91]},
      {stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage0_23[1]},
      {stage1_24[1],stage1_23[15],stage1_22[19],stage1_21[44],stage1_20[81]}
   );
   gpc1343_5 gpc402 (
      {stage0_20[44], stage0_20[45], stage0_20[46]},
      {stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage0_22[6], stage0_22[7], stage0_22[8]},
      {stage0_23[2]},
      {stage1_24[2],stage1_23[16],stage1_22[20],stage1_21[45],stage1_20[82]}
   );
   gpc1343_5 gpc403 (
      {stage0_20[47], stage0_20[48], stage0_20[49]},
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99]},
      {stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage0_23[3]},
      {stage1_24[3],stage1_23[17],stage1_22[21],stage1_21[46],stage1_20[83]}
   );
   gpc1343_5 gpc404 (
      {stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[100], stage0_21[101], stage0_21[102], stage0_21[103]},
      {stage0_22[12], stage0_22[13], stage0_22[14]},
      {stage0_23[4]},
      {stage1_24[4],stage1_23[18],stage1_22[22],stage1_21[47],stage1_20[84]}
   );
   gpc1343_5 gpc405 (
      {stage0_20[53], stage0_20[54], stage0_20[55]},
      {stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage0_23[5]},
      {stage1_24[5],stage1_23[19],stage1_22[23],stage1_21[48],stage1_20[85]}
   );
   gpc1343_5 gpc406 (
      {stage0_20[56], stage0_20[57], stage0_20[58]},
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111]},
      {stage0_22[18], stage0_22[19], stage0_22[20]},
      {stage0_23[6]},
      {stage1_24[6],stage1_23[20],stage1_22[24],stage1_21[49],stage1_20[86]}
   );
   gpc1343_5 gpc407 (
      {stage0_20[59], stage0_20[60], stage0_20[61]},
      {stage0_21[112], stage0_21[113], stage0_21[114], stage0_21[115]},
      {stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage0_23[7]},
      {stage1_24[7],stage1_23[21],stage1_22[25],stage1_21[50],stage1_20[87]}
   );
   gpc1343_5 gpc408 (
      {stage0_20[62], stage0_20[63], stage0_20[64]},
      {stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage0_22[24], stage0_22[25], stage0_22[26]},
      {stage0_23[8]},
      {stage1_24[8],stage1_23[22],stage1_22[26],stage1_21[51],stage1_20[88]}
   );
   gpc606_5 gpc409 (
      {stage0_20[65], stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69], stage0_20[70]},
      {stage0_22[27], stage0_22[28], stage0_22[29], stage0_22[30], stage0_22[31], stage0_22[32]},
      {stage1_24[9],stage1_23[23],stage1_22[27],stage1_21[52],stage1_20[89]}
   );
   gpc606_5 gpc410 (
      {stage0_20[71], stage0_20[72], stage0_20[73], stage0_20[74], stage0_20[75], stage0_20[76]},
      {stage0_22[33], stage0_22[34], stage0_22[35], stage0_22[36], stage0_22[37], stage0_22[38]},
      {stage1_24[10],stage1_23[24],stage1_22[28],stage1_21[53],stage1_20[90]}
   );
   gpc606_5 gpc411 (
      {stage0_20[77], stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81], stage0_20[82]},
      {stage0_22[39], stage0_22[40], stage0_22[41], stage0_22[42], stage0_22[43], stage0_22[44]},
      {stage1_24[11],stage1_23[25],stage1_22[29],stage1_21[54],stage1_20[91]}
   );
   gpc606_5 gpc412 (
      {stage0_20[83], stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88]},
      {stage0_22[45], stage0_22[46], stage0_22[47], stage0_22[48], stage0_22[49], stage0_22[50]},
      {stage1_24[12],stage1_23[26],stage1_22[30],stage1_21[55],stage1_20[92]}
   );
   gpc606_5 gpc413 (
      {stage0_20[89], stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94]},
      {stage0_22[51], stage0_22[52], stage0_22[53], stage0_22[54], stage0_22[55], stage0_22[56]},
      {stage1_24[13],stage1_23[27],stage1_22[31],stage1_21[56],stage1_20[93]}
   );
   gpc606_5 gpc414 (
      {stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99], stage0_20[100]},
      {stage0_22[57], stage0_22[58], stage0_22[59], stage0_22[60], stage0_22[61], stage0_22[62]},
      {stage1_24[14],stage1_23[28],stage1_22[32],stage1_21[57],stage1_20[94]}
   );
   gpc606_5 gpc415 (
      {stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105], stage0_20[106]},
      {stage0_22[63], stage0_22[64], stage0_22[65], stage0_22[66], stage0_22[67], stage0_22[68]},
      {stage1_24[15],stage1_23[29],stage1_22[33],stage1_21[58],stage1_20[95]}
   );
   gpc606_5 gpc416 (
      {stage0_20[107], stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111], stage0_20[112]},
      {stage0_22[69], stage0_22[70], stage0_22[71], stage0_22[72], stage0_22[73], stage0_22[74]},
      {stage1_24[16],stage1_23[30],stage1_22[34],stage1_21[59],stage1_20[96]}
   );
   gpc606_5 gpc417 (
      {stage0_20[113], stage0_20[114], stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118]},
      {stage0_22[75], stage0_22[76], stage0_22[77], stage0_22[78], stage0_22[79], stage0_22[80]},
      {stage1_24[17],stage1_23[31],stage1_22[35],stage1_21[60],stage1_20[97]}
   );
   gpc606_5 gpc418 (
      {stage0_20[119], stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124]},
      {stage0_22[81], stage0_22[82], stage0_22[83], stage0_22[84], stage0_22[85], stage0_22[86]},
      {stage1_24[18],stage1_23[32],stage1_22[36],stage1_21[61],stage1_20[98]}
   );
   gpc606_5 gpc419 (
      {stage0_20[125], stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130]},
      {stage0_22[87], stage0_22[88], stage0_22[89], stage0_22[90], stage0_22[91], stage0_22[92]},
      {stage1_24[19],stage1_23[33],stage1_22[37],stage1_21[62],stage1_20[99]}
   );
   gpc606_5 gpc420 (
      {stage0_20[131], stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136]},
      {stage0_22[93], stage0_22[94], stage0_22[95], stage0_22[96], stage0_22[97], stage0_22[98]},
      {stage1_24[20],stage1_23[34],stage1_22[38],stage1_21[63],stage1_20[100]}
   );
   gpc606_5 gpc421 (
      {stage0_20[137], stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141], stage0_20[142]},
      {stage0_22[99], stage0_22[100], stage0_22[101], stage0_22[102], stage0_22[103], stage0_22[104]},
      {stage1_24[21],stage1_23[35],stage1_22[39],stage1_21[64],stage1_20[101]}
   );
   gpc606_5 gpc422 (
      {stage0_20[143], stage0_20[144], stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148]},
      {stage0_22[105], stage0_22[106], stage0_22[107], stage0_22[108], stage0_22[109], stage0_22[110]},
      {stage1_24[22],stage1_23[36],stage1_22[40],stage1_21[65],stage1_20[102]}
   );
   gpc606_5 gpc423 (
      {stage0_20[149], stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154]},
      {stage0_22[111], stage0_22[112], stage0_22[113], stage0_22[114], stage0_22[115], stage0_22[116]},
      {stage1_24[23],stage1_23[37],stage1_22[41],stage1_21[66],stage1_20[103]}
   );
   gpc606_5 gpc424 (
      {stage0_20[155], stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160]},
      {stage0_22[117], stage0_22[118], stage0_22[119], stage0_22[120], stage0_22[121], stage0_22[122]},
      {stage1_24[24],stage1_23[38],stage1_22[42],stage1_21[67],stage1_20[104]}
   );
   gpc606_5 gpc425 (
      {stage0_20[161], stage0_20[162], stage0_20[163], stage0_20[164], stage0_20[165], stage0_20[166]},
      {stage0_22[123], stage0_22[124], stage0_22[125], stage0_22[126], stage0_22[127], stage0_22[128]},
      {stage1_24[25],stage1_23[39],stage1_22[43],stage1_21[68],stage1_20[105]}
   );
   gpc606_5 gpc426 (
      {stage0_20[167], stage0_20[168], stage0_20[169], stage0_20[170], stage0_20[171], stage0_20[172]},
      {stage0_22[129], stage0_22[130], stage0_22[131], stage0_22[132], stage0_22[133], stage0_22[134]},
      {stage1_24[26],stage1_23[40],stage1_22[44],stage1_21[69],stage1_20[106]}
   );
   gpc606_5 gpc427 (
      {stage0_20[173], stage0_20[174], stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178]},
      {stage0_22[135], stage0_22[136], stage0_22[137], stage0_22[138], stage0_22[139], stage0_22[140]},
      {stage1_24[27],stage1_23[41],stage1_22[45],stage1_21[70],stage1_20[107]}
   );
   gpc606_5 gpc428 (
      {stage0_20[179], stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184]},
      {stage0_22[141], stage0_22[142], stage0_22[143], stage0_22[144], stage0_22[145], stage0_22[146]},
      {stage1_24[28],stage1_23[42],stage1_22[46],stage1_21[71],stage1_20[108]}
   );
   gpc606_5 gpc429 (
      {stage0_20[185], stage0_20[186], stage0_20[187], stage0_20[188], stage0_20[189], stage0_20[190]},
      {stage0_22[147], stage0_22[148], stage0_22[149], stage0_22[150], stage0_22[151], stage0_22[152]},
      {stage1_24[29],stage1_23[43],stage1_22[47],stage1_21[72],stage1_20[109]}
   );
   gpc606_5 gpc430 (
      {stage0_20[191], stage0_20[192], stage0_20[193], stage0_20[194], stage0_20[195], stage0_20[196]},
      {stage0_22[153], stage0_22[154], stage0_22[155], stage0_22[156], stage0_22[157], stage0_22[158]},
      {stage1_24[30],stage1_23[44],stage1_22[48],stage1_21[73],stage1_20[110]}
   );
   gpc606_5 gpc431 (
      {stage0_20[197], stage0_20[198], stage0_20[199], stage0_20[200], stage0_20[201], stage0_20[202]},
      {stage0_22[159], stage0_22[160], stage0_22[161], stage0_22[162], stage0_22[163], stage0_22[164]},
      {stage1_24[31],stage1_23[45],stage1_22[49],stage1_21[74],stage1_20[111]}
   );
   gpc606_5 gpc432 (
      {stage0_20[203], stage0_20[204], stage0_20[205], stage0_20[206], stage0_20[207], stage0_20[208]},
      {stage0_22[165], stage0_22[166], stage0_22[167], stage0_22[168], stage0_22[169], stage0_22[170]},
      {stage1_24[32],stage1_23[46],stage1_22[50],stage1_21[75],stage1_20[112]}
   );
   gpc606_5 gpc433 (
      {stage0_20[209], stage0_20[210], stage0_20[211], stage0_20[212], stage0_20[213], stage0_20[214]},
      {stage0_22[171], stage0_22[172], stage0_22[173], stage0_22[174], stage0_22[175], stage0_22[176]},
      {stage1_24[33],stage1_23[47],stage1_22[51],stage1_21[76],stage1_20[113]}
   );
   gpc606_5 gpc434 (
      {stage0_20[215], stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219], stage0_20[220]},
      {stage0_22[177], stage0_22[178], stage0_22[179], stage0_22[180], stage0_22[181], stage0_22[182]},
      {stage1_24[34],stage1_23[48],stage1_22[52],stage1_21[77],stage1_20[114]}
   );
   gpc606_5 gpc435 (
      {stage0_20[221], stage0_20[222], stage0_20[223], stage0_20[224], stage0_20[225], stage0_20[226]},
      {stage0_22[183], stage0_22[184], stage0_22[185], stage0_22[186], stage0_22[187], stage0_22[188]},
      {stage1_24[35],stage1_23[49],stage1_22[53],stage1_21[78],stage1_20[115]}
   );
   gpc606_5 gpc436 (
      {stage0_20[227], stage0_20[228], stage0_20[229], stage0_20[230], stage0_20[231], stage0_20[232]},
      {stage0_22[189], stage0_22[190], stage0_22[191], stage0_22[192], stage0_22[193], stage0_22[194]},
      {stage1_24[36],stage1_23[50],stage1_22[54],stage1_21[79],stage1_20[116]}
   );
   gpc606_5 gpc437 (
      {stage0_20[233], stage0_20[234], stage0_20[235], stage0_20[236], stage0_20[237], stage0_20[238]},
      {stage0_22[195], stage0_22[196], stage0_22[197], stage0_22[198], stage0_22[199], stage0_22[200]},
      {stage1_24[37],stage1_23[51],stage1_22[55],stage1_21[80],stage1_20[117]}
   );
   gpc606_5 gpc438 (
      {stage0_20[239], stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243], stage0_20[244]},
      {stage0_22[201], stage0_22[202], stage0_22[203], stage0_22[204], stage0_22[205], stage0_22[206]},
      {stage1_24[38],stage1_23[52],stage1_22[56],stage1_21[81],stage1_20[118]}
   );
   gpc606_5 gpc439 (
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage0_23[9], stage0_23[10], stage0_23[11], stage0_23[12], stage0_23[13], stage0_23[14]},
      {stage1_25[0],stage1_24[39],stage1_23[53],stage1_22[57],stage1_21[82]}
   );
   gpc606_5 gpc440 (
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage0_23[15], stage0_23[16], stage0_23[17], stage0_23[18], stage0_23[19], stage0_23[20]},
      {stage1_25[1],stage1_24[40],stage1_23[54],stage1_22[58],stage1_21[83]}
   );
   gpc606_5 gpc441 (
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage0_23[21], stage0_23[22], stage0_23[23], stage0_23[24], stage0_23[25], stage0_23[26]},
      {stage1_25[2],stage1_24[41],stage1_23[55],stage1_22[59],stage1_21[84]}
   );
   gpc606_5 gpc442 (
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage0_23[27], stage0_23[28], stage0_23[29], stage0_23[30], stage0_23[31], stage0_23[32]},
      {stage1_25[3],stage1_24[42],stage1_23[56],stage1_22[60],stage1_21[85]}
   );
   gpc606_5 gpc443 (
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage0_23[33], stage0_23[34], stage0_23[35], stage0_23[36], stage0_23[37], stage0_23[38]},
      {stage1_25[4],stage1_24[43],stage1_23[57],stage1_22[61],stage1_21[86]}
   );
   gpc606_5 gpc444 (
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage0_23[39], stage0_23[40], stage0_23[41], stage0_23[42], stage0_23[43], stage0_23[44]},
      {stage1_25[5],stage1_24[44],stage1_23[58],stage1_22[62],stage1_21[87]}
   );
   gpc606_5 gpc445 (
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage0_23[45], stage0_23[46], stage0_23[47], stage0_23[48], stage0_23[49], stage0_23[50]},
      {stage1_25[6],stage1_24[45],stage1_23[59],stage1_22[63],stage1_21[88]}
   );
   gpc606_5 gpc446 (
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage0_23[51], stage0_23[52], stage0_23[53], stage0_23[54], stage0_23[55], stage0_23[56]},
      {stage1_25[7],stage1_24[46],stage1_23[60],stage1_22[64],stage1_21[89]}
   );
   gpc606_5 gpc447 (
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage0_23[57], stage0_23[58], stage0_23[59], stage0_23[60], stage0_23[61], stage0_23[62]},
      {stage1_25[8],stage1_24[47],stage1_23[61],stage1_22[65],stage1_21[90]}
   );
   gpc606_5 gpc448 (
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage0_23[63], stage0_23[64], stage0_23[65], stage0_23[66], stage0_23[67], stage0_23[68]},
      {stage1_25[9],stage1_24[48],stage1_23[62],stage1_22[66],stage1_21[91]}
   );
   gpc606_5 gpc449 (
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage0_23[69], stage0_23[70], stage0_23[71], stage0_23[72], stage0_23[73], stage0_23[74]},
      {stage1_25[10],stage1_24[49],stage1_23[63],stage1_22[67],stage1_21[92]}
   );
   gpc606_5 gpc450 (
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage0_23[75], stage0_23[76], stage0_23[77], stage0_23[78], stage0_23[79], stage0_23[80]},
      {stage1_25[11],stage1_24[50],stage1_23[64],stage1_22[68],stage1_21[93]}
   );
   gpc606_5 gpc451 (
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage0_23[81], stage0_23[82], stage0_23[83], stage0_23[84], stage0_23[85], stage0_23[86]},
      {stage1_25[12],stage1_24[51],stage1_23[65],stage1_22[69],stage1_21[94]}
   );
   gpc606_5 gpc452 (
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage0_23[87], stage0_23[88], stage0_23[89], stage0_23[90], stage0_23[91], stage0_23[92]},
      {stage1_25[13],stage1_24[52],stage1_23[66],stage1_22[70],stage1_21[95]}
   );
   gpc606_5 gpc453 (
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage0_23[93], stage0_23[94], stage0_23[95], stage0_23[96], stage0_23[97], stage0_23[98]},
      {stage1_25[14],stage1_24[53],stage1_23[67],stage1_22[71],stage1_21[96]}
   );
   gpc606_5 gpc454 (
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage0_23[99], stage0_23[100], stage0_23[101], stage0_23[102], stage0_23[103], stage0_23[104]},
      {stage1_25[15],stage1_24[54],stage1_23[68],stage1_22[72],stage1_21[97]}
   );
   gpc606_5 gpc455 (
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage0_23[105], stage0_23[106], stage0_23[107], stage0_23[108], stage0_23[109], stage0_23[110]},
      {stage1_25[16],stage1_24[55],stage1_23[69],stage1_22[73],stage1_21[98]}
   );
   gpc606_5 gpc456 (
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage0_23[111], stage0_23[112], stage0_23[113], stage0_23[114], stage0_23[115], stage0_23[116]},
      {stage1_25[17],stage1_24[56],stage1_23[70],stage1_22[74],stage1_21[99]}
   );
   gpc606_5 gpc457 (
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage0_23[117], stage0_23[118], stage0_23[119], stage0_23[120], stage0_23[121], stage0_23[122]},
      {stage1_25[18],stage1_24[57],stage1_23[71],stage1_22[75],stage1_21[100]}
   );
   gpc606_5 gpc458 (
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage0_23[123], stage0_23[124], stage0_23[125], stage0_23[126], stage0_23[127], stage0_23[128]},
      {stage1_25[19],stage1_24[58],stage1_23[72],stage1_22[76],stage1_21[101]}
   );
   gpc606_5 gpc459 (
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage0_23[129], stage0_23[130], stage0_23[131], stage0_23[132], stage0_23[133], stage0_23[134]},
      {stage1_25[20],stage1_24[59],stage1_23[73],stage1_22[77],stage1_21[102]}
   );
   gpc606_5 gpc460 (
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249], stage0_21[250], stage0_21[251]},
      {stage0_23[135], stage0_23[136], stage0_23[137], stage0_23[138], stage0_23[139], stage0_23[140]},
      {stage1_25[21],stage1_24[60],stage1_23[74],stage1_22[78],stage1_21[103]}
   );
   gpc615_5 gpc461 (
      {stage0_22[207], stage0_22[208], stage0_22[209], stage0_22[210], stage0_22[211]},
      {stage0_23[141]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[22],stage1_24[61],stage1_23[75],stage1_22[79]}
   );
   gpc615_5 gpc462 (
      {stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215], stage0_22[216]},
      {stage0_23[142]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[23],stage1_24[62],stage1_23[76],stage1_22[80]}
   );
   gpc615_5 gpc463 (
      {stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage0_23[143]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[24],stage1_24[63],stage1_23[77],stage1_22[81]}
   );
   gpc615_5 gpc464 (
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226]},
      {stage0_23[144]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[25],stage1_24[64],stage1_23[78],stage1_22[82]}
   );
   gpc615_5 gpc465 (
      {stage0_22[227], stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231]},
      {stage0_23[145]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[26],stage1_24[65],stage1_23[79],stage1_22[83]}
   );
   gpc615_5 gpc466 (
      {stage0_22[232], stage0_22[233], stage0_22[234], stage0_22[235], stage0_22[236]},
      {stage0_23[146]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[27],stage1_24[66],stage1_23[80],stage1_22[84]}
   );
   gpc615_5 gpc467 (
      {stage0_22[237], stage0_22[238], stage0_22[239], stage0_22[240], stage0_22[241]},
      {stage0_23[147]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[28],stage1_24[67],stage1_23[81],stage1_22[85]}
   );
   gpc615_5 gpc468 (
      {stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245], stage0_22[246]},
      {stage0_23[148]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[29],stage1_24[68],stage1_23[82],stage1_22[86]}
   );
   gpc615_5 gpc469 (
      {stage0_22[247], stage0_22[248], stage0_22[249], stage0_22[250], stage0_22[251]},
      {stage0_23[149]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[30],stage1_24[69],stage1_23[83],stage1_22[87]}
   );
   gpc606_5 gpc470 (
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[9],stage1_25[31],stage1_24[70],stage1_23[84]}
   );
   gpc615_5 gpc471 (
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160]},
      {stage0_24[54]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[10],stage1_25[32],stage1_24[71],stage1_23[85]}
   );
   gpc615_5 gpc472 (
      {stage0_23[161], stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165]},
      {stage0_24[55]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[11],stage1_25[33],stage1_24[72],stage1_23[86]}
   );
   gpc615_5 gpc473 (
      {stage0_23[166], stage0_23[167], stage0_23[168], stage0_23[169], stage0_23[170]},
      {stage0_24[56]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[12],stage1_25[34],stage1_24[73],stage1_23[87]}
   );
   gpc615_5 gpc474 (
      {stage0_23[171], stage0_23[172], stage0_23[173], stage0_23[174], stage0_23[175]},
      {stage0_24[57]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[13],stage1_25[35],stage1_24[74],stage1_23[88]}
   );
   gpc615_5 gpc475 (
      {stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179], stage0_23[180]},
      {stage0_24[58]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[14],stage1_25[36],stage1_24[75],stage1_23[89]}
   );
   gpc615_5 gpc476 (
      {stage0_23[181], stage0_23[182], stage0_23[183], stage0_23[184], stage0_23[185]},
      {stage0_24[59]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[15],stage1_25[37],stage1_24[76],stage1_23[90]}
   );
   gpc615_5 gpc477 (
      {stage0_23[186], stage0_23[187], stage0_23[188], stage0_23[189], stage0_23[190]},
      {stage0_24[60]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[16],stage1_25[38],stage1_24[77],stage1_23[91]}
   );
   gpc615_5 gpc478 (
      {stage0_23[191], stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195]},
      {stage0_24[61]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[17],stage1_25[39],stage1_24[78],stage1_23[92]}
   );
   gpc615_5 gpc479 (
      {stage0_23[196], stage0_23[197], stage0_23[198], stage0_23[199], stage0_23[200]},
      {stage0_24[62]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[18],stage1_25[40],stage1_24[79],stage1_23[93]}
   );
   gpc615_5 gpc480 (
      {stage0_23[201], stage0_23[202], stage0_23[203], stage0_23[204], stage0_23[205]},
      {stage0_24[63]},
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage1_27[10],stage1_26[19],stage1_25[41],stage1_24[80],stage1_23[94]}
   );
   gpc615_5 gpc481 (
      {stage0_23[206], stage0_23[207], stage0_23[208], stage0_23[209], stage0_23[210]},
      {stage0_24[64]},
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage1_27[11],stage1_26[20],stage1_25[42],stage1_24[81],stage1_23[95]}
   );
   gpc615_5 gpc482 (
      {stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214], stage0_23[215]},
      {stage0_24[65]},
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage1_27[12],stage1_26[21],stage1_25[43],stage1_24[82],stage1_23[96]}
   );
   gpc615_5 gpc483 (
      {stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220]},
      {stage0_24[66]},
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage1_27[13],stage1_26[22],stage1_25[44],stage1_24[83],stage1_23[97]}
   );
   gpc615_5 gpc484 (
      {stage0_23[221], stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225]},
      {stage0_24[67]},
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage1_27[14],stage1_26[23],stage1_25[45],stage1_24[84],stage1_23[98]}
   );
   gpc606_5 gpc485 (
      {stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71], stage0_24[72], stage0_24[73]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[15],stage1_26[24],stage1_25[46],stage1_24[85]}
   );
   gpc606_5 gpc486 (
      {stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77], stage0_24[78], stage0_24[79]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[16],stage1_26[25],stage1_25[47],stage1_24[86]}
   );
   gpc606_5 gpc487 (
      {stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83], stage0_24[84], stage0_24[85]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[17],stage1_26[26],stage1_25[48],stage1_24[87]}
   );
   gpc606_5 gpc488 (
      {stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89], stage0_24[90], stage0_24[91]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[18],stage1_26[27],stage1_25[49],stage1_24[88]}
   );
   gpc606_5 gpc489 (
      {stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95], stage0_24[96], stage0_24[97]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[19],stage1_26[28],stage1_25[50],stage1_24[89]}
   );
   gpc606_5 gpc490 (
      {stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101], stage0_24[102], stage0_24[103]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[20],stage1_26[29],stage1_25[51],stage1_24[90]}
   );
   gpc606_5 gpc491 (
      {stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107], stage0_24[108], stage0_24[109]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[21],stage1_26[30],stage1_25[52],stage1_24[91]}
   );
   gpc606_5 gpc492 (
      {stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113], stage0_24[114], stage0_24[115]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[22],stage1_26[31],stage1_25[53],stage1_24[92]}
   );
   gpc606_5 gpc493 (
      {stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119], stage0_24[120], stage0_24[121]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[23],stage1_26[32],stage1_25[54],stage1_24[93]}
   );
   gpc606_5 gpc494 (
      {stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125], stage0_24[126], stage0_24[127]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[24],stage1_26[33],stage1_25[55],stage1_24[94]}
   );
   gpc606_5 gpc495 (
      {stage0_24[128], stage0_24[129], stage0_24[130], stage0_24[131], stage0_24[132], stage0_24[133]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[25],stage1_26[34],stage1_25[56],stage1_24[95]}
   );
   gpc606_5 gpc496 (
      {stage0_24[134], stage0_24[135], stage0_24[136], stage0_24[137], stage0_24[138], stage0_24[139]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[26],stage1_26[35],stage1_25[57],stage1_24[96]}
   );
   gpc606_5 gpc497 (
      {stage0_24[140], stage0_24[141], stage0_24[142], stage0_24[143], stage0_24[144], stage0_24[145]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[27],stage1_26[36],stage1_25[58],stage1_24[97]}
   );
   gpc615_5 gpc498 (
      {stage0_24[146], stage0_24[147], stage0_24[148], stage0_24[149], stage0_24[150]},
      {stage0_25[90]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[28],stage1_26[37],stage1_25[59],stage1_24[98]}
   );
   gpc615_5 gpc499 (
      {stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154], stage0_24[155]},
      {stage0_25[91]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[29],stage1_26[38],stage1_25[60],stage1_24[99]}
   );
   gpc615_5 gpc500 (
      {stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160]},
      {stage0_25[92]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[30],stage1_26[39],stage1_25[61],stage1_24[100]}
   );
   gpc615_5 gpc501 (
      {stage0_24[161], stage0_24[162], stage0_24[163], stage0_24[164], stage0_24[165]},
      {stage0_25[93]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[31],stage1_26[40],stage1_25[62],stage1_24[101]}
   );
   gpc615_5 gpc502 (
      {stage0_24[166], stage0_24[167], stage0_24[168], stage0_24[169], stage0_24[170]},
      {stage0_25[94]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[32],stage1_26[41],stage1_25[63],stage1_24[102]}
   );
   gpc615_5 gpc503 (
      {stage0_24[171], stage0_24[172], stage0_24[173], stage0_24[174], stage0_24[175]},
      {stage0_25[95]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[33],stage1_26[42],stage1_25[64],stage1_24[103]}
   );
   gpc615_5 gpc504 (
      {stage0_24[176], stage0_24[177], stage0_24[178], stage0_24[179], stage0_24[180]},
      {stage0_25[96]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[34],stage1_26[43],stage1_25[65],stage1_24[104]}
   );
   gpc615_5 gpc505 (
      {stage0_24[181], stage0_24[182], stage0_24[183], stage0_24[184], stage0_24[185]},
      {stage0_25[97]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[35],stage1_26[44],stage1_25[66],stage1_24[105]}
   );
   gpc615_5 gpc506 (
      {stage0_24[186], stage0_24[187], stage0_24[188], stage0_24[189], stage0_24[190]},
      {stage0_25[98]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[36],stage1_26[45],stage1_25[67],stage1_24[106]}
   );
   gpc615_5 gpc507 (
      {stage0_24[191], stage0_24[192], stage0_24[193], stage0_24[194], stage0_24[195]},
      {stage0_25[99]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[37],stage1_26[46],stage1_25[68],stage1_24[107]}
   );
   gpc615_5 gpc508 (
      {stage0_24[196], stage0_24[197], stage0_24[198], stage0_24[199], stage0_24[200]},
      {stage0_25[100]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[38],stage1_26[47],stage1_25[69],stage1_24[108]}
   );
   gpc615_5 gpc509 (
      {stage0_24[201], stage0_24[202], stage0_24[203], stage0_24[204], stage0_24[205]},
      {stage0_25[101]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[39],stage1_26[48],stage1_25[70],stage1_24[109]}
   );
   gpc615_5 gpc510 (
      {stage0_24[206], stage0_24[207], stage0_24[208], stage0_24[209], stage0_24[210]},
      {stage0_25[102]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[40],stage1_26[49],stage1_25[71],stage1_24[110]}
   );
   gpc615_5 gpc511 (
      {stage0_24[211], stage0_24[212], stage0_24[213], stage0_24[214], stage0_24[215]},
      {stage0_25[103]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[41],stage1_26[50],stage1_25[72],stage1_24[111]}
   );
   gpc615_5 gpc512 (
      {stage0_24[216], stage0_24[217], stage0_24[218], stage0_24[219], stage0_24[220]},
      {stage0_25[104]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[42],stage1_26[51],stage1_25[73],stage1_24[112]}
   );
   gpc615_5 gpc513 (
      {stage0_24[221], stage0_24[222], stage0_24[223], stage0_24[224], stage0_24[225]},
      {stage0_25[105]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[43],stage1_26[52],stage1_25[74],stage1_24[113]}
   );
   gpc615_5 gpc514 (
      {stage0_24[226], stage0_24[227], stage0_24[228], stage0_24[229], stage0_24[230]},
      {stage0_25[106]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[44],stage1_26[53],stage1_25[75],stage1_24[114]}
   );
   gpc606_5 gpc515 (
      {stage0_25[107], stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[30],stage1_27[45],stage1_26[54],stage1_25[76]}
   );
   gpc606_5 gpc516 (
      {stage0_25[113], stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117], stage0_25[118]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[31],stage1_27[46],stage1_26[55],stage1_25[77]}
   );
   gpc606_5 gpc517 (
      {stage0_25[119], stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123], stage0_25[124]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[32],stage1_27[47],stage1_26[56],stage1_25[78]}
   );
   gpc606_5 gpc518 (
      {stage0_25[125], stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129], stage0_25[130]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[33],stage1_27[48],stage1_26[57],stage1_25[79]}
   );
   gpc606_5 gpc519 (
      {stage0_25[131], stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[34],stage1_27[49],stage1_26[58],stage1_25[80]}
   );
   gpc606_5 gpc520 (
      {stage0_25[137], stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[35],stage1_27[50],stage1_26[59],stage1_25[81]}
   );
   gpc606_5 gpc521 (
      {stage0_25[143], stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147], stage0_25[148]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[36],stage1_27[51],stage1_26[60],stage1_25[82]}
   );
   gpc606_5 gpc522 (
      {stage0_25[149], stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153], stage0_25[154]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[37],stage1_27[52],stage1_26[61],stage1_25[83]}
   );
   gpc606_5 gpc523 (
      {stage0_25[155], stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159], stage0_25[160]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[38],stage1_27[53],stage1_26[62],stage1_25[84]}
   );
   gpc606_5 gpc524 (
      {stage0_25[161], stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165], stage0_25[166]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[39],stage1_27[54],stage1_26[63],stage1_25[85]}
   );
   gpc606_5 gpc525 (
      {stage0_25[167], stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171], stage0_25[172]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[40],stage1_27[55],stage1_26[64],stage1_25[86]}
   );
   gpc606_5 gpc526 (
      {stage0_25[173], stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177], stage0_25[178]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[41],stage1_27[56],stage1_26[65],stage1_25[87]}
   );
   gpc606_5 gpc527 (
      {stage0_25[179], stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183], stage0_25[184]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[42],stage1_27[57],stage1_26[66],stage1_25[88]}
   );
   gpc606_5 gpc528 (
      {stage0_25[185], stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189], stage0_25[190]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[43],stage1_27[58],stage1_26[67],stage1_25[89]}
   );
   gpc606_5 gpc529 (
      {stage0_25[191], stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195], stage0_25[196]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[44],stage1_27[59],stage1_26[68],stage1_25[90]}
   );
   gpc606_5 gpc530 (
      {stage0_25[197], stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201], stage0_25[202]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[45],stage1_27[60],stage1_26[69],stage1_25[91]}
   );
   gpc606_5 gpc531 (
      {stage0_25[203], stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207], stage0_25[208]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[46],stage1_27[61],stage1_26[70],stage1_25[92]}
   );
   gpc606_5 gpc532 (
      {stage0_25[209], stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213], stage0_25[214]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[47],stage1_27[62],stage1_26[71],stage1_25[93]}
   );
   gpc606_5 gpc533 (
      {stage0_25[215], stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219], stage0_25[220]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[48],stage1_27[63],stage1_26[72],stage1_25[94]}
   );
   gpc606_5 gpc534 (
      {stage0_25[221], stage0_25[222], stage0_25[223], stage0_25[224], stage0_25[225], stage0_25[226]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[49],stage1_27[64],stage1_26[73],stage1_25[95]}
   );
   gpc606_5 gpc535 (
      {stage0_25[227], stage0_25[228], stage0_25[229], stage0_25[230], stage0_25[231], stage0_25[232]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[50],stage1_27[65],stage1_26[74],stage1_25[96]}
   );
   gpc606_5 gpc536 (
      {stage0_25[233], stage0_25[234], stage0_25[235], stage0_25[236], stage0_25[237], stage0_25[238]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[51],stage1_27[66],stage1_26[75],stage1_25[97]}
   );
   gpc606_5 gpc537 (
      {stage0_25[239], stage0_25[240], stage0_25[241], stage0_25[242], stage0_25[243], stage0_25[244]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[52],stage1_27[67],stage1_26[76],stage1_25[98]}
   );
   gpc615_5 gpc538 (
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184]},
      {stage0_27[138]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[23],stage1_28[53],stage1_27[68],stage1_26[77]}
   );
   gpc615_5 gpc539 (
      {stage0_26[185], stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189]},
      {stage0_27[139]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[24],stage1_28[54],stage1_27[69],stage1_26[78]}
   );
   gpc615_5 gpc540 (
      {stage0_26[190], stage0_26[191], stage0_26[192], stage0_26[193], stage0_26[194]},
      {stage0_27[140]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[25],stage1_28[55],stage1_27[70],stage1_26[79]}
   );
   gpc606_5 gpc541 (
      {stage0_27[141], stage0_27[142], stage0_27[143], stage0_27[144], stage0_27[145], stage0_27[146]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[3],stage1_29[26],stage1_28[56],stage1_27[71]}
   );
   gpc606_5 gpc542 (
      {stage0_27[147], stage0_27[148], stage0_27[149], stage0_27[150], stage0_27[151], stage0_27[152]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[4],stage1_29[27],stage1_28[57],stage1_27[72]}
   );
   gpc606_5 gpc543 (
      {stage0_27[153], stage0_27[154], stage0_27[155], stage0_27[156], stage0_27[157], stage0_27[158]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[5],stage1_29[28],stage1_28[58],stage1_27[73]}
   );
   gpc615_5 gpc544 (
      {stage0_27[159], stage0_27[160], stage0_27[161], stage0_27[162], stage0_27[163]},
      {stage0_28[18]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[6],stage1_29[29],stage1_28[59],stage1_27[74]}
   );
   gpc615_5 gpc545 (
      {stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167], stage0_27[168]},
      {stage0_28[19]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[7],stage1_29[30],stage1_28[60],stage1_27[75]}
   );
   gpc615_5 gpc546 (
      {stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage0_28[20]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[8],stage1_29[31],stage1_28[61],stage1_27[76]}
   );
   gpc615_5 gpc547 (
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178]},
      {stage0_28[21]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[9],stage1_29[32],stage1_28[62],stage1_27[77]}
   );
   gpc615_5 gpc548 (
      {stage0_27[179], stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183]},
      {stage0_28[22]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[10],stage1_29[33],stage1_28[63],stage1_27[78]}
   );
   gpc615_5 gpc549 (
      {stage0_27[184], stage0_27[185], stage0_27[186], stage0_27[187], stage0_27[188]},
      {stage0_28[23]},
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage1_31[8],stage1_30[11],stage1_29[34],stage1_28[64],stage1_27[79]}
   );
   gpc615_5 gpc550 (
      {stage0_27[189], stage0_27[190], stage0_27[191], stage0_27[192], stage0_27[193]},
      {stage0_28[24]},
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage1_31[9],stage1_30[12],stage1_29[35],stage1_28[65],stage1_27[80]}
   );
   gpc615_5 gpc551 (
      {stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197], stage0_27[198]},
      {stage0_28[25]},
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage1_31[10],stage1_30[13],stage1_29[36],stage1_28[66],stage1_27[81]}
   );
   gpc615_5 gpc552 (
      {stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage0_28[26]},
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage1_31[11],stage1_30[14],stage1_29[37],stage1_28[67],stage1_27[82]}
   );
   gpc615_5 gpc553 (
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208]},
      {stage0_28[27]},
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage1_31[12],stage1_30[15],stage1_29[38],stage1_28[68],stage1_27[83]}
   );
   gpc615_5 gpc554 (
      {stage0_27[209], stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213]},
      {stage0_28[28]},
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage1_31[13],stage1_30[16],stage1_29[39],stage1_28[69],stage1_27[84]}
   );
   gpc615_5 gpc555 (
      {stage0_27[214], stage0_27[215], stage0_27[216], stage0_27[217], stage0_27[218]},
      {stage0_28[29]},
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage1_31[14],stage1_30[17],stage1_29[40],stage1_28[70],stage1_27[85]}
   );
   gpc615_5 gpc556 (
      {stage0_27[219], stage0_27[220], stage0_27[221], stage0_27[222], stage0_27[223]},
      {stage0_28[30]},
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage1_31[15],stage1_30[18],stage1_29[41],stage1_28[71],stage1_27[86]}
   );
   gpc2116_5 gpc557 (
      {stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35], stage0_28[36]},
      {stage0_29[96]},
      {stage0_30[0]},
      {stage0_31[0], stage0_31[1]},
      {stage1_32[0],stage1_31[16],stage1_30[19],stage1_29[42],stage1_28[72]}
   );
   gpc606_5 gpc558 (
      {stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41], stage0_28[42]},
      {stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5], stage0_30[6]},
      {stage1_32[1],stage1_31[17],stage1_30[20],stage1_29[43],stage1_28[73]}
   );
   gpc606_5 gpc559 (
      {stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47], stage0_28[48]},
      {stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11], stage0_30[12]},
      {stage1_32[2],stage1_31[18],stage1_30[21],stage1_29[44],stage1_28[74]}
   );
   gpc606_5 gpc560 (
      {stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53], stage0_28[54]},
      {stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17], stage0_30[18]},
      {stage1_32[3],stage1_31[19],stage1_30[22],stage1_29[45],stage1_28[75]}
   );
   gpc606_5 gpc561 (
      {stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59], stage0_28[60]},
      {stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23], stage0_30[24]},
      {stage1_32[4],stage1_31[20],stage1_30[23],stage1_29[46],stage1_28[76]}
   );
   gpc606_5 gpc562 (
      {stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65], stage0_28[66]},
      {stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29], stage0_30[30]},
      {stage1_32[5],stage1_31[21],stage1_30[24],stage1_29[47],stage1_28[77]}
   );
   gpc606_5 gpc563 (
      {stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71], stage0_28[72]},
      {stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35], stage0_30[36]},
      {stage1_32[6],stage1_31[22],stage1_30[25],stage1_29[48],stage1_28[78]}
   );
   gpc606_5 gpc564 (
      {stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77], stage0_28[78]},
      {stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41], stage0_30[42]},
      {stage1_32[7],stage1_31[23],stage1_30[26],stage1_29[49],stage1_28[79]}
   );
   gpc606_5 gpc565 (
      {stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83], stage0_28[84]},
      {stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47], stage0_30[48]},
      {stage1_32[8],stage1_31[24],stage1_30[27],stage1_29[50],stage1_28[80]}
   );
   gpc606_5 gpc566 (
      {stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89], stage0_28[90]},
      {stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53], stage0_30[54]},
      {stage1_32[9],stage1_31[25],stage1_30[28],stage1_29[51],stage1_28[81]}
   );
   gpc606_5 gpc567 (
      {stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95], stage0_28[96]},
      {stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59], stage0_30[60]},
      {stage1_32[10],stage1_31[26],stage1_30[29],stage1_29[52],stage1_28[82]}
   );
   gpc606_5 gpc568 (
      {stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101], stage0_28[102]},
      {stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65], stage0_30[66]},
      {stage1_32[11],stage1_31[27],stage1_30[30],stage1_29[53],stage1_28[83]}
   );
   gpc606_5 gpc569 (
      {stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107], stage0_28[108]},
      {stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71], stage0_30[72]},
      {stage1_32[12],stage1_31[28],stage1_30[31],stage1_29[54],stage1_28[84]}
   );
   gpc606_5 gpc570 (
      {stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114]},
      {stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77], stage0_30[78]},
      {stage1_32[13],stage1_31[29],stage1_30[32],stage1_29[55],stage1_28[85]}
   );
   gpc606_5 gpc571 (
      {stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120]},
      {stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83], stage0_30[84]},
      {stage1_32[14],stage1_31[30],stage1_30[33],stage1_29[56],stage1_28[86]}
   );
   gpc606_5 gpc572 (
      {stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126]},
      {stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89], stage0_30[90]},
      {stage1_32[15],stage1_31[31],stage1_30[34],stage1_29[57],stage1_28[87]}
   );
   gpc606_5 gpc573 (
      {stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132]},
      {stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95], stage0_30[96]},
      {stage1_32[16],stage1_31[32],stage1_30[35],stage1_29[58],stage1_28[88]}
   );
   gpc606_5 gpc574 (
      {stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138]},
      {stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101], stage0_30[102]},
      {stage1_32[17],stage1_31[33],stage1_30[36],stage1_29[59],stage1_28[89]}
   );
   gpc606_5 gpc575 (
      {stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143], stage0_28[144]},
      {stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107], stage0_30[108]},
      {stage1_32[18],stage1_31[34],stage1_30[37],stage1_29[60],stage1_28[90]}
   );
   gpc606_5 gpc576 (
      {stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149], stage0_28[150]},
      {stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113], stage0_30[114]},
      {stage1_32[19],stage1_31[35],stage1_30[38],stage1_29[61],stage1_28[91]}
   );
   gpc606_5 gpc577 (
      {stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155], stage0_28[156]},
      {stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119], stage0_30[120]},
      {stage1_32[20],stage1_31[36],stage1_30[39],stage1_29[62],stage1_28[92]}
   );
   gpc606_5 gpc578 (
      {stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161], stage0_28[162]},
      {stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125], stage0_30[126]},
      {stage1_32[21],stage1_31[37],stage1_30[40],stage1_29[63],stage1_28[93]}
   );
   gpc606_5 gpc579 (
      {stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167], stage0_28[168]},
      {stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131], stage0_30[132]},
      {stage1_32[22],stage1_31[38],stage1_30[41],stage1_29[64],stage1_28[94]}
   );
   gpc606_5 gpc580 (
      {stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173], stage0_28[174]},
      {stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137], stage0_30[138]},
      {stage1_32[23],stage1_31[39],stage1_30[42],stage1_29[65],stage1_28[95]}
   );
   gpc606_5 gpc581 (
      {stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179], stage0_28[180]},
      {stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143], stage0_30[144]},
      {stage1_32[24],stage1_31[40],stage1_30[43],stage1_29[66],stage1_28[96]}
   );
   gpc606_5 gpc582 (
      {stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185], stage0_28[186]},
      {stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149], stage0_30[150]},
      {stage1_32[25],stage1_31[41],stage1_30[44],stage1_29[67],stage1_28[97]}
   );
   gpc606_5 gpc583 (
      {stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191], stage0_28[192]},
      {stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155], stage0_30[156]},
      {stage1_32[26],stage1_31[42],stage1_30[45],stage1_29[68],stage1_28[98]}
   );
   gpc606_5 gpc584 (
      {stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197], stage0_28[198]},
      {stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161], stage0_30[162]},
      {stage1_32[27],stage1_31[43],stage1_30[46],stage1_29[69],stage1_28[99]}
   );
   gpc606_5 gpc585 (
      {stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203], stage0_28[204]},
      {stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167], stage0_30[168]},
      {stage1_32[28],stage1_31[44],stage1_30[47],stage1_29[70],stage1_28[100]}
   );
   gpc606_5 gpc586 (
      {stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209], stage0_28[210]},
      {stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173], stage0_30[174]},
      {stage1_32[29],stage1_31[45],stage1_30[48],stage1_29[71],stage1_28[101]}
   );
   gpc606_5 gpc587 (
      {stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215], stage0_28[216]},
      {stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179], stage0_30[180]},
      {stage1_32[30],stage1_31[46],stage1_30[49],stage1_29[72],stage1_28[102]}
   );
   gpc606_5 gpc588 (
      {stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221], stage0_28[222]},
      {stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185], stage0_30[186]},
      {stage1_32[31],stage1_31[47],stage1_30[50],stage1_29[73],stage1_28[103]}
   );
   gpc606_5 gpc589 (
      {stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227], stage0_28[228]},
      {stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191], stage0_30[192]},
      {stage1_32[32],stage1_31[48],stage1_30[51],stage1_29[74],stage1_28[104]}
   );
   gpc606_5 gpc590 (
      {stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233], stage0_28[234]},
      {stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197], stage0_30[198]},
      {stage1_32[33],stage1_31[49],stage1_30[52],stage1_29[75],stage1_28[105]}
   );
   gpc606_5 gpc591 (
      {stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101], stage0_29[102]},
      {stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5], stage0_31[6], stage0_31[7]},
      {stage1_33[0],stage1_32[34],stage1_31[50],stage1_30[53],stage1_29[76]}
   );
   gpc606_5 gpc592 (
      {stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107], stage0_29[108]},
      {stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11], stage0_31[12], stage0_31[13]},
      {stage1_33[1],stage1_32[35],stage1_31[51],stage1_30[54],stage1_29[77]}
   );
   gpc606_5 gpc593 (
      {stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113], stage0_29[114]},
      {stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17], stage0_31[18], stage0_31[19]},
      {stage1_33[2],stage1_32[36],stage1_31[52],stage1_30[55],stage1_29[78]}
   );
   gpc606_5 gpc594 (
      {stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119], stage0_29[120]},
      {stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23], stage0_31[24], stage0_31[25]},
      {stage1_33[3],stage1_32[37],stage1_31[53],stage1_30[56],stage1_29[79]}
   );
   gpc606_5 gpc595 (
      {stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125], stage0_29[126]},
      {stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29], stage0_31[30], stage0_31[31]},
      {stage1_33[4],stage1_32[38],stage1_31[54],stage1_30[57],stage1_29[80]}
   );
   gpc606_5 gpc596 (
      {stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131], stage0_29[132]},
      {stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35], stage0_31[36], stage0_31[37]},
      {stage1_33[5],stage1_32[39],stage1_31[55],stage1_30[58],stage1_29[81]}
   );
   gpc606_5 gpc597 (
      {stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137], stage0_29[138]},
      {stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41], stage0_31[42], stage0_31[43]},
      {stage1_33[6],stage1_32[40],stage1_31[56],stage1_30[59],stage1_29[82]}
   );
   gpc606_5 gpc598 (
      {stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143], stage0_29[144]},
      {stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47], stage0_31[48], stage0_31[49]},
      {stage1_33[7],stage1_32[41],stage1_31[57],stage1_30[60],stage1_29[83]}
   );
   gpc606_5 gpc599 (
      {stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149], stage0_29[150]},
      {stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53], stage0_31[54], stage0_31[55]},
      {stage1_33[8],stage1_32[42],stage1_31[58],stage1_30[61],stage1_29[84]}
   );
   gpc606_5 gpc600 (
      {stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155], stage0_29[156]},
      {stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59], stage0_31[60], stage0_31[61]},
      {stage1_33[9],stage1_32[43],stage1_31[59],stage1_30[62],stage1_29[85]}
   );
   gpc606_5 gpc601 (
      {stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161], stage0_29[162]},
      {stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65], stage0_31[66], stage0_31[67]},
      {stage1_33[10],stage1_32[44],stage1_31[60],stage1_30[63],stage1_29[86]}
   );
   gpc606_5 gpc602 (
      {stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167], stage0_29[168]},
      {stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71], stage0_31[72], stage0_31[73]},
      {stage1_33[11],stage1_32[45],stage1_31[61],stage1_30[64],stage1_29[87]}
   );
   gpc606_5 gpc603 (
      {stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173], stage0_29[174]},
      {stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77], stage0_31[78], stage0_31[79]},
      {stage1_33[12],stage1_32[46],stage1_31[62],stage1_30[65],stage1_29[88]}
   );
   gpc606_5 gpc604 (
      {stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179], stage0_29[180]},
      {stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83], stage0_31[84], stage0_31[85]},
      {stage1_33[13],stage1_32[47],stage1_31[63],stage1_30[66],stage1_29[89]}
   );
   gpc606_5 gpc605 (
      {stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185], stage0_29[186]},
      {stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89], stage0_31[90], stage0_31[91]},
      {stage1_33[14],stage1_32[48],stage1_31[64],stage1_30[67],stage1_29[90]}
   );
   gpc606_5 gpc606 (
      {stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190], stage0_29[191], stage0_29[192]},
      {stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95], stage0_31[96], stage0_31[97]},
      {stage1_33[15],stage1_32[49],stage1_31[65],stage1_30[68],stage1_29[91]}
   );
   gpc606_5 gpc607 (
      {stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196], stage0_29[197], stage0_29[198]},
      {stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101], stage0_31[102], stage0_31[103]},
      {stage1_33[16],stage1_32[50],stage1_31[66],stage1_30[69],stage1_29[92]}
   );
   gpc606_5 gpc608 (
      {stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202], stage0_29[203], stage0_29[204]},
      {stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107], stage0_31[108], stage0_31[109]},
      {stage1_33[17],stage1_32[51],stage1_31[67],stage1_30[70],stage1_29[93]}
   );
   gpc606_5 gpc609 (
      {stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209], stage0_29[210]},
      {stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113], stage0_31[114], stage0_31[115]},
      {stage1_33[18],stage1_32[52],stage1_31[68],stage1_30[71],stage1_29[94]}
   );
   gpc606_5 gpc610 (
      {stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215], stage0_29[216]},
      {stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119], stage0_31[120], stage0_31[121]},
      {stage1_33[19],stage1_32[53],stage1_31[69],stage1_30[72],stage1_29[95]}
   );
   gpc606_5 gpc611 (
      {stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220], stage0_29[221], stage0_29[222]},
      {stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125], stage0_31[126], stage0_31[127]},
      {stage1_33[20],stage1_32[54],stage1_31[70],stage1_30[73],stage1_29[96]}
   );
   gpc606_5 gpc612 (
      {stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226], stage0_29[227], stage0_29[228]},
      {stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131], stage0_31[132], stage0_31[133]},
      {stage1_33[21],stage1_32[55],stage1_31[71],stage1_30[74],stage1_29[97]}
   );
   gpc606_5 gpc613 (
      {stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232], stage0_29[233], stage0_29[234]},
      {stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137], stage0_31[138], stage0_31[139]},
      {stage1_33[22],stage1_32[56],stage1_31[72],stage1_30[75],stage1_29[98]}
   );
   gpc606_5 gpc614 (
      {stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239], stage0_29[240]},
      {stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143], stage0_31[144], stage0_31[145]},
      {stage1_33[23],stage1_32[57],stage1_31[73],stage1_30[76],stage1_29[99]}
   );
   gpc606_5 gpc615 (
      {stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245], stage0_29[246]},
      {stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149], stage0_31[150], stage0_31[151]},
      {stage1_33[24],stage1_32[58],stage1_31[74],stage1_30[77],stage1_29[100]}
   );
   gpc615_5 gpc616 (
      {stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage0_31[152]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[25],stage1_32[59],stage1_31[75],stage1_30[78]}
   );
   gpc615_5 gpc617 (
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208]},
      {stage0_31[153]},
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage1_34[1],stage1_33[26],stage1_32[60],stage1_31[76],stage1_30[79]}
   );
   gpc615_5 gpc618 (
      {stage0_30[209], stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213]},
      {stage0_31[154]},
      {stage0_32[12], stage0_32[13], stage0_32[14], stage0_32[15], stage0_32[16], stage0_32[17]},
      {stage1_34[2],stage1_33[27],stage1_32[61],stage1_31[77],stage1_30[80]}
   );
   gpc615_5 gpc619 (
      {stage0_30[214], stage0_30[215], stage0_30[216], stage0_30[217], stage0_30[218]},
      {stage0_31[155]},
      {stage0_32[18], stage0_32[19], stage0_32[20], stage0_32[21], stage0_32[22], stage0_32[23]},
      {stage1_34[3],stage1_33[28],stage1_32[62],stage1_31[78],stage1_30[81]}
   );
   gpc615_5 gpc620 (
      {stage0_30[219], stage0_30[220], stage0_30[221], stage0_30[222], stage0_30[223]},
      {stage0_31[156]},
      {stage0_32[24], stage0_32[25], stage0_32[26], stage0_32[27], stage0_32[28], stage0_32[29]},
      {stage1_34[4],stage1_33[29],stage1_32[63],stage1_31[79],stage1_30[82]}
   );
   gpc615_5 gpc621 (
      {stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227], stage0_30[228]},
      {stage0_31[157]},
      {stage0_32[30], stage0_32[31], stage0_32[32], stage0_32[33], stage0_32[34], stage0_32[35]},
      {stage1_34[5],stage1_33[30],stage1_32[64],stage1_31[80],stage1_30[83]}
   );
   gpc615_5 gpc622 (
      {stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage0_31[158]},
      {stage0_32[36], stage0_32[37], stage0_32[38], stage0_32[39], stage0_32[40], stage0_32[41]},
      {stage1_34[6],stage1_33[31],stage1_32[65],stage1_31[81],stage1_30[84]}
   );
   gpc615_5 gpc623 (
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238]},
      {stage0_31[159]},
      {stage0_32[42], stage0_32[43], stage0_32[44], stage0_32[45], stage0_32[46], stage0_32[47]},
      {stage1_34[7],stage1_33[32],stage1_32[66],stage1_31[82],stage1_30[85]}
   );
   gpc615_5 gpc624 (
      {stage0_30[239], stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243]},
      {stage0_31[160]},
      {stage0_32[48], stage0_32[49], stage0_32[50], stage0_32[51], stage0_32[52], stage0_32[53]},
      {stage1_34[8],stage1_33[33],stage1_32[67],stage1_31[83],stage1_30[86]}
   );
   gpc615_5 gpc625 (
      {stage0_30[244], stage0_30[245], stage0_30[246], stage0_30[247], stage0_30[248]},
      {stage0_31[161]},
      {stage0_32[54], stage0_32[55], stage0_32[56], stage0_32[57], stage0_32[58], stage0_32[59]},
      {stage1_34[9],stage1_33[34],stage1_32[68],stage1_31[84],stage1_30[87]}
   );
   gpc615_5 gpc626 (
      {stage0_30[249], stage0_30[250], stage0_30[251], stage0_30[252], stage0_30[253]},
      {stage0_31[162]},
      {stage0_32[60], stage0_32[61], stage0_32[62], stage0_32[63], stage0_32[64], stage0_32[65]},
      {stage1_34[10],stage1_33[35],stage1_32[69],stage1_31[85],stage1_30[88]}
   );
   gpc615_5 gpc627 (
      {stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage0_32[66]},
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage1_35[0],stage1_34[11],stage1_33[36],stage1_32[70],stage1_31[86]}
   );
   gpc615_5 gpc628 (
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172]},
      {stage0_32[67]},
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage1_35[1],stage1_34[12],stage1_33[37],stage1_32[71],stage1_31[87]}
   );
   gpc615_5 gpc629 (
      {stage0_31[173], stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177]},
      {stage0_32[68]},
      {stage0_33[12], stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17]},
      {stage1_35[2],stage1_34[13],stage1_33[38],stage1_32[72],stage1_31[88]}
   );
   gpc615_5 gpc630 (
      {stage0_31[178], stage0_31[179], stage0_31[180], stage0_31[181], stage0_31[182]},
      {stage0_32[69]},
      {stage0_33[18], stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23]},
      {stage1_35[3],stage1_34[14],stage1_33[39],stage1_32[73],stage1_31[89]}
   );
   gpc615_5 gpc631 (
      {stage0_31[183], stage0_31[184], stage0_31[185], stage0_31[186], stage0_31[187]},
      {stage0_32[70]},
      {stage0_33[24], stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29]},
      {stage1_35[4],stage1_34[15],stage1_33[40],stage1_32[74],stage1_31[90]}
   );
   gpc615_5 gpc632 (
      {stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191], stage0_31[192]},
      {stage0_32[71]},
      {stage0_33[30], stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35]},
      {stage1_35[5],stage1_34[16],stage1_33[41],stage1_32[75],stage1_31[91]}
   );
   gpc615_5 gpc633 (
      {stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage0_32[72]},
      {stage0_33[36], stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41]},
      {stage1_35[6],stage1_34[17],stage1_33[42],stage1_32[76],stage1_31[92]}
   );
   gpc615_5 gpc634 (
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202]},
      {stage0_32[73]},
      {stage0_33[42], stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47]},
      {stage1_35[7],stage1_34[18],stage1_33[43],stage1_32[77],stage1_31[93]}
   );
   gpc615_5 gpc635 (
      {stage0_31[203], stage0_31[204], stage0_31[205], stage0_31[206], stage0_31[207]},
      {stage0_32[74]},
      {stage0_33[48], stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52], stage0_33[53]},
      {stage1_35[8],stage1_34[19],stage1_33[44],stage1_32[78],stage1_31[94]}
   );
   gpc615_5 gpc636 (
      {stage0_31[208], stage0_31[209], stage0_31[210], stage0_31[211], stage0_31[212]},
      {stage0_32[75]},
      {stage0_33[54], stage0_33[55], stage0_33[56], stage0_33[57], stage0_33[58], stage0_33[59]},
      {stage1_35[9],stage1_34[20],stage1_33[45],stage1_32[79],stage1_31[95]}
   );
   gpc615_5 gpc637 (
      {stage0_31[213], stage0_31[214], stage0_31[215], stage0_31[216], stage0_31[217]},
      {stage0_32[76]},
      {stage0_33[60], stage0_33[61], stage0_33[62], stage0_33[63], stage0_33[64], stage0_33[65]},
      {stage1_35[10],stage1_34[21],stage1_33[46],stage1_32[80],stage1_31[96]}
   );
   gpc615_5 gpc638 (
      {stage0_31[218], stage0_31[219], stage0_31[220], stage0_31[221], stage0_31[222]},
      {stage0_32[77]},
      {stage0_33[66], stage0_33[67], stage0_33[68], stage0_33[69], stage0_33[70], stage0_33[71]},
      {stage1_35[11],stage1_34[22],stage1_33[47],stage1_32[81],stage1_31[97]}
   );
   gpc615_5 gpc639 (
      {stage0_31[223], stage0_31[224], stage0_31[225], stage0_31[226], stage0_31[227]},
      {stage0_32[78]},
      {stage0_33[72], stage0_33[73], stage0_33[74], stage0_33[75], stage0_33[76], stage0_33[77]},
      {stage1_35[12],stage1_34[23],stage1_33[48],stage1_32[82],stage1_31[98]}
   );
   gpc615_5 gpc640 (
      {stage0_31[228], stage0_31[229], stage0_31[230], stage0_31[231], stage0_31[232]},
      {stage0_32[79]},
      {stage0_33[78], stage0_33[79], stage0_33[80], stage0_33[81], stage0_33[82], stage0_33[83]},
      {stage1_35[13],stage1_34[24],stage1_33[49],stage1_32[83],stage1_31[99]}
   );
   gpc615_5 gpc641 (
      {stage0_31[233], stage0_31[234], stage0_31[235], stage0_31[236], stage0_31[237]},
      {stage0_32[80]},
      {stage0_33[84], stage0_33[85], stage0_33[86], stage0_33[87], stage0_33[88], stage0_33[89]},
      {stage1_35[14],stage1_34[25],stage1_33[50],stage1_32[84],stage1_31[100]}
   );
   gpc615_5 gpc642 (
      {stage0_31[238], stage0_31[239], stage0_31[240], stage0_31[241], stage0_31[242]},
      {stage0_32[81]},
      {stage0_33[90], stage0_33[91], stage0_33[92], stage0_33[93], stage0_33[94], stage0_33[95]},
      {stage1_35[15],stage1_34[26],stage1_33[51],stage1_32[85],stage1_31[101]}
   );
   gpc606_5 gpc643 (
      {stage0_32[82], stage0_32[83], stage0_32[84], stage0_32[85], stage0_32[86], stage0_32[87]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[16],stage1_34[27],stage1_33[52],stage1_32[86]}
   );
   gpc606_5 gpc644 (
      {stage0_32[88], stage0_32[89], stage0_32[90], stage0_32[91], stage0_32[92], stage0_32[93]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[17],stage1_34[28],stage1_33[53],stage1_32[87]}
   );
   gpc606_5 gpc645 (
      {stage0_32[94], stage0_32[95], stage0_32[96], stage0_32[97], stage0_32[98], stage0_32[99]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[18],stage1_34[29],stage1_33[54],stage1_32[88]}
   );
   gpc606_5 gpc646 (
      {stage0_32[100], stage0_32[101], stage0_32[102], stage0_32[103], stage0_32[104], stage0_32[105]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[19],stage1_34[30],stage1_33[55],stage1_32[89]}
   );
   gpc606_5 gpc647 (
      {stage0_32[106], stage0_32[107], stage0_32[108], stage0_32[109], stage0_32[110], stage0_32[111]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[20],stage1_34[31],stage1_33[56],stage1_32[90]}
   );
   gpc606_5 gpc648 (
      {stage0_32[112], stage0_32[113], stage0_32[114], stage0_32[115], stage0_32[116], stage0_32[117]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[21],stage1_34[32],stage1_33[57],stage1_32[91]}
   );
   gpc606_5 gpc649 (
      {stage0_32[118], stage0_32[119], stage0_32[120], stage0_32[121], stage0_32[122], stage0_32[123]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[22],stage1_34[33],stage1_33[58],stage1_32[92]}
   );
   gpc606_5 gpc650 (
      {stage0_32[124], stage0_32[125], stage0_32[126], stage0_32[127], stage0_32[128], stage0_32[129]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[23],stage1_34[34],stage1_33[59],stage1_32[93]}
   );
   gpc606_5 gpc651 (
      {stage0_32[130], stage0_32[131], stage0_32[132], stage0_32[133], stage0_32[134], stage0_32[135]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[24],stage1_34[35],stage1_33[60],stage1_32[94]}
   );
   gpc606_5 gpc652 (
      {stage0_32[136], stage0_32[137], stage0_32[138], stage0_32[139], stage0_32[140], stage0_32[141]},
      {stage0_34[54], stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage1_36[9],stage1_35[25],stage1_34[36],stage1_33[61],stage1_32[95]}
   );
   gpc606_5 gpc653 (
      {stage0_32[142], stage0_32[143], stage0_32[144], stage0_32[145], stage0_32[146], stage0_32[147]},
      {stage0_34[60], stage0_34[61], stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65]},
      {stage1_36[10],stage1_35[26],stage1_34[37],stage1_33[62],stage1_32[96]}
   );
   gpc606_5 gpc654 (
      {stage0_32[148], stage0_32[149], stage0_32[150], stage0_32[151], stage0_32[152], stage0_32[153]},
      {stage0_34[66], stage0_34[67], stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71]},
      {stage1_36[11],stage1_35[27],stage1_34[38],stage1_33[63],stage1_32[97]}
   );
   gpc606_5 gpc655 (
      {stage0_32[154], stage0_32[155], stage0_32[156], stage0_32[157], stage0_32[158], stage0_32[159]},
      {stage0_34[72], stage0_34[73], stage0_34[74], stage0_34[75], stage0_34[76], stage0_34[77]},
      {stage1_36[12],stage1_35[28],stage1_34[39],stage1_33[64],stage1_32[98]}
   );
   gpc606_5 gpc656 (
      {stage0_32[160], stage0_32[161], stage0_32[162], stage0_32[163], stage0_32[164], stage0_32[165]},
      {stage0_34[78], stage0_34[79], stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83]},
      {stage1_36[13],stage1_35[29],stage1_34[40],stage1_33[65],stage1_32[99]}
   );
   gpc606_5 gpc657 (
      {stage0_32[166], stage0_32[167], stage0_32[168], stage0_32[169], stage0_32[170], stage0_32[171]},
      {stage0_34[84], stage0_34[85], stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89]},
      {stage1_36[14],stage1_35[30],stage1_34[41],stage1_33[66],stage1_32[100]}
   );
   gpc606_5 gpc658 (
      {stage0_32[172], stage0_32[173], stage0_32[174], stage0_32[175], stage0_32[176], stage0_32[177]},
      {stage0_34[90], stage0_34[91], stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95]},
      {stage1_36[15],stage1_35[31],stage1_34[42],stage1_33[67],stage1_32[101]}
   );
   gpc606_5 gpc659 (
      {stage0_32[178], stage0_32[179], stage0_32[180], stage0_32[181], stage0_32[182], stage0_32[183]},
      {stage0_34[96], stage0_34[97], stage0_34[98], stage0_34[99], stage0_34[100], stage0_34[101]},
      {stage1_36[16],stage1_35[32],stage1_34[43],stage1_33[68],stage1_32[102]}
   );
   gpc606_5 gpc660 (
      {stage0_32[184], stage0_32[185], stage0_32[186], stage0_32[187], stage0_32[188], stage0_32[189]},
      {stage0_34[102], stage0_34[103], stage0_34[104], stage0_34[105], stage0_34[106], stage0_34[107]},
      {stage1_36[17],stage1_35[33],stage1_34[44],stage1_33[69],stage1_32[103]}
   );
   gpc606_5 gpc661 (
      {stage0_32[190], stage0_32[191], stage0_32[192], stage0_32[193], stage0_32[194], stage0_32[195]},
      {stage0_34[108], stage0_34[109], stage0_34[110], stage0_34[111], stage0_34[112], stage0_34[113]},
      {stage1_36[18],stage1_35[34],stage1_34[45],stage1_33[70],stage1_32[104]}
   );
   gpc606_5 gpc662 (
      {stage0_32[196], stage0_32[197], stage0_32[198], stage0_32[199], stage0_32[200], stage0_32[201]},
      {stage0_34[114], stage0_34[115], stage0_34[116], stage0_34[117], stage0_34[118], stage0_34[119]},
      {stage1_36[19],stage1_35[35],stage1_34[46],stage1_33[71],stage1_32[105]}
   );
   gpc606_5 gpc663 (
      {stage0_32[202], stage0_32[203], stage0_32[204], stage0_32[205], stage0_32[206], stage0_32[207]},
      {stage0_34[120], stage0_34[121], stage0_34[122], stage0_34[123], stage0_34[124], stage0_34[125]},
      {stage1_36[20],stage1_35[36],stage1_34[47],stage1_33[72],stage1_32[106]}
   );
   gpc606_5 gpc664 (
      {stage0_32[208], stage0_32[209], stage0_32[210], stage0_32[211], stage0_32[212], stage0_32[213]},
      {stage0_34[126], stage0_34[127], stage0_34[128], stage0_34[129], stage0_34[130], stage0_34[131]},
      {stage1_36[21],stage1_35[37],stage1_34[48],stage1_33[73],stage1_32[107]}
   );
   gpc606_5 gpc665 (
      {stage0_32[214], stage0_32[215], stage0_32[216], stage0_32[217], stage0_32[218], stage0_32[219]},
      {stage0_34[132], stage0_34[133], stage0_34[134], stage0_34[135], stage0_34[136], stage0_34[137]},
      {stage1_36[22],stage1_35[38],stage1_34[49],stage1_33[74],stage1_32[108]}
   );
   gpc606_5 gpc666 (
      {stage0_32[220], stage0_32[221], stage0_32[222], stage0_32[223], stage0_32[224], stage0_32[225]},
      {stage0_34[138], stage0_34[139], stage0_34[140], stage0_34[141], stage0_34[142], stage0_34[143]},
      {stage1_36[23],stage1_35[39],stage1_34[50],stage1_33[75],stage1_32[109]}
   );
   gpc606_5 gpc667 (
      {stage0_32[226], stage0_32[227], stage0_32[228], stage0_32[229], stage0_32[230], stage0_32[231]},
      {stage0_34[144], stage0_34[145], stage0_34[146], stage0_34[147], stage0_34[148], stage0_34[149]},
      {stage1_36[24],stage1_35[40],stage1_34[51],stage1_33[76],stage1_32[110]}
   );
   gpc606_5 gpc668 (
      {stage0_32[232], stage0_32[233], stage0_32[234], stage0_32[235], stage0_32[236], stage0_32[237]},
      {stage0_34[150], stage0_34[151], stage0_34[152], stage0_34[153], stage0_34[154], stage0_34[155]},
      {stage1_36[25],stage1_35[41],stage1_34[52],stage1_33[77],stage1_32[111]}
   );
   gpc606_5 gpc669 (
      {stage0_32[238], stage0_32[239], stage0_32[240], stage0_32[241], stage0_32[242], stage0_32[243]},
      {stage0_34[156], stage0_34[157], stage0_34[158], stage0_34[159], stage0_34[160], stage0_34[161]},
      {stage1_36[26],stage1_35[42],stage1_34[53],stage1_33[78],stage1_32[112]}
   );
   gpc606_5 gpc670 (
      {stage0_32[244], stage0_32[245], stage0_32[246], stage0_32[247], stage0_32[248], stage0_32[249]},
      {stage0_34[162], stage0_34[163], stage0_34[164], stage0_34[165], stage0_34[166], stage0_34[167]},
      {stage1_36[27],stage1_35[43],stage1_34[54],stage1_33[79],stage1_32[113]}
   );
   gpc606_5 gpc671 (
      {stage0_32[250], stage0_32[251], stage0_32[252], stage0_32[253], stage0_32[254], stage0_32[255]},
      {stage0_34[168], stage0_34[169], stage0_34[170], stage0_34[171], stage0_34[172], stage0_34[173]},
      {stage1_36[28],stage1_35[44],stage1_34[55],stage1_33[80],stage1_32[114]}
   );
   gpc606_5 gpc672 (
      {stage0_33[96], stage0_33[97], stage0_33[98], stage0_33[99], stage0_33[100], stage0_33[101]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[29],stage1_35[45],stage1_34[56],stage1_33[81]}
   );
   gpc606_5 gpc673 (
      {stage0_33[102], stage0_33[103], stage0_33[104], stage0_33[105], stage0_33[106], stage0_33[107]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[30],stage1_35[46],stage1_34[57],stage1_33[82]}
   );
   gpc606_5 gpc674 (
      {stage0_33[108], stage0_33[109], stage0_33[110], stage0_33[111], stage0_33[112], stage0_33[113]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[31],stage1_35[47],stage1_34[58],stage1_33[83]}
   );
   gpc606_5 gpc675 (
      {stage0_33[114], stage0_33[115], stage0_33[116], stage0_33[117], stage0_33[118], stage0_33[119]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[32],stage1_35[48],stage1_34[59],stage1_33[84]}
   );
   gpc606_5 gpc676 (
      {stage0_33[120], stage0_33[121], stage0_33[122], stage0_33[123], stage0_33[124], stage0_33[125]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[33],stage1_35[49],stage1_34[60],stage1_33[85]}
   );
   gpc606_5 gpc677 (
      {stage0_33[126], stage0_33[127], stage0_33[128], stage0_33[129], stage0_33[130], stage0_33[131]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[34],stage1_35[50],stage1_34[61],stage1_33[86]}
   );
   gpc606_5 gpc678 (
      {stage0_33[132], stage0_33[133], stage0_33[134], stage0_33[135], stage0_33[136], stage0_33[137]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[35],stage1_35[51],stage1_34[62],stage1_33[87]}
   );
   gpc606_5 gpc679 (
      {stage0_33[138], stage0_33[139], stage0_33[140], stage0_33[141], stage0_33[142], stage0_33[143]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[36],stage1_35[52],stage1_34[63],stage1_33[88]}
   );
   gpc606_5 gpc680 (
      {stage0_33[144], stage0_33[145], stage0_33[146], stage0_33[147], stage0_33[148], stage0_33[149]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[37],stage1_35[53],stage1_34[64],stage1_33[89]}
   );
   gpc606_5 gpc681 (
      {stage0_33[150], stage0_33[151], stage0_33[152], stage0_33[153], stage0_33[154], stage0_33[155]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[38],stage1_35[54],stage1_34[65],stage1_33[90]}
   );
   gpc606_5 gpc682 (
      {stage0_33[156], stage0_33[157], stage0_33[158], stage0_33[159], stage0_33[160], stage0_33[161]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[39],stage1_35[55],stage1_34[66],stage1_33[91]}
   );
   gpc606_5 gpc683 (
      {stage0_33[162], stage0_33[163], stage0_33[164], stage0_33[165], stage0_33[166], stage0_33[167]},
      {stage0_35[66], stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage1_37[11],stage1_36[40],stage1_35[56],stage1_34[67],stage1_33[92]}
   );
   gpc606_5 gpc684 (
      {stage0_33[168], stage0_33[169], stage0_33[170], stage0_33[171], stage0_33[172], stage0_33[173]},
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76], stage0_35[77]},
      {stage1_37[12],stage1_36[41],stage1_35[57],stage1_34[68],stage1_33[93]}
   );
   gpc606_5 gpc685 (
      {stage0_33[174], stage0_33[175], stage0_33[176], stage0_33[177], stage0_33[178], stage0_33[179]},
      {stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81], stage0_35[82], stage0_35[83]},
      {stage1_37[13],stage1_36[42],stage1_35[58],stage1_34[69],stage1_33[94]}
   );
   gpc606_5 gpc686 (
      {stage0_33[180], stage0_33[181], stage0_33[182], stage0_33[183], stage0_33[184], stage0_33[185]},
      {stage0_35[84], stage0_35[85], stage0_35[86], stage0_35[87], stage0_35[88], stage0_35[89]},
      {stage1_37[14],stage1_36[43],stage1_35[59],stage1_34[70],stage1_33[95]}
   );
   gpc606_5 gpc687 (
      {stage0_33[186], stage0_33[187], stage0_33[188], stage0_33[189], stage0_33[190], stage0_33[191]},
      {stage0_35[90], stage0_35[91], stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95]},
      {stage1_37[15],stage1_36[44],stage1_35[60],stage1_34[71],stage1_33[96]}
   );
   gpc606_5 gpc688 (
      {stage0_33[192], stage0_33[193], stage0_33[194], stage0_33[195], stage0_33[196], stage0_33[197]},
      {stage0_35[96], stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage1_37[16],stage1_36[45],stage1_35[61],stage1_34[72],stage1_33[97]}
   );
   gpc606_5 gpc689 (
      {stage0_33[198], stage0_33[199], stage0_33[200], stage0_33[201], stage0_33[202], stage0_33[203]},
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106], stage0_35[107]},
      {stage1_37[17],stage1_36[46],stage1_35[62],stage1_34[73],stage1_33[98]}
   );
   gpc606_5 gpc690 (
      {stage0_33[204], stage0_33[205], stage0_33[206], stage0_33[207], stage0_33[208], stage0_33[209]},
      {stage0_35[108], stage0_35[109], stage0_35[110], stage0_35[111], stage0_35[112], stage0_35[113]},
      {stage1_37[18],stage1_36[47],stage1_35[63],stage1_34[74],stage1_33[99]}
   );
   gpc606_5 gpc691 (
      {stage0_33[210], stage0_33[211], stage0_33[212], stage0_33[213], stage0_33[214], stage0_33[215]},
      {stage0_35[114], stage0_35[115], stage0_35[116], stage0_35[117], stage0_35[118], stage0_35[119]},
      {stage1_37[19],stage1_36[48],stage1_35[64],stage1_34[75],stage1_33[100]}
   );
   gpc606_5 gpc692 (
      {stage0_33[216], stage0_33[217], stage0_33[218], stage0_33[219], stage0_33[220], stage0_33[221]},
      {stage0_35[120], stage0_35[121], stage0_35[122], stage0_35[123], stage0_35[124], stage0_35[125]},
      {stage1_37[20],stage1_36[49],stage1_35[65],stage1_34[76],stage1_33[101]}
   );
   gpc606_5 gpc693 (
      {stage0_33[222], stage0_33[223], stage0_33[224], stage0_33[225], stage0_33[226], stage0_33[227]},
      {stage0_35[126], stage0_35[127], stage0_35[128], stage0_35[129], stage0_35[130], stage0_35[131]},
      {stage1_37[21],stage1_36[50],stage1_35[66],stage1_34[77],stage1_33[102]}
   );
   gpc606_5 gpc694 (
      {stage0_33[228], stage0_33[229], stage0_33[230], stage0_33[231], stage0_33[232], stage0_33[233]},
      {stage0_35[132], stage0_35[133], stage0_35[134], stage0_35[135], stage0_35[136], stage0_35[137]},
      {stage1_37[22],stage1_36[51],stage1_35[67],stage1_34[78],stage1_33[103]}
   );
   gpc606_5 gpc695 (
      {stage0_33[234], stage0_33[235], stage0_33[236], stage0_33[237], stage0_33[238], stage0_33[239]},
      {stage0_35[138], stage0_35[139], stage0_35[140], stage0_35[141], stage0_35[142], stage0_35[143]},
      {stage1_37[23],stage1_36[52],stage1_35[68],stage1_34[79],stage1_33[104]}
   );
   gpc606_5 gpc696 (
      {stage0_33[240], stage0_33[241], stage0_33[242], stage0_33[243], stage0_33[244], stage0_33[245]},
      {stage0_35[144], stage0_35[145], stage0_35[146], stage0_35[147], stage0_35[148], stage0_35[149]},
      {stage1_37[24],stage1_36[53],stage1_35[69],stage1_34[80],stage1_33[105]}
   );
   gpc606_5 gpc697 (
      {stage0_33[246], stage0_33[247], stage0_33[248], stage0_33[249], stage0_33[250], stage0_33[251]},
      {stage0_35[150], stage0_35[151], stage0_35[152], stage0_35[153], stage0_35[154], stage0_35[155]},
      {stage1_37[25],stage1_36[54],stage1_35[70],stage1_34[81],stage1_33[106]}
   );
   gpc615_5 gpc698 (
      {stage0_34[174], stage0_34[175], stage0_34[176], stage0_34[177], stage0_34[178]},
      {stage0_35[156]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[26],stage1_36[55],stage1_35[71],stage1_34[82]}
   );
   gpc615_5 gpc699 (
      {stage0_34[179], stage0_34[180], stage0_34[181], stage0_34[182], stage0_34[183]},
      {stage0_35[157]},
      {stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11]},
      {stage1_38[1],stage1_37[27],stage1_36[56],stage1_35[72],stage1_34[83]}
   );
   gpc615_5 gpc700 (
      {stage0_34[184], stage0_34[185], stage0_34[186], stage0_34[187], stage0_34[188]},
      {stage0_35[158]},
      {stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16], stage0_36[17]},
      {stage1_38[2],stage1_37[28],stage1_36[57],stage1_35[73],stage1_34[84]}
   );
   gpc615_5 gpc701 (
      {stage0_34[189], stage0_34[190], stage0_34[191], stage0_34[192], stage0_34[193]},
      {stage0_35[159]},
      {stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21], stage0_36[22], stage0_36[23]},
      {stage1_38[3],stage1_37[29],stage1_36[58],stage1_35[74],stage1_34[85]}
   );
   gpc615_5 gpc702 (
      {stage0_34[194], stage0_34[195], stage0_34[196], stage0_34[197], stage0_34[198]},
      {stage0_35[160]},
      {stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27], stage0_36[28], stage0_36[29]},
      {stage1_38[4],stage1_37[30],stage1_36[59],stage1_35[75],stage1_34[86]}
   );
   gpc615_5 gpc703 (
      {stage0_34[199], stage0_34[200], stage0_34[201], stage0_34[202], stage0_34[203]},
      {stage0_35[161]},
      {stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33], stage0_36[34], stage0_36[35]},
      {stage1_38[5],stage1_37[31],stage1_36[60],stage1_35[76],stage1_34[87]}
   );
   gpc615_5 gpc704 (
      {stage0_34[204], stage0_34[205], stage0_34[206], stage0_34[207], stage0_34[208]},
      {stage0_35[162]},
      {stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39], stage0_36[40], stage0_36[41]},
      {stage1_38[6],stage1_37[32],stage1_36[61],stage1_35[77],stage1_34[88]}
   );
   gpc615_5 gpc705 (
      {stage0_34[209], stage0_34[210], stage0_34[211], stage0_34[212], stage0_34[213]},
      {stage0_35[163]},
      {stage0_36[42], stage0_36[43], stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47]},
      {stage1_38[7],stage1_37[33],stage1_36[62],stage1_35[78],stage1_34[89]}
   );
   gpc615_5 gpc706 (
      {stage0_34[214], stage0_34[215], stage0_34[216], stage0_34[217], stage0_34[218]},
      {stage0_35[164]},
      {stage0_36[48], stage0_36[49], stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53]},
      {stage1_38[8],stage1_37[34],stage1_36[63],stage1_35[79],stage1_34[90]}
   );
   gpc615_5 gpc707 (
      {stage0_34[219], stage0_34[220], stage0_34[221], stage0_34[222], stage0_34[223]},
      {stage0_35[165]},
      {stage0_36[54], stage0_36[55], stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59]},
      {stage1_38[9],stage1_37[35],stage1_36[64],stage1_35[80],stage1_34[91]}
   );
   gpc615_5 gpc708 (
      {stage0_34[224], stage0_34[225], stage0_34[226], stage0_34[227], stage0_34[228]},
      {stage0_35[166]},
      {stage0_36[60], stage0_36[61], stage0_36[62], stage0_36[63], stage0_36[64], stage0_36[65]},
      {stage1_38[10],stage1_37[36],stage1_36[65],stage1_35[81],stage1_34[92]}
   );
   gpc615_5 gpc709 (
      {stage0_34[229], stage0_34[230], stage0_34[231], stage0_34[232], stage0_34[233]},
      {stage0_35[167]},
      {stage0_36[66], stage0_36[67], stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71]},
      {stage1_38[11],stage1_37[37],stage1_36[66],stage1_35[82],stage1_34[93]}
   );
   gpc615_5 gpc710 (
      {stage0_34[234], stage0_34[235], stage0_34[236], stage0_34[237], stage0_34[238]},
      {stage0_35[168]},
      {stage0_36[72], stage0_36[73], stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77]},
      {stage1_38[12],stage1_37[38],stage1_36[67],stage1_35[83],stage1_34[94]}
   );
   gpc615_5 gpc711 (
      {stage0_34[239], stage0_34[240], stage0_34[241], stage0_34[242], stage0_34[243]},
      {stage0_35[169]},
      {stage0_36[78], stage0_36[79], stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83]},
      {stage1_38[13],stage1_37[39],stage1_36[68],stage1_35[84],stage1_34[95]}
   );
   gpc615_5 gpc712 (
      {stage0_34[244], stage0_34[245], stage0_34[246], stage0_34[247], stage0_34[248]},
      {stage0_35[170]},
      {stage0_36[84], stage0_36[85], stage0_36[86], stage0_36[87], stage0_36[88], stage0_36[89]},
      {stage1_38[14],stage1_37[40],stage1_36[69],stage1_35[85],stage1_34[96]}
   );
   gpc615_5 gpc713 (
      {stage0_35[171], stage0_35[172], stage0_35[173], stage0_35[174], stage0_35[175]},
      {stage0_36[90]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[15],stage1_37[41],stage1_36[70],stage1_35[86]}
   );
   gpc615_5 gpc714 (
      {stage0_35[176], stage0_35[177], stage0_35[178], stage0_35[179], stage0_35[180]},
      {stage0_36[91]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[16],stage1_37[42],stage1_36[71],stage1_35[87]}
   );
   gpc615_5 gpc715 (
      {stage0_35[181], stage0_35[182], stage0_35[183], stage0_35[184], stage0_35[185]},
      {stage0_36[92]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[17],stage1_37[43],stage1_36[72],stage1_35[88]}
   );
   gpc615_5 gpc716 (
      {stage0_35[186], stage0_35[187], stage0_35[188], stage0_35[189], stage0_35[190]},
      {stage0_36[93]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[18],stage1_37[44],stage1_36[73],stage1_35[89]}
   );
   gpc615_5 gpc717 (
      {stage0_35[191], stage0_35[192], stage0_35[193], stage0_35[194], stage0_35[195]},
      {stage0_36[94]},
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage1_39[4],stage1_38[19],stage1_37[45],stage1_36[74],stage1_35[90]}
   );
   gpc615_5 gpc718 (
      {stage0_35[196], stage0_35[197], stage0_35[198], stage0_35[199], stage0_35[200]},
      {stage0_36[95]},
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage1_39[5],stage1_38[20],stage1_37[46],stage1_36[75],stage1_35[91]}
   );
   gpc615_5 gpc719 (
      {stage0_35[201], stage0_35[202], stage0_35[203], stage0_35[204], stage0_35[205]},
      {stage0_36[96]},
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage1_39[6],stage1_38[21],stage1_37[47],stage1_36[76],stage1_35[92]}
   );
   gpc615_5 gpc720 (
      {stage0_35[206], stage0_35[207], stage0_35[208], stage0_35[209], stage0_35[210]},
      {stage0_36[97]},
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage1_39[7],stage1_38[22],stage1_37[48],stage1_36[77],stage1_35[93]}
   );
   gpc615_5 gpc721 (
      {stage0_35[211], stage0_35[212], stage0_35[213], stage0_35[214], stage0_35[215]},
      {stage0_36[98]},
      {stage0_37[48], stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53]},
      {stage1_39[8],stage1_38[23],stage1_37[49],stage1_36[78],stage1_35[94]}
   );
   gpc615_5 gpc722 (
      {stage0_35[216], stage0_35[217], stage0_35[218], stage0_35[219], stage0_35[220]},
      {stage0_36[99]},
      {stage0_37[54], stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59]},
      {stage1_39[9],stage1_38[24],stage1_37[50],stage1_36[79],stage1_35[95]}
   );
   gpc615_5 gpc723 (
      {stage0_35[221], stage0_35[222], stage0_35[223], stage0_35[224], stage0_35[225]},
      {stage0_36[100]},
      {stage0_37[60], stage0_37[61], stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65]},
      {stage1_39[10],stage1_38[25],stage1_37[51],stage1_36[80],stage1_35[96]}
   );
   gpc615_5 gpc724 (
      {stage0_35[226], stage0_35[227], stage0_35[228], stage0_35[229], stage0_35[230]},
      {stage0_36[101]},
      {stage0_37[66], stage0_37[67], stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71]},
      {stage1_39[11],stage1_38[26],stage1_37[52],stage1_36[81],stage1_35[97]}
   );
   gpc615_5 gpc725 (
      {stage0_35[231], stage0_35[232], stage0_35[233], stage0_35[234], stage0_35[235]},
      {stage0_36[102]},
      {stage0_37[72], stage0_37[73], stage0_37[74], stage0_37[75], stage0_37[76], stage0_37[77]},
      {stage1_39[12],stage1_38[27],stage1_37[53],stage1_36[82],stage1_35[98]}
   );
   gpc207_4 gpc726 (
      {stage0_36[103], stage0_36[104], stage0_36[105], stage0_36[106], stage0_36[107], stage0_36[108], stage0_36[109]},
      {stage0_38[0], stage0_38[1]},
      {stage1_39[13],stage1_38[28],stage1_37[54],stage1_36[83]}
   );
   gpc606_5 gpc727 (
      {stage0_36[110], stage0_36[111], stage0_36[112], stage0_36[113], stage0_36[114], stage0_36[115]},
      {stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5], stage0_38[6], stage0_38[7]},
      {stage1_40[0],stage1_39[14],stage1_38[29],stage1_37[55],stage1_36[84]}
   );
   gpc606_5 gpc728 (
      {stage0_36[116], stage0_36[117], stage0_36[118], stage0_36[119], stage0_36[120], stage0_36[121]},
      {stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11], stage0_38[12], stage0_38[13]},
      {stage1_40[1],stage1_39[15],stage1_38[30],stage1_37[56],stage1_36[85]}
   );
   gpc606_5 gpc729 (
      {stage0_36[122], stage0_36[123], stage0_36[124], stage0_36[125], stage0_36[126], stage0_36[127]},
      {stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17], stage0_38[18], stage0_38[19]},
      {stage1_40[2],stage1_39[16],stage1_38[31],stage1_37[57],stage1_36[86]}
   );
   gpc606_5 gpc730 (
      {stage0_36[128], stage0_36[129], stage0_36[130], stage0_36[131], stage0_36[132], stage0_36[133]},
      {stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23], stage0_38[24], stage0_38[25]},
      {stage1_40[3],stage1_39[17],stage1_38[32],stage1_37[58],stage1_36[87]}
   );
   gpc606_5 gpc731 (
      {stage0_36[134], stage0_36[135], stage0_36[136], stage0_36[137], stage0_36[138], stage0_36[139]},
      {stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29], stage0_38[30], stage0_38[31]},
      {stage1_40[4],stage1_39[18],stage1_38[33],stage1_37[59],stage1_36[88]}
   );
   gpc606_5 gpc732 (
      {stage0_36[140], stage0_36[141], stage0_36[142], stage0_36[143], stage0_36[144], stage0_36[145]},
      {stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35], stage0_38[36], stage0_38[37]},
      {stage1_40[5],stage1_39[19],stage1_38[34],stage1_37[60],stage1_36[89]}
   );
   gpc606_5 gpc733 (
      {stage0_36[146], stage0_36[147], stage0_36[148], stage0_36[149], stage0_36[150], stage0_36[151]},
      {stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41], stage0_38[42], stage0_38[43]},
      {stage1_40[6],stage1_39[20],stage1_38[35],stage1_37[61],stage1_36[90]}
   );
   gpc606_5 gpc734 (
      {stage0_36[152], stage0_36[153], stage0_36[154], stage0_36[155], stage0_36[156], stage0_36[157]},
      {stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47], stage0_38[48], stage0_38[49]},
      {stage1_40[7],stage1_39[21],stage1_38[36],stage1_37[62],stage1_36[91]}
   );
   gpc606_5 gpc735 (
      {stage0_36[158], stage0_36[159], stage0_36[160], stage0_36[161], stage0_36[162], stage0_36[163]},
      {stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53], stage0_38[54], stage0_38[55]},
      {stage1_40[8],stage1_39[22],stage1_38[37],stage1_37[63],stage1_36[92]}
   );
   gpc606_5 gpc736 (
      {stage0_36[164], stage0_36[165], stage0_36[166], stage0_36[167], stage0_36[168], stage0_36[169]},
      {stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59], stage0_38[60], stage0_38[61]},
      {stage1_40[9],stage1_39[23],stage1_38[38],stage1_37[64],stage1_36[93]}
   );
   gpc606_5 gpc737 (
      {stage0_36[170], stage0_36[171], stage0_36[172], stage0_36[173], stage0_36[174], stage0_36[175]},
      {stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65], stage0_38[66], stage0_38[67]},
      {stage1_40[10],stage1_39[24],stage1_38[39],stage1_37[65],stage1_36[94]}
   );
   gpc606_5 gpc738 (
      {stage0_36[176], stage0_36[177], stage0_36[178], stage0_36[179], stage0_36[180], stage0_36[181]},
      {stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71], stage0_38[72], stage0_38[73]},
      {stage1_40[11],stage1_39[25],stage1_38[40],stage1_37[66],stage1_36[95]}
   );
   gpc606_5 gpc739 (
      {stage0_36[182], stage0_36[183], stage0_36[184], stage0_36[185], stage0_36[186], stage0_36[187]},
      {stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77], stage0_38[78], stage0_38[79]},
      {stage1_40[12],stage1_39[26],stage1_38[41],stage1_37[67],stage1_36[96]}
   );
   gpc606_5 gpc740 (
      {stage0_36[188], stage0_36[189], stage0_36[190], stage0_36[191], stage0_36[192], stage0_36[193]},
      {stage0_38[80], stage0_38[81], stage0_38[82], stage0_38[83], stage0_38[84], stage0_38[85]},
      {stage1_40[13],stage1_39[27],stage1_38[42],stage1_37[68],stage1_36[97]}
   );
   gpc606_5 gpc741 (
      {stage0_36[194], stage0_36[195], stage0_36[196], stage0_36[197], stage0_36[198], stage0_36[199]},
      {stage0_38[86], stage0_38[87], stage0_38[88], stage0_38[89], stage0_38[90], stage0_38[91]},
      {stage1_40[14],stage1_39[28],stage1_38[43],stage1_37[69],stage1_36[98]}
   );
   gpc606_5 gpc742 (
      {stage0_36[200], stage0_36[201], stage0_36[202], stage0_36[203], stage0_36[204], stage0_36[205]},
      {stage0_38[92], stage0_38[93], stage0_38[94], stage0_38[95], stage0_38[96], stage0_38[97]},
      {stage1_40[15],stage1_39[29],stage1_38[44],stage1_37[70],stage1_36[99]}
   );
   gpc606_5 gpc743 (
      {stage0_36[206], stage0_36[207], stage0_36[208], stage0_36[209], stage0_36[210], stage0_36[211]},
      {stage0_38[98], stage0_38[99], stage0_38[100], stage0_38[101], stage0_38[102], stage0_38[103]},
      {stage1_40[16],stage1_39[30],stage1_38[45],stage1_37[71],stage1_36[100]}
   );
   gpc606_5 gpc744 (
      {stage0_37[78], stage0_37[79], stage0_37[80], stage0_37[81], stage0_37[82], stage0_37[83]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[17],stage1_39[31],stage1_38[46],stage1_37[72]}
   );
   gpc606_5 gpc745 (
      {stage0_37[84], stage0_37[85], stage0_37[86], stage0_37[87], stage0_37[88], stage0_37[89]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[18],stage1_39[32],stage1_38[47],stage1_37[73]}
   );
   gpc606_5 gpc746 (
      {stage0_37[90], stage0_37[91], stage0_37[92], stage0_37[93], stage0_37[94], stage0_37[95]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[19],stage1_39[33],stage1_38[48],stage1_37[74]}
   );
   gpc606_5 gpc747 (
      {stage0_37[96], stage0_37[97], stage0_37[98], stage0_37[99], stage0_37[100], stage0_37[101]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[20],stage1_39[34],stage1_38[49],stage1_37[75]}
   );
   gpc606_5 gpc748 (
      {stage0_37[102], stage0_37[103], stage0_37[104], stage0_37[105], stage0_37[106], stage0_37[107]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[21],stage1_39[35],stage1_38[50],stage1_37[76]}
   );
   gpc606_5 gpc749 (
      {stage0_37[108], stage0_37[109], stage0_37[110], stage0_37[111], stage0_37[112], stage0_37[113]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[22],stage1_39[36],stage1_38[51],stage1_37[77]}
   );
   gpc606_5 gpc750 (
      {stage0_37[114], stage0_37[115], stage0_37[116], stage0_37[117], stage0_37[118], stage0_37[119]},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[23],stage1_39[37],stage1_38[52],stage1_37[78]}
   );
   gpc606_5 gpc751 (
      {stage0_37[120], stage0_37[121], stage0_37[122], stage0_37[123], stage0_37[124], stage0_37[125]},
      {stage0_39[42], stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage1_41[7],stage1_40[24],stage1_39[38],stage1_38[53],stage1_37[79]}
   );
   gpc606_5 gpc752 (
      {stage0_37[126], stage0_37[127], stage0_37[128], stage0_37[129], stage0_37[130], stage0_37[131]},
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52], stage0_39[53]},
      {stage1_41[8],stage1_40[25],stage1_39[39],stage1_38[54],stage1_37[80]}
   );
   gpc606_5 gpc753 (
      {stage0_37[132], stage0_37[133], stage0_37[134], stage0_37[135], stage0_37[136], stage0_37[137]},
      {stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57], stage0_39[58], stage0_39[59]},
      {stage1_41[9],stage1_40[26],stage1_39[40],stage1_38[55],stage1_37[81]}
   );
   gpc606_5 gpc754 (
      {stage0_37[138], stage0_37[139], stage0_37[140], stage0_37[141], stage0_37[142], stage0_37[143]},
      {stage0_39[60], stage0_39[61], stage0_39[62], stage0_39[63], stage0_39[64], stage0_39[65]},
      {stage1_41[10],stage1_40[27],stage1_39[41],stage1_38[56],stage1_37[82]}
   );
   gpc606_5 gpc755 (
      {stage0_37[144], stage0_37[145], stage0_37[146], stage0_37[147], stage0_37[148], stage0_37[149]},
      {stage0_39[66], stage0_39[67], stage0_39[68], stage0_39[69], stage0_39[70], stage0_39[71]},
      {stage1_41[11],stage1_40[28],stage1_39[42],stage1_38[57],stage1_37[83]}
   );
   gpc606_5 gpc756 (
      {stage0_37[150], stage0_37[151], stage0_37[152], stage0_37[153], stage0_37[154], stage0_37[155]},
      {stage0_39[72], stage0_39[73], stage0_39[74], stage0_39[75], stage0_39[76], stage0_39[77]},
      {stage1_41[12],stage1_40[29],stage1_39[43],stage1_38[58],stage1_37[84]}
   );
   gpc606_5 gpc757 (
      {stage0_37[156], stage0_37[157], stage0_37[158], stage0_37[159], stage0_37[160], stage0_37[161]},
      {stage0_39[78], stage0_39[79], stage0_39[80], stage0_39[81], stage0_39[82], stage0_39[83]},
      {stage1_41[13],stage1_40[30],stage1_39[44],stage1_38[59],stage1_37[85]}
   );
   gpc606_5 gpc758 (
      {stage0_37[162], stage0_37[163], stage0_37[164], stage0_37[165], stage0_37[166], stage0_37[167]},
      {stage0_39[84], stage0_39[85], stage0_39[86], stage0_39[87], stage0_39[88], stage0_39[89]},
      {stage1_41[14],stage1_40[31],stage1_39[45],stage1_38[60],stage1_37[86]}
   );
   gpc606_5 gpc759 (
      {stage0_37[168], stage0_37[169], stage0_37[170], stage0_37[171], stage0_37[172], stage0_37[173]},
      {stage0_39[90], stage0_39[91], stage0_39[92], stage0_39[93], stage0_39[94], stage0_39[95]},
      {stage1_41[15],stage1_40[32],stage1_39[46],stage1_38[61],stage1_37[87]}
   );
   gpc606_5 gpc760 (
      {stage0_37[174], stage0_37[175], stage0_37[176], stage0_37[177], stage0_37[178], stage0_37[179]},
      {stage0_39[96], stage0_39[97], stage0_39[98], stage0_39[99], stage0_39[100], stage0_39[101]},
      {stage1_41[16],stage1_40[33],stage1_39[47],stage1_38[62],stage1_37[88]}
   );
   gpc606_5 gpc761 (
      {stage0_37[180], stage0_37[181], stage0_37[182], stage0_37[183], stage0_37[184], stage0_37[185]},
      {stage0_39[102], stage0_39[103], stage0_39[104], stage0_39[105], stage0_39[106], stage0_39[107]},
      {stage1_41[17],stage1_40[34],stage1_39[48],stage1_38[63],stage1_37[89]}
   );
   gpc606_5 gpc762 (
      {stage0_37[186], stage0_37[187], stage0_37[188], stage0_37[189], stage0_37[190], stage0_37[191]},
      {stage0_39[108], stage0_39[109], stage0_39[110], stage0_39[111], stage0_39[112], stage0_39[113]},
      {stage1_41[18],stage1_40[35],stage1_39[49],stage1_38[64],stage1_37[90]}
   );
   gpc606_5 gpc763 (
      {stage0_37[192], stage0_37[193], stage0_37[194], stage0_37[195], stage0_37[196], stage0_37[197]},
      {stage0_39[114], stage0_39[115], stage0_39[116], stage0_39[117], stage0_39[118], stage0_39[119]},
      {stage1_41[19],stage1_40[36],stage1_39[50],stage1_38[65],stage1_37[91]}
   );
   gpc606_5 gpc764 (
      {stage0_37[198], stage0_37[199], stage0_37[200], stage0_37[201], stage0_37[202], stage0_37[203]},
      {stage0_39[120], stage0_39[121], stage0_39[122], stage0_39[123], stage0_39[124], stage0_39[125]},
      {stage1_41[20],stage1_40[37],stage1_39[51],stage1_38[66],stage1_37[92]}
   );
   gpc606_5 gpc765 (
      {stage0_37[204], stage0_37[205], stage0_37[206], stage0_37[207], stage0_37[208], stage0_37[209]},
      {stage0_39[126], stage0_39[127], stage0_39[128], stage0_39[129], stage0_39[130], stage0_39[131]},
      {stage1_41[21],stage1_40[38],stage1_39[52],stage1_38[67],stage1_37[93]}
   );
   gpc606_5 gpc766 (
      {stage0_37[210], stage0_37[211], stage0_37[212], stage0_37[213], stage0_37[214], stage0_37[215]},
      {stage0_39[132], stage0_39[133], stage0_39[134], stage0_39[135], stage0_39[136], stage0_39[137]},
      {stage1_41[22],stage1_40[39],stage1_39[53],stage1_38[68],stage1_37[94]}
   );
   gpc606_5 gpc767 (
      {stage0_37[216], stage0_37[217], stage0_37[218], stage0_37[219], stage0_37[220], stage0_37[221]},
      {stage0_39[138], stage0_39[139], stage0_39[140], stage0_39[141], stage0_39[142], stage0_39[143]},
      {stage1_41[23],stage1_40[40],stage1_39[54],stage1_38[69],stage1_37[95]}
   );
   gpc606_5 gpc768 (
      {stage0_37[222], stage0_37[223], stage0_37[224], stage0_37[225], stage0_37[226], stage0_37[227]},
      {stage0_39[144], stage0_39[145], stage0_39[146], stage0_39[147], stage0_39[148], stage0_39[149]},
      {stage1_41[24],stage1_40[41],stage1_39[55],stage1_38[70],stage1_37[96]}
   );
   gpc606_5 gpc769 (
      {stage0_37[228], stage0_37[229], stage0_37[230], stage0_37[231], stage0_37[232], stage0_37[233]},
      {stage0_39[150], stage0_39[151], stage0_39[152], stage0_39[153], stage0_39[154], stage0_39[155]},
      {stage1_41[25],stage1_40[42],stage1_39[56],stage1_38[71],stage1_37[97]}
   );
   gpc606_5 gpc770 (
      {stage0_37[234], stage0_37[235], stage0_37[236], stage0_37[237], stage0_37[238], stage0_37[239]},
      {stage0_39[156], stage0_39[157], stage0_39[158], stage0_39[159], stage0_39[160], stage0_39[161]},
      {stage1_41[26],stage1_40[43],stage1_39[57],stage1_38[72],stage1_37[98]}
   );
   gpc606_5 gpc771 (
      {stage0_37[240], stage0_37[241], stage0_37[242], stage0_37[243], stage0_37[244], stage0_37[245]},
      {stage0_39[162], stage0_39[163], stage0_39[164], stage0_39[165], stage0_39[166], stage0_39[167]},
      {stage1_41[27],stage1_40[44],stage1_39[58],stage1_38[73],stage1_37[99]}
   );
   gpc606_5 gpc772 (
      {stage0_37[246], stage0_37[247], stage0_37[248], stage0_37[249], stage0_37[250], stage0_37[251]},
      {stage0_39[168], stage0_39[169], stage0_39[170], stage0_39[171], stage0_39[172], stage0_39[173]},
      {stage1_41[28],stage1_40[45],stage1_39[59],stage1_38[74],stage1_37[100]}
   );
   gpc615_5 gpc773 (
      {stage0_38[104], stage0_38[105], stage0_38[106], stage0_38[107], stage0_38[108]},
      {stage0_39[174]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[29],stage1_40[46],stage1_39[60],stage1_38[75]}
   );
   gpc615_5 gpc774 (
      {stage0_38[109], stage0_38[110], stage0_38[111], stage0_38[112], stage0_38[113]},
      {stage0_39[175]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[30],stage1_40[47],stage1_39[61],stage1_38[76]}
   );
   gpc615_5 gpc775 (
      {stage0_38[114], stage0_38[115], stage0_38[116], stage0_38[117], stage0_38[118]},
      {stage0_39[176]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[31],stage1_40[48],stage1_39[62],stage1_38[77]}
   );
   gpc615_5 gpc776 (
      {stage0_38[119], stage0_38[120], stage0_38[121], stage0_38[122], stage0_38[123]},
      {stage0_39[177]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[32],stage1_40[49],stage1_39[63],stage1_38[78]}
   );
   gpc615_5 gpc777 (
      {stage0_38[124], stage0_38[125], stage0_38[126], stage0_38[127], stage0_38[128]},
      {stage0_39[178]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[33],stage1_40[50],stage1_39[64],stage1_38[79]}
   );
   gpc615_5 gpc778 (
      {stage0_38[129], stage0_38[130], stage0_38[131], stage0_38[132], stage0_38[133]},
      {stage0_39[179]},
      {stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33], stage0_40[34], stage0_40[35]},
      {stage1_42[5],stage1_41[34],stage1_40[51],stage1_39[65],stage1_38[80]}
   );
   gpc615_5 gpc779 (
      {stage0_38[134], stage0_38[135], stage0_38[136], stage0_38[137], stage0_38[138]},
      {stage0_39[180]},
      {stage0_40[36], stage0_40[37], stage0_40[38], stage0_40[39], stage0_40[40], stage0_40[41]},
      {stage1_42[6],stage1_41[35],stage1_40[52],stage1_39[66],stage1_38[81]}
   );
   gpc615_5 gpc780 (
      {stage0_38[139], stage0_38[140], stage0_38[141], stage0_38[142], stage0_38[143]},
      {stage0_39[181]},
      {stage0_40[42], stage0_40[43], stage0_40[44], stage0_40[45], stage0_40[46], stage0_40[47]},
      {stage1_42[7],stage1_41[36],stage1_40[53],stage1_39[67],stage1_38[82]}
   );
   gpc615_5 gpc781 (
      {stage0_38[144], stage0_38[145], stage0_38[146], stage0_38[147], stage0_38[148]},
      {stage0_39[182]},
      {stage0_40[48], stage0_40[49], stage0_40[50], stage0_40[51], stage0_40[52], stage0_40[53]},
      {stage1_42[8],stage1_41[37],stage1_40[54],stage1_39[68],stage1_38[83]}
   );
   gpc615_5 gpc782 (
      {stage0_38[149], stage0_38[150], stage0_38[151], stage0_38[152], stage0_38[153]},
      {stage0_39[183]},
      {stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57], stage0_40[58], stage0_40[59]},
      {stage1_42[9],stage1_41[38],stage1_40[55],stage1_39[69],stage1_38[84]}
   );
   gpc615_5 gpc783 (
      {stage0_38[154], stage0_38[155], stage0_38[156], stage0_38[157], stage0_38[158]},
      {stage0_39[184]},
      {stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63], stage0_40[64], stage0_40[65]},
      {stage1_42[10],stage1_41[39],stage1_40[56],stage1_39[70],stage1_38[85]}
   );
   gpc615_5 gpc784 (
      {stage0_38[159], stage0_38[160], stage0_38[161], stage0_38[162], stage0_38[163]},
      {stage0_39[185]},
      {stage0_40[66], stage0_40[67], stage0_40[68], stage0_40[69], stage0_40[70], stage0_40[71]},
      {stage1_42[11],stage1_41[40],stage1_40[57],stage1_39[71],stage1_38[86]}
   );
   gpc615_5 gpc785 (
      {stage0_38[164], stage0_38[165], stage0_38[166], stage0_38[167], stage0_38[168]},
      {stage0_39[186]},
      {stage0_40[72], stage0_40[73], stage0_40[74], stage0_40[75], stage0_40[76], stage0_40[77]},
      {stage1_42[12],stage1_41[41],stage1_40[58],stage1_39[72],stage1_38[87]}
   );
   gpc615_5 gpc786 (
      {stage0_38[169], stage0_38[170], stage0_38[171], stage0_38[172], stage0_38[173]},
      {stage0_39[187]},
      {stage0_40[78], stage0_40[79], stage0_40[80], stage0_40[81], stage0_40[82], stage0_40[83]},
      {stage1_42[13],stage1_41[42],stage1_40[59],stage1_39[73],stage1_38[88]}
   );
   gpc615_5 gpc787 (
      {stage0_38[174], stage0_38[175], stage0_38[176], stage0_38[177], stage0_38[178]},
      {stage0_39[188]},
      {stage0_40[84], stage0_40[85], stage0_40[86], stage0_40[87], stage0_40[88], stage0_40[89]},
      {stage1_42[14],stage1_41[43],stage1_40[60],stage1_39[74],stage1_38[89]}
   );
   gpc615_5 gpc788 (
      {stage0_38[179], stage0_38[180], stage0_38[181], stage0_38[182], stage0_38[183]},
      {stage0_39[189]},
      {stage0_40[90], stage0_40[91], stage0_40[92], stage0_40[93], stage0_40[94], stage0_40[95]},
      {stage1_42[15],stage1_41[44],stage1_40[61],stage1_39[75],stage1_38[90]}
   );
   gpc615_5 gpc789 (
      {stage0_38[184], stage0_38[185], stage0_38[186], stage0_38[187], stage0_38[188]},
      {stage0_39[190]},
      {stage0_40[96], stage0_40[97], stage0_40[98], stage0_40[99], stage0_40[100], stage0_40[101]},
      {stage1_42[16],stage1_41[45],stage1_40[62],stage1_39[76],stage1_38[91]}
   );
   gpc615_5 gpc790 (
      {stage0_38[189], stage0_38[190], stage0_38[191], stage0_38[192], stage0_38[193]},
      {stage0_39[191]},
      {stage0_40[102], stage0_40[103], stage0_40[104], stage0_40[105], stage0_40[106], stage0_40[107]},
      {stage1_42[17],stage1_41[46],stage1_40[63],stage1_39[77],stage1_38[92]}
   );
   gpc615_5 gpc791 (
      {stage0_38[194], stage0_38[195], stage0_38[196], stage0_38[197], stage0_38[198]},
      {stage0_39[192]},
      {stage0_40[108], stage0_40[109], stage0_40[110], stage0_40[111], stage0_40[112], stage0_40[113]},
      {stage1_42[18],stage1_41[47],stage1_40[64],stage1_39[78],stage1_38[93]}
   );
   gpc615_5 gpc792 (
      {stage0_38[199], stage0_38[200], stage0_38[201], stage0_38[202], stage0_38[203]},
      {stage0_39[193]},
      {stage0_40[114], stage0_40[115], stage0_40[116], stage0_40[117], stage0_40[118], stage0_40[119]},
      {stage1_42[19],stage1_41[48],stage1_40[65],stage1_39[79],stage1_38[94]}
   );
   gpc615_5 gpc793 (
      {stage0_38[204], stage0_38[205], stage0_38[206], stage0_38[207], stage0_38[208]},
      {stage0_39[194]},
      {stage0_40[120], stage0_40[121], stage0_40[122], stage0_40[123], stage0_40[124], stage0_40[125]},
      {stage1_42[20],stage1_41[49],stage1_40[66],stage1_39[80],stage1_38[95]}
   );
   gpc615_5 gpc794 (
      {stage0_38[209], stage0_38[210], stage0_38[211], stage0_38[212], stage0_38[213]},
      {stage0_39[195]},
      {stage0_40[126], stage0_40[127], stage0_40[128], stage0_40[129], stage0_40[130], stage0_40[131]},
      {stage1_42[21],stage1_41[50],stage1_40[67],stage1_39[81],stage1_38[96]}
   );
   gpc623_5 gpc795 (
      {stage0_38[214], stage0_38[215], stage0_38[216]},
      {stage0_39[196], stage0_39[197]},
      {stage0_40[132], stage0_40[133], stage0_40[134], stage0_40[135], stage0_40[136], stage0_40[137]},
      {stage1_42[22],stage1_41[51],stage1_40[68],stage1_39[82],stage1_38[97]}
   );
   gpc615_5 gpc796 (
      {stage0_39[198], stage0_39[199], stage0_39[200], stage0_39[201], stage0_39[202]},
      {stage0_40[138]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[23],stage1_41[52],stage1_40[69],stage1_39[83]}
   );
   gpc615_5 gpc797 (
      {stage0_39[203], stage0_39[204], stage0_39[205], stage0_39[206], stage0_39[207]},
      {stage0_40[139]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[24],stage1_41[53],stage1_40[70],stage1_39[84]}
   );
   gpc615_5 gpc798 (
      {stage0_39[208], stage0_39[209], stage0_39[210], stage0_39[211], stage0_39[212]},
      {stage0_40[140]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[25],stage1_41[54],stage1_40[71],stage1_39[85]}
   );
   gpc615_5 gpc799 (
      {stage0_39[213], stage0_39[214], stage0_39[215], stage0_39[216], stage0_39[217]},
      {stage0_40[141]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[26],stage1_41[55],stage1_40[72],stage1_39[86]}
   );
   gpc606_5 gpc800 (
      {stage0_40[142], stage0_40[143], stage0_40[144], stage0_40[145], stage0_40[146], stage0_40[147]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[4],stage1_42[27],stage1_41[56],stage1_40[73]}
   );
   gpc606_5 gpc801 (
      {stage0_40[148], stage0_40[149], stage0_40[150], stage0_40[151], stage0_40[152], stage0_40[153]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[5],stage1_42[28],stage1_41[57],stage1_40[74]}
   );
   gpc606_5 gpc802 (
      {stage0_40[154], stage0_40[155], stage0_40[156], stage0_40[157], stage0_40[158], stage0_40[159]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[6],stage1_42[29],stage1_41[58],stage1_40[75]}
   );
   gpc606_5 gpc803 (
      {stage0_40[160], stage0_40[161], stage0_40[162], stage0_40[163], stage0_40[164], stage0_40[165]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[7],stage1_42[30],stage1_41[59],stage1_40[76]}
   );
   gpc606_5 gpc804 (
      {stage0_40[166], stage0_40[167], stage0_40[168], stage0_40[169], stage0_40[170], stage0_40[171]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[8],stage1_42[31],stage1_41[60],stage1_40[77]}
   );
   gpc606_5 gpc805 (
      {stage0_40[172], stage0_40[173], stage0_40[174], stage0_40[175], stage0_40[176], stage0_40[177]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[9],stage1_42[32],stage1_41[61],stage1_40[78]}
   );
   gpc606_5 gpc806 (
      {stage0_40[178], stage0_40[179], stage0_40[180], stage0_40[181], stage0_40[182], stage0_40[183]},
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage1_44[6],stage1_43[10],stage1_42[33],stage1_41[62],stage1_40[79]}
   );
   gpc606_5 gpc807 (
      {stage0_40[184], stage0_40[185], stage0_40[186], stage0_40[187], stage0_40[188], stage0_40[189]},
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage1_44[7],stage1_43[11],stage1_42[34],stage1_41[63],stage1_40[80]}
   );
   gpc606_5 gpc808 (
      {stage0_40[190], stage0_40[191], stage0_40[192], stage0_40[193], stage0_40[194], stage0_40[195]},
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage1_44[8],stage1_43[12],stage1_42[35],stage1_41[64],stage1_40[81]}
   );
   gpc606_5 gpc809 (
      {stage0_40[196], stage0_40[197], stage0_40[198], stage0_40[199], stage0_40[200], stage0_40[201]},
      {stage0_42[54], stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59]},
      {stage1_44[9],stage1_43[13],stage1_42[36],stage1_41[65],stage1_40[82]}
   );
   gpc606_5 gpc810 (
      {stage0_40[202], stage0_40[203], stage0_40[204], stage0_40[205], stage0_40[206], stage0_40[207]},
      {stage0_42[60], stage0_42[61], stage0_42[62], stage0_42[63], stage0_42[64], stage0_42[65]},
      {stage1_44[10],stage1_43[14],stage1_42[37],stage1_41[66],stage1_40[83]}
   );
   gpc606_5 gpc811 (
      {stage0_40[208], stage0_40[209], stage0_40[210], stage0_40[211], stage0_40[212], stage0_40[213]},
      {stage0_42[66], stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70], stage0_42[71]},
      {stage1_44[11],stage1_43[15],stage1_42[38],stage1_41[67],stage1_40[84]}
   );
   gpc606_5 gpc812 (
      {stage0_40[214], stage0_40[215], stage0_40[216], stage0_40[217], stage0_40[218], stage0_40[219]},
      {stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75], stage0_42[76], stage0_42[77]},
      {stage1_44[12],stage1_43[16],stage1_42[39],stage1_41[68],stage1_40[85]}
   );
   gpc606_5 gpc813 (
      {stage0_40[220], stage0_40[221], stage0_40[222], stage0_40[223], stage0_40[224], stage0_40[225]},
      {stage0_42[78], stage0_42[79], stage0_42[80], stage0_42[81], stage0_42[82], stage0_42[83]},
      {stage1_44[13],stage1_43[17],stage1_42[40],stage1_41[69],stage1_40[86]}
   );
   gpc606_5 gpc814 (
      {stage0_40[226], stage0_40[227], stage0_40[228], stage0_40[229], stage0_40[230], stage0_40[231]},
      {stage0_42[84], stage0_42[85], stage0_42[86], stage0_42[87], stage0_42[88], stage0_42[89]},
      {stage1_44[14],stage1_43[18],stage1_42[41],stage1_41[70],stage1_40[87]}
   );
   gpc606_5 gpc815 (
      {stage0_40[232], stage0_40[233], stage0_40[234], stage0_40[235], stage0_40[236], stage0_40[237]},
      {stage0_42[90], stage0_42[91], stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95]},
      {stage1_44[15],stage1_43[19],stage1_42[42],stage1_41[71],stage1_40[88]}
   );
   gpc606_5 gpc816 (
      {stage0_40[238], stage0_40[239], stage0_40[240], stage0_40[241], stage0_40[242], stage0_40[243]},
      {stage0_42[96], stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100], stage0_42[101]},
      {stage1_44[16],stage1_43[20],stage1_42[43],stage1_41[72],stage1_40[89]}
   );
   gpc606_5 gpc817 (
      {stage0_40[244], stage0_40[245], stage0_40[246], stage0_40[247], stage0_40[248], stage0_40[249]},
      {stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105], stage0_42[106], stage0_42[107]},
      {stage1_44[17],stage1_43[21],stage1_42[44],stage1_41[73],stage1_40[90]}
   );
   gpc606_5 gpc818 (
      {stage0_40[250], stage0_40[251], stage0_40[252], stage0_40[253], stage0_40[254], stage0_40[255]},
      {stage0_42[108], stage0_42[109], stage0_42[110], stage0_42[111], stage0_42[112], stage0_42[113]},
      {stage1_44[18],stage1_43[22],stage1_42[45],stage1_41[74],stage1_40[91]}
   );
   gpc606_5 gpc819 (
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[19],stage1_43[23],stage1_42[46],stage1_41[75]}
   );
   gpc606_5 gpc820 (
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[20],stage1_43[24],stage1_42[47],stage1_41[76]}
   );
   gpc606_5 gpc821 (
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[21],stage1_43[25],stage1_42[48],stage1_41[77]}
   );
   gpc606_5 gpc822 (
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage0_43[18], stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage1_45[3],stage1_44[22],stage1_43[26],stage1_42[49],stage1_41[78]}
   );
   gpc606_5 gpc823 (
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage1_45[4],stage1_44[23],stage1_43[27],stage1_42[50],stage1_41[79]}
   );
   gpc606_5 gpc824 (
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35]},
      {stage1_45[5],stage1_44[24],stage1_43[28],stage1_42[51],stage1_41[80]}
   );
   gpc606_5 gpc825 (
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39], stage0_43[40], stage0_43[41]},
      {stage1_45[6],stage1_44[25],stage1_43[29],stage1_42[52],stage1_41[81]}
   );
   gpc606_5 gpc826 (
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage0_43[42], stage0_43[43], stage0_43[44], stage0_43[45], stage0_43[46], stage0_43[47]},
      {stage1_45[7],stage1_44[26],stage1_43[30],stage1_42[53],stage1_41[82]}
   );
   gpc606_5 gpc827 (
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage0_43[48], stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage1_45[8],stage1_44[27],stage1_43[31],stage1_42[54],stage1_41[83]}
   );
   gpc606_5 gpc828 (
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58], stage0_43[59]},
      {stage1_45[9],stage1_44[28],stage1_43[32],stage1_42[55],stage1_41[84]}
   );
   gpc606_5 gpc829 (
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63], stage0_43[64], stage0_43[65]},
      {stage1_45[10],stage1_44[29],stage1_43[33],stage1_42[56],stage1_41[85]}
   );
   gpc606_5 gpc830 (
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage0_43[66], stage0_43[67], stage0_43[68], stage0_43[69], stage0_43[70], stage0_43[71]},
      {stage1_45[11],stage1_44[30],stage1_43[34],stage1_42[57],stage1_41[86]}
   );
   gpc606_5 gpc831 (
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100], stage0_41[101]},
      {stage0_43[72], stage0_43[73], stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77]},
      {stage1_45[12],stage1_44[31],stage1_43[35],stage1_42[58],stage1_41[87]}
   );
   gpc606_5 gpc832 (
      {stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105], stage0_41[106], stage0_41[107]},
      {stage0_43[78], stage0_43[79], stage0_43[80], stage0_43[81], stage0_43[82], stage0_43[83]},
      {stage1_45[13],stage1_44[32],stage1_43[36],stage1_42[59],stage1_41[88]}
   );
   gpc606_5 gpc833 (
      {stage0_41[108], stage0_41[109], stage0_41[110], stage0_41[111], stage0_41[112], stage0_41[113]},
      {stage0_43[84], stage0_43[85], stage0_43[86], stage0_43[87], stage0_43[88], stage0_43[89]},
      {stage1_45[14],stage1_44[33],stage1_43[37],stage1_42[60],stage1_41[89]}
   );
   gpc606_5 gpc834 (
      {stage0_41[114], stage0_41[115], stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119]},
      {stage0_43[90], stage0_43[91], stage0_43[92], stage0_43[93], stage0_43[94], stage0_43[95]},
      {stage1_45[15],stage1_44[34],stage1_43[38],stage1_42[61],stage1_41[90]}
   );
   gpc606_5 gpc835 (
      {stage0_41[120], stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage0_43[96], stage0_43[97], stage0_43[98], stage0_43[99], stage0_43[100], stage0_43[101]},
      {stage1_45[16],stage1_44[35],stage1_43[39],stage1_42[62],stage1_41[91]}
   );
   gpc606_5 gpc836 (
      {stage0_41[126], stage0_41[127], stage0_41[128], stage0_41[129], stage0_41[130], stage0_41[131]},
      {stage0_43[102], stage0_43[103], stage0_43[104], stage0_43[105], stage0_43[106], stage0_43[107]},
      {stage1_45[17],stage1_44[36],stage1_43[40],stage1_42[63],stage1_41[92]}
   );
   gpc606_5 gpc837 (
      {stage0_41[132], stage0_41[133], stage0_41[134], stage0_41[135], stage0_41[136], stage0_41[137]},
      {stage0_43[108], stage0_43[109], stage0_43[110], stage0_43[111], stage0_43[112], stage0_43[113]},
      {stage1_45[18],stage1_44[37],stage1_43[41],stage1_42[64],stage1_41[93]}
   );
   gpc606_5 gpc838 (
      {stage0_41[138], stage0_41[139], stage0_41[140], stage0_41[141], stage0_41[142], stage0_41[143]},
      {stage0_43[114], stage0_43[115], stage0_43[116], stage0_43[117], stage0_43[118], stage0_43[119]},
      {stage1_45[19],stage1_44[38],stage1_43[42],stage1_42[65],stage1_41[94]}
   );
   gpc615_5 gpc839 (
      {stage0_41[144], stage0_41[145], stage0_41[146], stage0_41[147], stage0_41[148]},
      {stage0_42[114]},
      {stage0_43[120], stage0_43[121], stage0_43[122], stage0_43[123], stage0_43[124], stage0_43[125]},
      {stage1_45[20],stage1_44[39],stage1_43[43],stage1_42[66],stage1_41[95]}
   );
   gpc615_5 gpc840 (
      {stage0_41[149], stage0_41[150], stage0_41[151], stage0_41[152], stage0_41[153]},
      {stage0_42[115]},
      {stage0_43[126], stage0_43[127], stage0_43[128], stage0_43[129], stage0_43[130], stage0_43[131]},
      {stage1_45[21],stage1_44[40],stage1_43[44],stage1_42[67],stage1_41[96]}
   );
   gpc615_5 gpc841 (
      {stage0_41[154], stage0_41[155], stage0_41[156], stage0_41[157], stage0_41[158]},
      {stage0_42[116]},
      {stage0_43[132], stage0_43[133], stage0_43[134], stage0_43[135], stage0_43[136], stage0_43[137]},
      {stage1_45[22],stage1_44[41],stage1_43[45],stage1_42[68],stage1_41[97]}
   );
   gpc615_5 gpc842 (
      {stage0_41[159], stage0_41[160], stage0_41[161], stage0_41[162], stage0_41[163]},
      {stage0_42[117]},
      {stage0_43[138], stage0_43[139], stage0_43[140], stage0_43[141], stage0_43[142], stage0_43[143]},
      {stage1_45[23],stage1_44[42],stage1_43[46],stage1_42[69],stage1_41[98]}
   );
   gpc615_5 gpc843 (
      {stage0_41[164], stage0_41[165], stage0_41[166], stage0_41[167], stage0_41[168]},
      {stage0_42[118]},
      {stage0_43[144], stage0_43[145], stage0_43[146], stage0_43[147], stage0_43[148], stage0_43[149]},
      {stage1_45[24],stage1_44[43],stage1_43[47],stage1_42[70],stage1_41[99]}
   );
   gpc615_5 gpc844 (
      {stage0_41[169], stage0_41[170], stage0_41[171], stage0_41[172], stage0_41[173]},
      {stage0_42[119]},
      {stage0_43[150], stage0_43[151], stage0_43[152], stage0_43[153], stage0_43[154], stage0_43[155]},
      {stage1_45[25],stage1_44[44],stage1_43[48],stage1_42[71],stage1_41[100]}
   );
   gpc615_5 gpc845 (
      {stage0_41[174], stage0_41[175], stage0_41[176], stage0_41[177], stage0_41[178]},
      {stage0_42[120]},
      {stage0_43[156], stage0_43[157], stage0_43[158], stage0_43[159], stage0_43[160], stage0_43[161]},
      {stage1_45[26],stage1_44[45],stage1_43[49],stage1_42[72],stage1_41[101]}
   );
   gpc615_5 gpc846 (
      {stage0_41[179], stage0_41[180], stage0_41[181], stage0_41[182], stage0_41[183]},
      {stage0_42[121]},
      {stage0_43[162], stage0_43[163], stage0_43[164], stage0_43[165], stage0_43[166], stage0_43[167]},
      {stage1_45[27],stage1_44[46],stage1_43[50],stage1_42[73],stage1_41[102]}
   );
   gpc615_5 gpc847 (
      {stage0_41[184], stage0_41[185], stage0_41[186], stage0_41[187], stage0_41[188]},
      {stage0_42[122]},
      {stage0_43[168], stage0_43[169], stage0_43[170], stage0_43[171], stage0_43[172], stage0_43[173]},
      {stage1_45[28],stage1_44[47],stage1_43[51],stage1_42[74],stage1_41[103]}
   );
   gpc615_5 gpc848 (
      {stage0_41[189], stage0_41[190], stage0_41[191], stage0_41[192], stage0_41[193]},
      {stage0_42[123]},
      {stage0_43[174], stage0_43[175], stage0_43[176], stage0_43[177], stage0_43[178], stage0_43[179]},
      {stage1_45[29],stage1_44[48],stage1_43[52],stage1_42[75],stage1_41[104]}
   );
   gpc615_5 gpc849 (
      {stage0_41[194], stage0_41[195], stage0_41[196], stage0_41[197], stage0_41[198]},
      {stage0_42[124]},
      {stage0_43[180], stage0_43[181], stage0_43[182], stage0_43[183], stage0_43[184], stage0_43[185]},
      {stage1_45[30],stage1_44[49],stage1_43[53],stage1_42[76],stage1_41[105]}
   );
   gpc615_5 gpc850 (
      {stage0_41[199], stage0_41[200], stage0_41[201], stage0_41[202], stage0_41[203]},
      {stage0_42[125]},
      {stage0_43[186], stage0_43[187], stage0_43[188], stage0_43[189], stage0_43[190], stage0_43[191]},
      {stage1_45[31],stage1_44[50],stage1_43[54],stage1_42[77],stage1_41[106]}
   );
   gpc615_5 gpc851 (
      {stage0_41[204], stage0_41[205], stage0_41[206], stage0_41[207], stage0_41[208]},
      {stage0_42[126]},
      {stage0_43[192], stage0_43[193], stage0_43[194], stage0_43[195], stage0_43[196], stage0_43[197]},
      {stage1_45[32],stage1_44[51],stage1_43[55],stage1_42[78],stage1_41[107]}
   );
   gpc615_5 gpc852 (
      {stage0_41[209], stage0_41[210], stage0_41[211], stage0_41[212], stage0_41[213]},
      {stage0_42[127]},
      {stage0_43[198], stage0_43[199], stage0_43[200], stage0_43[201], stage0_43[202], stage0_43[203]},
      {stage1_45[33],stage1_44[52],stage1_43[56],stage1_42[79],stage1_41[108]}
   );
   gpc615_5 gpc853 (
      {stage0_41[214], stage0_41[215], stage0_41[216], stage0_41[217], stage0_41[218]},
      {stage0_42[128]},
      {stage0_43[204], stage0_43[205], stage0_43[206], stage0_43[207], stage0_43[208], stage0_43[209]},
      {stage1_45[34],stage1_44[53],stage1_43[57],stage1_42[80],stage1_41[109]}
   );
   gpc615_5 gpc854 (
      {stage0_41[219], stage0_41[220], stage0_41[221], stage0_41[222], stage0_41[223]},
      {stage0_42[129]},
      {stage0_43[210], stage0_43[211], stage0_43[212], stage0_43[213], stage0_43[214], stage0_43[215]},
      {stage1_45[35],stage1_44[54],stage1_43[58],stage1_42[81],stage1_41[110]}
   );
   gpc615_5 gpc855 (
      {stage0_42[130], stage0_42[131], stage0_42[132], stage0_42[133], stage0_42[134]},
      {stage0_43[216]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[36],stage1_44[55],stage1_43[59],stage1_42[82]}
   );
   gpc615_5 gpc856 (
      {stage0_42[135], stage0_42[136], stage0_42[137], stage0_42[138], stage0_42[139]},
      {stage0_43[217]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[37],stage1_44[56],stage1_43[60],stage1_42[83]}
   );
   gpc615_5 gpc857 (
      {stage0_42[140], stage0_42[141], stage0_42[142], stage0_42[143], stage0_42[144]},
      {stage0_43[218]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[38],stage1_44[57],stage1_43[61],stage1_42[84]}
   );
   gpc615_5 gpc858 (
      {stage0_42[145], stage0_42[146], stage0_42[147], stage0_42[148], stage0_42[149]},
      {stage0_43[219]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[39],stage1_44[58],stage1_43[62],stage1_42[85]}
   );
   gpc615_5 gpc859 (
      {stage0_42[150], stage0_42[151], stage0_42[152], stage0_42[153], stage0_42[154]},
      {stage0_43[220]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[40],stage1_44[59],stage1_43[63],stage1_42[86]}
   );
   gpc615_5 gpc860 (
      {stage0_42[155], stage0_42[156], stage0_42[157], stage0_42[158], stage0_42[159]},
      {stage0_43[221]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[41],stage1_44[60],stage1_43[64],stage1_42[87]}
   );
   gpc615_5 gpc861 (
      {stage0_42[160], stage0_42[161], stage0_42[162], stage0_42[163], stage0_42[164]},
      {stage0_43[222]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[42],stage1_44[61],stage1_43[65],stage1_42[88]}
   );
   gpc615_5 gpc862 (
      {stage0_42[165], stage0_42[166], stage0_42[167], stage0_42[168], stage0_42[169]},
      {stage0_43[223]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[43],stage1_44[62],stage1_43[66],stage1_42[89]}
   );
   gpc615_5 gpc863 (
      {stage0_42[170], stage0_42[171], stage0_42[172], stage0_42[173], stage0_42[174]},
      {stage0_43[224]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[44],stage1_44[63],stage1_43[67],stage1_42[90]}
   );
   gpc615_5 gpc864 (
      {stage0_43[225], stage0_43[226], stage0_43[227], stage0_43[228], stage0_43[229]},
      {stage0_44[54]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[9],stage1_45[45],stage1_44[64],stage1_43[68]}
   );
   gpc615_5 gpc865 (
      {stage0_43[230], stage0_43[231], stage0_43[232], stage0_43[233], stage0_43[234]},
      {stage0_44[55]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[10],stage1_45[46],stage1_44[65],stage1_43[69]}
   );
   gpc615_5 gpc866 (
      {stage0_43[235], stage0_43[236], stage0_43[237], stage0_43[238], stage0_43[239]},
      {stage0_44[56]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[11],stage1_45[47],stage1_44[66],stage1_43[70]}
   );
   gpc615_5 gpc867 (
      {stage0_43[240], stage0_43[241], stage0_43[242], stage0_43[243], stage0_43[244]},
      {stage0_44[57]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[12],stage1_45[48],stage1_44[67],stage1_43[71]}
   );
   gpc615_5 gpc868 (
      {stage0_43[245], stage0_43[246], stage0_43[247], stage0_43[248], stage0_43[249]},
      {stage0_44[58]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[13],stage1_45[49],stage1_44[68],stage1_43[72]}
   );
   gpc606_5 gpc869 (
      {stage0_44[59], stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[5],stage1_46[14],stage1_45[50],stage1_44[69]}
   );
   gpc606_5 gpc870 (
      {stage0_44[65], stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[6],stage1_46[15],stage1_45[51],stage1_44[70]}
   );
   gpc606_5 gpc871 (
      {stage0_44[71], stage0_44[72], stage0_44[73], stage0_44[74], stage0_44[75], stage0_44[76]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[7],stage1_46[16],stage1_45[52],stage1_44[71]}
   );
   gpc606_5 gpc872 (
      {stage0_44[77], stage0_44[78], stage0_44[79], stage0_44[80], stage0_44[81], stage0_44[82]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[8],stage1_46[17],stage1_45[53],stage1_44[72]}
   );
   gpc606_5 gpc873 (
      {stage0_44[83], stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[9],stage1_46[18],stage1_45[54],stage1_44[73]}
   );
   gpc606_5 gpc874 (
      {stage0_44[89], stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[10],stage1_46[19],stage1_45[55],stage1_44[74]}
   );
   gpc606_5 gpc875 (
      {stage0_44[95], stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[11],stage1_46[20],stage1_45[56],stage1_44[75]}
   );
   gpc606_5 gpc876 (
      {stage0_44[101], stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[12],stage1_46[21],stage1_45[57],stage1_44[76]}
   );
   gpc606_5 gpc877 (
      {stage0_44[107], stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[13],stage1_46[22],stage1_45[58],stage1_44[77]}
   );
   gpc606_5 gpc878 (
      {stage0_44[113], stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118]},
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage1_48[9],stage1_47[14],stage1_46[23],stage1_45[59],stage1_44[78]}
   );
   gpc606_5 gpc879 (
      {stage0_44[119], stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124]},
      {stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63], stage0_46[64], stage0_46[65]},
      {stage1_48[10],stage1_47[15],stage1_46[24],stage1_45[60],stage1_44[79]}
   );
   gpc606_5 gpc880 (
      {stage0_44[125], stage0_44[126], stage0_44[127], stage0_44[128], stage0_44[129], stage0_44[130]},
      {stage0_46[66], stage0_46[67], stage0_46[68], stage0_46[69], stage0_46[70], stage0_46[71]},
      {stage1_48[11],stage1_47[16],stage1_46[25],stage1_45[61],stage1_44[80]}
   );
   gpc606_5 gpc881 (
      {stage0_44[131], stage0_44[132], stage0_44[133], stage0_44[134], stage0_44[135], stage0_44[136]},
      {stage0_46[72], stage0_46[73], stage0_46[74], stage0_46[75], stage0_46[76], stage0_46[77]},
      {stage1_48[12],stage1_47[17],stage1_46[26],stage1_45[62],stage1_44[81]}
   );
   gpc606_5 gpc882 (
      {stage0_44[137], stage0_44[138], stage0_44[139], stage0_44[140], stage0_44[141], stage0_44[142]},
      {stage0_46[78], stage0_46[79], stage0_46[80], stage0_46[81], stage0_46[82], stage0_46[83]},
      {stage1_48[13],stage1_47[18],stage1_46[27],stage1_45[63],stage1_44[82]}
   );
   gpc606_5 gpc883 (
      {stage0_44[143], stage0_44[144], stage0_44[145], stage0_44[146], stage0_44[147], stage0_44[148]},
      {stage0_46[84], stage0_46[85], stage0_46[86], stage0_46[87], stage0_46[88], stage0_46[89]},
      {stage1_48[14],stage1_47[19],stage1_46[28],stage1_45[64],stage1_44[83]}
   );
   gpc606_5 gpc884 (
      {stage0_44[149], stage0_44[150], stage0_44[151], stage0_44[152], stage0_44[153], stage0_44[154]},
      {stage0_46[90], stage0_46[91], stage0_46[92], stage0_46[93], stage0_46[94], stage0_46[95]},
      {stage1_48[15],stage1_47[20],stage1_46[29],stage1_45[65],stage1_44[84]}
   );
   gpc606_5 gpc885 (
      {stage0_44[155], stage0_44[156], stage0_44[157], stage0_44[158], stage0_44[159], stage0_44[160]},
      {stage0_46[96], stage0_46[97], stage0_46[98], stage0_46[99], stage0_46[100], stage0_46[101]},
      {stage1_48[16],stage1_47[21],stage1_46[30],stage1_45[66],stage1_44[85]}
   );
   gpc606_5 gpc886 (
      {stage0_44[161], stage0_44[162], stage0_44[163], stage0_44[164], stage0_44[165], stage0_44[166]},
      {stage0_46[102], stage0_46[103], stage0_46[104], stage0_46[105], stage0_46[106], stage0_46[107]},
      {stage1_48[17],stage1_47[22],stage1_46[31],stage1_45[67],stage1_44[86]}
   );
   gpc606_5 gpc887 (
      {stage0_44[167], stage0_44[168], stage0_44[169], stage0_44[170], stage0_44[171], stage0_44[172]},
      {stage0_46[108], stage0_46[109], stage0_46[110], stage0_46[111], stage0_46[112], stage0_46[113]},
      {stage1_48[18],stage1_47[23],stage1_46[32],stage1_45[68],stage1_44[87]}
   );
   gpc606_5 gpc888 (
      {stage0_44[173], stage0_44[174], stage0_44[175], stage0_44[176], stage0_44[177], stage0_44[178]},
      {stage0_46[114], stage0_46[115], stage0_46[116], stage0_46[117], stage0_46[118], stage0_46[119]},
      {stage1_48[19],stage1_47[24],stage1_46[33],stage1_45[69],stage1_44[88]}
   );
   gpc606_5 gpc889 (
      {stage0_44[179], stage0_44[180], stage0_44[181], stage0_44[182], stage0_44[183], stage0_44[184]},
      {stage0_46[120], stage0_46[121], stage0_46[122], stage0_46[123], stage0_46[124], stage0_46[125]},
      {stage1_48[20],stage1_47[25],stage1_46[34],stage1_45[70],stage1_44[89]}
   );
   gpc606_5 gpc890 (
      {stage0_44[185], stage0_44[186], stage0_44[187], stage0_44[188], stage0_44[189], stage0_44[190]},
      {stage0_46[126], stage0_46[127], stage0_46[128], stage0_46[129], stage0_46[130], stage0_46[131]},
      {stage1_48[21],stage1_47[26],stage1_46[35],stage1_45[71],stage1_44[90]}
   );
   gpc606_5 gpc891 (
      {stage0_44[191], stage0_44[192], stage0_44[193], stage0_44[194], stage0_44[195], stage0_44[196]},
      {stage0_46[132], stage0_46[133], stage0_46[134], stage0_46[135], stage0_46[136], stage0_46[137]},
      {stage1_48[22],stage1_47[27],stage1_46[36],stage1_45[72],stage1_44[91]}
   );
   gpc606_5 gpc892 (
      {stage0_44[197], stage0_44[198], stage0_44[199], stage0_44[200], stage0_44[201], stage0_44[202]},
      {stage0_46[138], stage0_46[139], stage0_46[140], stage0_46[141], stage0_46[142], stage0_46[143]},
      {stage1_48[23],stage1_47[28],stage1_46[37],stage1_45[73],stage1_44[92]}
   );
   gpc606_5 gpc893 (
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[24],stage1_47[29],stage1_46[38],stage1_45[74]}
   );
   gpc606_5 gpc894 (
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[25],stage1_47[30],stage1_46[39],stage1_45[75]}
   );
   gpc606_5 gpc895 (
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[26],stage1_47[31],stage1_46[40],stage1_45[76]}
   );
   gpc606_5 gpc896 (
      {stage0_45[48], stage0_45[49], stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[27],stage1_47[32],stage1_46[41],stage1_45[77]}
   );
   gpc606_5 gpc897 (
      {stage0_45[54], stage0_45[55], stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[28],stage1_47[33],stage1_46[42],stage1_45[78]}
   );
   gpc606_5 gpc898 (
      {stage0_45[60], stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[29],stage1_47[34],stage1_46[43],stage1_45[79]}
   );
   gpc606_5 gpc899 (
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70], stage0_45[71]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[30],stage1_47[35],stage1_46[44],stage1_45[80]}
   );
   gpc606_5 gpc900 (
      {stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75], stage0_45[76], stage0_45[77]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[31],stage1_47[36],stage1_46[45],stage1_45[81]}
   );
   gpc606_5 gpc901 (
      {stage0_45[78], stage0_45[79], stage0_45[80], stage0_45[81], stage0_45[82], stage0_45[83]},
      {stage0_47[48], stage0_47[49], stage0_47[50], stage0_47[51], stage0_47[52], stage0_47[53]},
      {stage1_49[8],stage1_48[32],stage1_47[37],stage1_46[46],stage1_45[82]}
   );
   gpc606_5 gpc902 (
      {stage0_45[84], stage0_45[85], stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89]},
      {stage0_47[54], stage0_47[55], stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59]},
      {stage1_49[9],stage1_48[33],stage1_47[38],stage1_46[47],stage1_45[83]}
   );
   gpc606_5 gpc903 (
      {stage0_45[90], stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage0_47[60], stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65]},
      {stage1_49[10],stage1_48[34],stage1_47[39],stage1_46[48],stage1_45[84]}
   );
   gpc606_5 gpc904 (
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100], stage0_45[101]},
      {stage0_47[66], stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71]},
      {stage1_49[11],stage1_48[35],stage1_47[40],stage1_46[49],stage1_45[85]}
   );
   gpc606_5 gpc905 (
      {stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105], stage0_45[106], stage0_45[107]},
      {stage0_47[72], stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage1_49[12],stage1_48[36],stage1_47[41],stage1_46[50],stage1_45[86]}
   );
   gpc606_5 gpc906 (
      {stage0_45[108], stage0_45[109], stage0_45[110], stage0_45[111], stage0_45[112], stage0_45[113]},
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82], stage0_47[83]},
      {stage1_49[13],stage1_48[37],stage1_47[42],stage1_46[51],stage1_45[87]}
   );
   gpc606_5 gpc907 (
      {stage0_45[114], stage0_45[115], stage0_45[116], stage0_45[117], stage0_45[118], stage0_45[119]},
      {stage0_47[84], stage0_47[85], stage0_47[86], stage0_47[87], stage0_47[88], stage0_47[89]},
      {stage1_49[14],stage1_48[38],stage1_47[43],stage1_46[52],stage1_45[88]}
   );
   gpc606_5 gpc908 (
      {stage0_45[120], stage0_45[121], stage0_45[122], stage0_45[123], stage0_45[124], stage0_45[125]},
      {stage0_47[90], stage0_47[91], stage0_47[92], stage0_47[93], stage0_47[94], stage0_47[95]},
      {stage1_49[15],stage1_48[39],stage1_47[44],stage1_46[53],stage1_45[89]}
   );
   gpc606_5 gpc909 (
      {stage0_45[126], stage0_45[127], stage0_45[128], stage0_45[129], stage0_45[130], stage0_45[131]},
      {stage0_47[96], stage0_47[97], stage0_47[98], stage0_47[99], stage0_47[100], stage0_47[101]},
      {stage1_49[16],stage1_48[40],stage1_47[45],stage1_46[54],stage1_45[90]}
   );
   gpc606_5 gpc910 (
      {stage0_45[132], stage0_45[133], stage0_45[134], stage0_45[135], stage0_45[136], stage0_45[137]},
      {stage0_47[102], stage0_47[103], stage0_47[104], stage0_47[105], stage0_47[106], stage0_47[107]},
      {stage1_49[17],stage1_48[41],stage1_47[46],stage1_46[55],stage1_45[91]}
   );
   gpc606_5 gpc911 (
      {stage0_45[138], stage0_45[139], stage0_45[140], stage0_45[141], stage0_45[142], stage0_45[143]},
      {stage0_47[108], stage0_47[109], stage0_47[110], stage0_47[111], stage0_47[112], stage0_47[113]},
      {stage1_49[18],stage1_48[42],stage1_47[47],stage1_46[56],stage1_45[92]}
   );
   gpc606_5 gpc912 (
      {stage0_45[144], stage0_45[145], stage0_45[146], stage0_45[147], stage0_45[148], stage0_45[149]},
      {stage0_47[114], stage0_47[115], stage0_47[116], stage0_47[117], stage0_47[118], stage0_47[119]},
      {stage1_49[19],stage1_48[43],stage1_47[48],stage1_46[57],stage1_45[93]}
   );
   gpc606_5 gpc913 (
      {stage0_45[150], stage0_45[151], stage0_45[152], stage0_45[153], stage0_45[154], stage0_45[155]},
      {stage0_47[120], stage0_47[121], stage0_47[122], stage0_47[123], stage0_47[124], stage0_47[125]},
      {stage1_49[20],stage1_48[44],stage1_47[49],stage1_46[58],stage1_45[94]}
   );
   gpc606_5 gpc914 (
      {stage0_45[156], stage0_45[157], stage0_45[158], stage0_45[159], stage0_45[160], stage0_45[161]},
      {stage0_47[126], stage0_47[127], stage0_47[128], stage0_47[129], stage0_47[130], stage0_47[131]},
      {stage1_49[21],stage1_48[45],stage1_47[50],stage1_46[59],stage1_45[95]}
   );
   gpc606_5 gpc915 (
      {stage0_45[162], stage0_45[163], stage0_45[164], stage0_45[165], stage0_45[166], stage0_45[167]},
      {stage0_47[132], stage0_47[133], stage0_47[134], stage0_47[135], stage0_47[136], stage0_47[137]},
      {stage1_49[22],stage1_48[46],stage1_47[51],stage1_46[60],stage1_45[96]}
   );
   gpc606_5 gpc916 (
      {stage0_45[168], stage0_45[169], stage0_45[170], stage0_45[171], stage0_45[172], stage0_45[173]},
      {stage0_47[138], stage0_47[139], stage0_47[140], stage0_47[141], stage0_47[142], stage0_47[143]},
      {stage1_49[23],stage1_48[47],stage1_47[52],stage1_46[61],stage1_45[97]}
   );
   gpc606_5 gpc917 (
      {stage0_45[174], stage0_45[175], stage0_45[176], stage0_45[177], stage0_45[178], stage0_45[179]},
      {stage0_47[144], stage0_47[145], stage0_47[146], stage0_47[147], stage0_47[148], stage0_47[149]},
      {stage1_49[24],stage1_48[48],stage1_47[53],stage1_46[62],stage1_45[98]}
   );
   gpc615_5 gpc918 (
      {stage0_45[180], stage0_45[181], stage0_45[182], stage0_45[183], stage0_45[184]},
      {stage0_46[144]},
      {stage0_47[150], stage0_47[151], stage0_47[152], stage0_47[153], stage0_47[154], stage0_47[155]},
      {stage1_49[25],stage1_48[49],stage1_47[54],stage1_46[63],stage1_45[99]}
   );
   gpc615_5 gpc919 (
      {stage0_45[185], stage0_45[186], stage0_45[187], stage0_45[188], stage0_45[189]},
      {stage0_46[145]},
      {stage0_47[156], stage0_47[157], stage0_47[158], stage0_47[159], stage0_47[160], stage0_47[161]},
      {stage1_49[26],stage1_48[50],stage1_47[55],stage1_46[64],stage1_45[100]}
   );
   gpc615_5 gpc920 (
      {stage0_45[190], stage0_45[191], stage0_45[192], stage0_45[193], stage0_45[194]},
      {stage0_46[146]},
      {stage0_47[162], stage0_47[163], stage0_47[164], stage0_47[165], stage0_47[166], stage0_47[167]},
      {stage1_49[27],stage1_48[51],stage1_47[56],stage1_46[65],stage1_45[101]}
   );
   gpc615_5 gpc921 (
      {stage0_45[195], stage0_45[196], stage0_45[197], stage0_45[198], stage0_45[199]},
      {stage0_46[147]},
      {stage0_47[168], stage0_47[169], stage0_47[170], stage0_47[171], stage0_47[172], stage0_47[173]},
      {stage1_49[28],stage1_48[52],stage1_47[57],stage1_46[66],stage1_45[102]}
   );
   gpc606_5 gpc922 (
      {stage0_46[148], stage0_46[149], stage0_46[150], stage0_46[151], stage0_46[152], stage0_46[153]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[29],stage1_48[53],stage1_47[58],stage1_46[67]}
   );
   gpc606_5 gpc923 (
      {stage0_46[154], stage0_46[155], stage0_46[156], stage0_46[157], stage0_46[158], stage0_46[159]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[30],stage1_48[54],stage1_47[59],stage1_46[68]}
   );
   gpc606_5 gpc924 (
      {stage0_46[160], stage0_46[161], stage0_46[162], stage0_46[163], stage0_46[164], stage0_46[165]},
      {stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17]},
      {stage1_50[2],stage1_49[31],stage1_48[55],stage1_47[60],stage1_46[69]}
   );
   gpc606_5 gpc925 (
      {stage0_46[166], stage0_46[167], stage0_46[168], stage0_46[169], stage0_46[170], stage0_46[171]},
      {stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23]},
      {stage1_50[3],stage1_49[32],stage1_48[56],stage1_47[61],stage1_46[70]}
   );
   gpc606_5 gpc926 (
      {stage0_46[172], stage0_46[173], stage0_46[174], stage0_46[175], stage0_46[176], stage0_46[177]},
      {stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29]},
      {stage1_50[4],stage1_49[33],stage1_48[57],stage1_47[62],stage1_46[71]}
   );
   gpc606_5 gpc927 (
      {stage0_46[178], stage0_46[179], stage0_46[180], stage0_46[181], stage0_46[182], stage0_46[183]},
      {stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33], stage0_48[34], stage0_48[35]},
      {stage1_50[5],stage1_49[34],stage1_48[58],stage1_47[63],stage1_46[72]}
   );
   gpc606_5 gpc928 (
      {stage0_46[184], stage0_46[185], stage0_46[186], stage0_46[187], stage0_46[188], stage0_46[189]},
      {stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41]},
      {stage1_50[6],stage1_49[35],stage1_48[59],stage1_47[64],stage1_46[73]}
   );
   gpc606_5 gpc929 (
      {stage0_46[190], stage0_46[191], stage0_46[192], stage0_46[193], stage0_46[194], stage0_46[195]},
      {stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47]},
      {stage1_50[7],stage1_49[36],stage1_48[60],stage1_47[65],stage1_46[74]}
   );
   gpc606_5 gpc930 (
      {stage0_46[196], stage0_46[197], stage0_46[198], stage0_46[199], stage0_46[200], stage0_46[201]},
      {stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51], stage0_48[52], stage0_48[53]},
      {stage1_50[8],stage1_49[37],stage1_48[61],stage1_47[66],stage1_46[75]}
   );
   gpc606_5 gpc931 (
      {stage0_46[202], stage0_46[203], stage0_46[204], stage0_46[205], stage0_46[206], stage0_46[207]},
      {stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57], stage0_48[58], stage0_48[59]},
      {stage1_50[9],stage1_49[38],stage1_48[62],stage1_47[67],stage1_46[76]}
   );
   gpc606_5 gpc932 (
      {stage0_46[208], stage0_46[209], stage0_46[210], stage0_46[211], stage0_46[212], stage0_46[213]},
      {stage0_48[60], stage0_48[61], stage0_48[62], stage0_48[63], stage0_48[64], stage0_48[65]},
      {stage1_50[10],stage1_49[39],stage1_48[63],stage1_47[68],stage1_46[77]}
   );
   gpc606_5 gpc933 (
      {stage0_46[214], stage0_46[215], stage0_46[216], stage0_46[217], stage0_46[218], stage0_46[219]},
      {stage0_48[66], stage0_48[67], stage0_48[68], stage0_48[69], stage0_48[70], stage0_48[71]},
      {stage1_50[11],stage1_49[40],stage1_48[64],stage1_47[69],stage1_46[78]}
   );
   gpc606_5 gpc934 (
      {stage0_46[220], stage0_46[221], stage0_46[222], stage0_46[223], stage0_46[224], stage0_46[225]},
      {stage0_48[72], stage0_48[73], stage0_48[74], stage0_48[75], stage0_48[76], stage0_48[77]},
      {stage1_50[12],stage1_49[41],stage1_48[65],stage1_47[70],stage1_46[79]}
   );
   gpc606_5 gpc935 (
      {stage0_46[226], stage0_46[227], stage0_46[228], stage0_46[229], stage0_46[230], stage0_46[231]},
      {stage0_48[78], stage0_48[79], stage0_48[80], stage0_48[81], stage0_48[82], stage0_48[83]},
      {stage1_50[13],stage1_49[42],stage1_48[66],stage1_47[71],stage1_46[80]}
   );
   gpc615_5 gpc936 (
      {stage0_46[232], stage0_46[233], stage0_46[234], stage0_46[235], stage0_46[236]},
      {stage0_47[174]},
      {stage0_48[84], stage0_48[85], stage0_48[86], stage0_48[87], stage0_48[88], stage0_48[89]},
      {stage1_50[14],stage1_49[43],stage1_48[67],stage1_47[72],stage1_46[81]}
   );
   gpc615_5 gpc937 (
      {stage0_47[175], stage0_47[176], stage0_47[177], stage0_47[178], stage0_47[179]},
      {stage0_48[90]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[15],stage1_49[44],stage1_48[68],stage1_47[73]}
   );
   gpc615_5 gpc938 (
      {stage0_47[180], stage0_47[181], stage0_47[182], stage0_47[183], stage0_47[184]},
      {stage0_48[91]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[16],stage1_49[45],stage1_48[69],stage1_47[74]}
   );
   gpc615_5 gpc939 (
      {stage0_47[185], stage0_47[186], stage0_47[187], stage0_47[188], stage0_47[189]},
      {stage0_48[92]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[17],stage1_49[46],stage1_48[70],stage1_47[75]}
   );
   gpc615_5 gpc940 (
      {stage0_47[190], stage0_47[191], stage0_47[192], stage0_47[193], stage0_47[194]},
      {stage0_48[93]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[18],stage1_49[47],stage1_48[71],stage1_47[76]}
   );
   gpc615_5 gpc941 (
      {stage0_47[195], stage0_47[196], stage0_47[197], stage0_47[198], stage0_47[199]},
      {stage0_48[94]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[19],stage1_49[48],stage1_48[72],stage1_47[77]}
   );
   gpc615_5 gpc942 (
      {stage0_47[200], stage0_47[201], stage0_47[202], stage0_47[203], stage0_47[204]},
      {stage0_48[95]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[20],stage1_49[49],stage1_48[73],stage1_47[78]}
   );
   gpc606_5 gpc943 (
      {stage0_48[96], stage0_48[97], stage0_48[98], stage0_48[99], stage0_48[100], stage0_48[101]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[6],stage1_50[21],stage1_49[50],stage1_48[74]}
   );
   gpc606_5 gpc944 (
      {stage0_48[102], stage0_48[103], stage0_48[104], stage0_48[105], stage0_48[106], stage0_48[107]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[7],stage1_50[22],stage1_49[51],stage1_48[75]}
   );
   gpc615_5 gpc945 (
      {stage0_48[108], stage0_48[109], stage0_48[110], stage0_48[111], stage0_48[112]},
      {stage0_49[36]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[8],stage1_50[23],stage1_49[52],stage1_48[76]}
   );
   gpc615_5 gpc946 (
      {stage0_48[113], stage0_48[114], stage0_48[115], stage0_48[116], stage0_48[117]},
      {stage0_49[37]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[9],stage1_50[24],stage1_49[53],stage1_48[77]}
   );
   gpc615_5 gpc947 (
      {stage0_48[118], stage0_48[119], stage0_48[120], stage0_48[121], stage0_48[122]},
      {stage0_49[38]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[10],stage1_50[25],stage1_49[54],stage1_48[78]}
   );
   gpc615_5 gpc948 (
      {stage0_48[123], stage0_48[124], stage0_48[125], stage0_48[126], stage0_48[127]},
      {stage0_49[39]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[11],stage1_50[26],stage1_49[55],stage1_48[79]}
   );
   gpc615_5 gpc949 (
      {stage0_48[128], stage0_48[129], stage0_48[130], stage0_48[131], stage0_48[132]},
      {stage0_49[40]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[12],stage1_50[27],stage1_49[56],stage1_48[80]}
   );
   gpc615_5 gpc950 (
      {stage0_48[133], stage0_48[134], stage0_48[135], stage0_48[136], stage0_48[137]},
      {stage0_49[41]},
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47]},
      {stage1_52[7],stage1_51[13],stage1_50[28],stage1_49[57],stage1_48[81]}
   );
   gpc615_5 gpc951 (
      {stage0_48[138], stage0_48[139], stage0_48[140], stage0_48[141], stage0_48[142]},
      {stage0_49[42]},
      {stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53]},
      {stage1_52[8],stage1_51[14],stage1_50[29],stage1_49[58],stage1_48[82]}
   );
   gpc615_5 gpc952 (
      {stage0_48[143], stage0_48[144], stage0_48[145], stage0_48[146], stage0_48[147]},
      {stage0_49[43]},
      {stage0_50[54], stage0_50[55], stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59]},
      {stage1_52[9],stage1_51[15],stage1_50[30],stage1_49[59],stage1_48[83]}
   );
   gpc615_5 gpc953 (
      {stage0_48[148], stage0_48[149], stage0_48[150], stage0_48[151], stage0_48[152]},
      {stage0_49[44]},
      {stage0_50[60], stage0_50[61], stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65]},
      {stage1_52[10],stage1_51[16],stage1_50[31],stage1_49[60],stage1_48[84]}
   );
   gpc615_5 gpc954 (
      {stage0_48[153], stage0_48[154], stage0_48[155], stage0_48[156], stage0_48[157]},
      {stage0_49[45]},
      {stage0_50[66], stage0_50[67], stage0_50[68], stage0_50[69], stage0_50[70], stage0_50[71]},
      {stage1_52[11],stage1_51[17],stage1_50[32],stage1_49[61],stage1_48[85]}
   );
   gpc615_5 gpc955 (
      {stage0_48[158], stage0_48[159], stage0_48[160], stage0_48[161], stage0_48[162]},
      {stage0_49[46]},
      {stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75], stage0_50[76], stage0_50[77]},
      {stage1_52[12],stage1_51[18],stage1_50[33],stage1_49[62],stage1_48[86]}
   );
   gpc615_5 gpc956 (
      {stage0_48[163], stage0_48[164], stage0_48[165], stage0_48[166], stage0_48[167]},
      {stage0_49[47]},
      {stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81], stage0_50[82], stage0_50[83]},
      {stage1_52[13],stage1_51[19],stage1_50[34],stage1_49[63],stage1_48[87]}
   );
   gpc615_5 gpc957 (
      {stage0_48[168], stage0_48[169], stage0_48[170], stage0_48[171], stage0_48[172]},
      {stage0_49[48]},
      {stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87], stage0_50[88], stage0_50[89]},
      {stage1_52[14],stage1_51[20],stage1_50[35],stage1_49[64],stage1_48[88]}
   );
   gpc615_5 gpc958 (
      {stage0_48[173], stage0_48[174], stage0_48[175], stage0_48[176], stage0_48[177]},
      {stage0_49[49]},
      {stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93], stage0_50[94], stage0_50[95]},
      {stage1_52[15],stage1_51[21],stage1_50[36],stage1_49[65],stage1_48[89]}
   );
   gpc615_5 gpc959 (
      {stage0_48[178], stage0_48[179], stage0_48[180], stage0_48[181], stage0_48[182]},
      {stage0_49[50]},
      {stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99], stage0_50[100], stage0_50[101]},
      {stage1_52[16],stage1_51[22],stage1_50[37],stage1_49[66],stage1_48[90]}
   );
   gpc615_5 gpc960 (
      {stage0_48[183], stage0_48[184], stage0_48[185], stage0_48[186], stage0_48[187]},
      {stage0_49[51]},
      {stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105], stage0_50[106], stage0_50[107]},
      {stage1_52[17],stage1_51[23],stage1_50[38],stage1_49[67],stage1_48[91]}
   );
   gpc615_5 gpc961 (
      {stage0_48[188], stage0_48[189], stage0_48[190], stage0_48[191], stage0_48[192]},
      {stage0_49[52]},
      {stage0_50[108], stage0_50[109], stage0_50[110], stage0_50[111], stage0_50[112], stage0_50[113]},
      {stage1_52[18],stage1_51[24],stage1_50[39],stage1_49[68],stage1_48[92]}
   );
   gpc615_5 gpc962 (
      {stage0_48[193], stage0_48[194], stage0_48[195], stage0_48[196], stage0_48[197]},
      {stage0_49[53]},
      {stage0_50[114], stage0_50[115], stage0_50[116], stage0_50[117], stage0_50[118], stage0_50[119]},
      {stage1_52[19],stage1_51[25],stage1_50[40],stage1_49[69],stage1_48[93]}
   );
   gpc615_5 gpc963 (
      {stage0_48[198], stage0_48[199], stage0_48[200], stage0_48[201], stage0_48[202]},
      {stage0_49[54]},
      {stage0_50[120], stage0_50[121], stage0_50[122], stage0_50[123], stage0_50[124], stage0_50[125]},
      {stage1_52[20],stage1_51[26],stage1_50[41],stage1_49[70],stage1_48[94]}
   );
   gpc615_5 gpc964 (
      {stage0_48[203], stage0_48[204], stage0_48[205], stage0_48[206], stage0_48[207]},
      {stage0_49[55]},
      {stage0_50[126], stage0_50[127], stage0_50[128], stage0_50[129], stage0_50[130], stage0_50[131]},
      {stage1_52[21],stage1_51[27],stage1_50[42],stage1_49[71],stage1_48[95]}
   );
   gpc615_5 gpc965 (
      {stage0_48[208], stage0_48[209], stage0_48[210], stage0_48[211], stage0_48[212]},
      {stage0_49[56]},
      {stage0_50[132], stage0_50[133], stage0_50[134], stage0_50[135], stage0_50[136], stage0_50[137]},
      {stage1_52[22],stage1_51[28],stage1_50[43],stage1_49[72],stage1_48[96]}
   );
   gpc615_5 gpc966 (
      {stage0_48[213], stage0_48[214], stage0_48[215], stage0_48[216], stage0_48[217]},
      {stage0_49[57]},
      {stage0_50[138], stage0_50[139], stage0_50[140], stage0_50[141], stage0_50[142], stage0_50[143]},
      {stage1_52[23],stage1_51[29],stage1_50[44],stage1_49[73],stage1_48[97]}
   );
   gpc615_5 gpc967 (
      {stage0_48[218], stage0_48[219], stage0_48[220], stage0_48[221], stage0_48[222]},
      {stage0_49[58]},
      {stage0_50[144], stage0_50[145], stage0_50[146], stage0_50[147], stage0_50[148], stage0_50[149]},
      {stage1_52[24],stage1_51[30],stage1_50[45],stage1_49[74],stage1_48[98]}
   );
   gpc615_5 gpc968 (
      {stage0_48[223], stage0_48[224], stage0_48[225], stage0_48[226], stage0_48[227]},
      {stage0_49[59]},
      {stage0_50[150], stage0_50[151], stage0_50[152], stage0_50[153], stage0_50[154], stage0_50[155]},
      {stage1_52[25],stage1_51[31],stage1_50[46],stage1_49[75],stage1_48[99]}
   );
   gpc615_5 gpc969 (
      {stage0_48[228], stage0_48[229], stage0_48[230], stage0_48[231], stage0_48[232]},
      {stage0_49[60]},
      {stage0_50[156], stage0_50[157], stage0_50[158], stage0_50[159], stage0_50[160], stage0_50[161]},
      {stage1_52[26],stage1_51[32],stage1_50[47],stage1_49[76],stage1_48[100]}
   );
   gpc615_5 gpc970 (
      {stage0_48[233], stage0_48[234], stage0_48[235], stage0_48[236], stage0_48[237]},
      {stage0_49[61]},
      {stage0_50[162], stage0_50[163], stage0_50[164], stage0_50[165], stage0_50[166], stage0_50[167]},
      {stage1_52[27],stage1_51[33],stage1_50[48],stage1_49[77],stage1_48[101]}
   );
   gpc615_5 gpc971 (
      {stage0_48[238], stage0_48[239], stage0_48[240], stage0_48[241], stage0_48[242]},
      {stage0_49[62]},
      {stage0_50[168], stage0_50[169], stage0_50[170], stage0_50[171], stage0_50[172], stage0_50[173]},
      {stage1_52[28],stage1_51[34],stage1_50[49],stage1_49[78],stage1_48[102]}
   );
   gpc615_5 gpc972 (
      {stage0_48[243], stage0_48[244], stage0_48[245], stage0_48[246], stage0_48[247]},
      {stage0_49[63]},
      {stage0_50[174], stage0_50[175], stage0_50[176], stage0_50[177], stage0_50[178], stage0_50[179]},
      {stage1_52[29],stage1_51[35],stage1_50[50],stage1_49[79],stage1_48[103]}
   );
   gpc615_5 gpc973 (
      {stage0_48[248], stage0_48[249], stage0_48[250], stage0_48[251], stage0_48[252]},
      {stage0_49[64]},
      {stage0_50[180], stage0_50[181], stage0_50[182], stage0_50[183], stage0_50[184], stage0_50[185]},
      {stage1_52[30],stage1_51[36],stage1_50[51],stage1_49[80],stage1_48[104]}
   );
   gpc606_5 gpc974 (
      {stage0_49[65], stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[31],stage1_51[37],stage1_50[52],stage1_49[81]}
   );
   gpc606_5 gpc975 (
      {stage0_49[71], stage0_49[72], stage0_49[73], stage0_49[74], stage0_49[75], stage0_49[76]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[32],stage1_51[38],stage1_50[53],stage1_49[82]}
   );
   gpc606_5 gpc976 (
      {stage0_49[77], stage0_49[78], stage0_49[79], stage0_49[80], stage0_49[81], stage0_49[82]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[33],stage1_51[39],stage1_50[54],stage1_49[83]}
   );
   gpc606_5 gpc977 (
      {stage0_49[83], stage0_49[84], stage0_49[85], stage0_49[86], stage0_49[87], stage0_49[88]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[34],stage1_51[40],stage1_50[55],stage1_49[84]}
   );
   gpc606_5 gpc978 (
      {stage0_49[89], stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[35],stage1_51[41],stage1_50[56],stage1_49[85]}
   );
   gpc606_5 gpc979 (
      {stage0_49[95], stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[36],stage1_51[42],stage1_50[57],stage1_49[86]}
   );
   gpc606_5 gpc980 (
      {stage0_49[101], stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[37],stage1_51[43],stage1_50[58],stage1_49[87]}
   );
   gpc606_5 gpc981 (
      {stage0_49[107], stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111], stage0_49[112]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[38],stage1_51[44],stage1_50[59],stage1_49[88]}
   );
   gpc606_5 gpc982 (
      {stage0_49[113], stage0_49[114], stage0_49[115], stage0_49[116], stage0_49[117], stage0_49[118]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[39],stage1_51[45],stage1_50[60],stage1_49[89]}
   );
   gpc606_5 gpc983 (
      {stage0_49[119], stage0_49[120], stage0_49[121], stage0_49[122], stage0_49[123], stage0_49[124]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[40],stage1_51[46],stage1_50[61],stage1_49[90]}
   );
   gpc606_5 gpc984 (
      {stage0_49[125], stage0_49[126], stage0_49[127], stage0_49[128], stage0_49[129], stage0_49[130]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[41],stage1_51[47],stage1_50[62],stage1_49[91]}
   );
   gpc606_5 gpc985 (
      {stage0_49[131], stage0_49[132], stage0_49[133], stage0_49[134], stage0_49[135], stage0_49[136]},
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage1_53[11],stage1_52[42],stage1_51[48],stage1_50[63],stage1_49[92]}
   );
   gpc606_5 gpc986 (
      {stage0_49[137], stage0_49[138], stage0_49[139], stage0_49[140], stage0_49[141], stage0_49[142]},
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage1_53[12],stage1_52[43],stage1_51[49],stage1_50[64],stage1_49[93]}
   );
   gpc606_5 gpc987 (
      {stage0_49[143], stage0_49[144], stage0_49[145], stage0_49[146], stage0_49[147], stage0_49[148]},
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage1_53[13],stage1_52[44],stage1_51[50],stage1_50[65],stage1_49[94]}
   );
   gpc606_5 gpc988 (
      {stage0_49[149], stage0_49[150], stage0_49[151], stage0_49[152], stage0_49[153], stage0_49[154]},
      {stage0_51[84], stage0_51[85], stage0_51[86], stage0_51[87], stage0_51[88], stage0_51[89]},
      {stage1_53[14],stage1_52[45],stage1_51[51],stage1_50[66],stage1_49[95]}
   );
   gpc606_5 gpc989 (
      {stage0_49[155], stage0_49[156], stage0_49[157], stage0_49[158], stage0_49[159], stage0_49[160]},
      {stage0_51[90], stage0_51[91], stage0_51[92], stage0_51[93], stage0_51[94], stage0_51[95]},
      {stage1_53[15],stage1_52[46],stage1_51[52],stage1_50[67],stage1_49[96]}
   );
   gpc606_5 gpc990 (
      {stage0_49[161], stage0_49[162], stage0_49[163], stage0_49[164], stage0_49[165], stage0_49[166]},
      {stage0_51[96], stage0_51[97], stage0_51[98], stage0_51[99], stage0_51[100], stage0_51[101]},
      {stage1_53[16],stage1_52[47],stage1_51[53],stage1_50[68],stage1_49[97]}
   );
   gpc606_5 gpc991 (
      {stage0_49[167], stage0_49[168], stage0_49[169], stage0_49[170], stage0_49[171], stage0_49[172]},
      {stage0_51[102], stage0_51[103], stage0_51[104], stage0_51[105], stage0_51[106], stage0_51[107]},
      {stage1_53[17],stage1_52[48],stage1_51[54],stage1_50[69],stage1_49[98]}
   );
   gpc606_5 gpc992 (
      {stage0_49[173], stage0_49[174], stage0_49[175], stage0_49[176], stage0_49[177], stage0_49[178]},
      {stage0_51[108], stage0_51[109], stage0_51[110], stage0_51[111], stage0_51[112], stage0_51[113]},
      {stage1_53[18],stage1_52[49],stage1_51[55],stage1_50[70],stage1_49[99]}
   );
   gpc606_5 gpc993 (
      {stage0_49[179], stage0_49[180], stage0_49[181], stage0_49[182], stage0_49[183], stage0_49[184]},
      {stage0_51[114], stage0_51[115], stage0_51[116], stage0_51[117], stage0_51[118], stage0_51[119]},
      {stage1_53[19],stage1_52[50],stage1_51[56],stage1_50[71],stage1_49[100]}
   );
   gpc606_5 gpc994 (
      {stage0_49[185], stage0_49[186], stage0_49[187], stage0_49[188], stage0_49[189], stage0_49[190]},
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124], stage0_51[125]},
      {stage1_53[20],stage1_52[51],stage1_51[57],stage1_50[72],stage1_49[101]}
   );
   gpc606_5 gpc995 (
      {stage0_49[191], stage0_49[192], stage0_49[193], stage0_49[194], stage0_49[195], stage0_49[196]},
      {stage0_51[126], stage0_51[127], stage0_51[128], stage0_51[129], stage0_51[130], stage0_51[131]},
      {stage1_53[21],stage1_52[52],stage1_51[58],stage1_50[73],stage1_49[102]}
   );
   gpc606_5 gpc996 (
      {stage0_49[197], stage0_49[198], stage0_49[199], stage0_49[200], stage0_49[201], stage0_49[202]},
      {stage0_51[132], stage0_51[133], stage0_51[134], stage0_51[135], stage0_51[136], stage0_51[137]},
      {stage1_53[22],stage1_52[53],stage1_51[59],stage1_50[74],stage1_49[103]}
   );
   gpc606_5 gpc997 (
      {stage0_49[203], stage0_49[204], stage0_49[205], stage0_49[206], stage0_49[207], stage0_49[208]},
      {stage0_51[138], stage0_51[139], stage0_51[140], stage0_51[141], stage0_51[142], stage0_51[143]},
      {stage1_53[23],stage1_52[54],stage1_51[60],stage1_50[75],stage1_49[104]}
   );
   gpc606_5 gpc998 (
      {stage0_50[186], stage0_50[187], stage0_50[188], stage0_50[189], stage0_50[190], stage0_50[191]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[24],stage1_52[55],stage1_51[61],stage1_50[76]}
   );
   gpc606_5 gpc999 (
      {stage0_50[192], stage0_50[193], stage0_50[194], stage0_50[195], stage0_50[196], stage0_50[197]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[25],stage1_52[56],stage1_51[62],stage1_50[77]}
   );
   gpc606_5 gpc1000 (
      {stage0_50[198], stage0_50[199], stage0_50[200], stage0_50[201], stage0_50[202], stage0_50[203]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[26],stage1_52[57],stage1_51[63],stage1_50[78]}
   );
   gpc606_5 gpc1001 (
      {stage0_50[204], stage0_50[205], stage0_50[206], stage0_50[207], stage0_50[208], stage0_50[209]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[27],stage1_52[58],stage1_51[64],stage1_50[79]}
   );
   gpc606_5 gpc1002 (
      {stage0_50[210], stage0_50[211], stage0_50[212], stage0_50[213], stage0_50[214], stage0_50[215]},
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage1_54[4],stage1_53[28],stage1_52[59],stage1_51[65],stage1_50[80]}
   );
   gpc606_5 gpc1003 (
      {stage0_50[216], stage0_50[217], stage0_50[218], stage0_50[219], stage0_50[220], stage0_50[221]},
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage1_54[5],stage1_53[29],stage1_52[60],stage1_51[66],stage1_50[81]}
   );
   gpc606_5 gpc1004 (
      {stage0_50[222], stage0_50[223], stage0_50[224], stage0_50[225], stage0_50[226], stage0_50[227]},
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage1_54[6],stage1_53[30],stage1_52[61],stage1_51[67],stage1_50[82]}
   );
   gpc615_5 gpc1005 (
      {stage0_50[228], stage0_50[229], stage0_50[230], stage0_50[231], stage0_50[232]},
      {stage0_51[144]},
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage1_54[7],stage1_53[31],stage1_52[62],stage1_51[68],stage1_50[83]}
   );
   gpc615_5 gpc1006 (
      {stage0_50[233], stage0_50[234], stage0_50[235], stage0_50[236], stage0_50[237]},
      {stage0_51[145]},
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage1_54[8],stage1_53[32],stage1_52[63],stage1_51[69],stage1_50[84]}
   );
   gpc615_5 gpc1007 (
      {stage0_50[238], stage0_50[239], stage0_50[240], stage0_50[241], stage0_50[242]},
      {stage0_51[146]},
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage1_54[9],stage1_53[33],stage1_52[64],stage1_51[70],stage1_50[85]}
   );
   gpc606_5 gpc1008 (
      {stage0_51[147], stage0_51[148], stage0_51[149], stage0_51[150], stage0_51[151], stage0_51[152]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[10],stage1_53[34],stage1_52[65],stage1_51[71]}
   );
   gpc606_5 gpc1009 (
      {stage0_51[153], stage0_51[154], stage0_51[155], stage0_51[156], stage0_51[157], stage0_51[158]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[11],stage1_53[35],stage1_52[66],stage1_51[72]}
   );
   gpc606_5 gpc1010 (
      {stage0_51[159], stage0_51[160], stage0_51[161], stage0_51[162], stage0_51[163], stage0_51[164]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[12],stage1_53[36],stage1_52[67],stage1_51[73]}
   );
   gpc606_5 gpc1011 (
      {stage0_51[165], stage0_51[166], stage0_51[167], stage0_51[168], stage0_51[169], stage0_51[170]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[13],stage1_53[37],stage1_52[68],stage1_51[74]}
   );
   gpc606_5 gpc1012 (
      {stage0_51[171], stage0_51[172], stage0_51[173], stage0_51[174], stage0_51[175], stage0_51[176]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[14],stage1_53[38],stage1_52[69],stage1_51[75]}
   );
   gpc606_5 gpc1013 (
      {stage0_51[177], stage0_51[178], stage0_51[179], stage0_51[180], stage0_51[181], stage0_51[182]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[15],stage1_53[39],stage1_52[70],stage1_51[76]}
   );
   gpc606_5 gpc1014 (
      {stage0_51[183], stage0_51[184], stage0_51[185], stage0_51[186], stage0_51[187], stage0_51[188]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[16],stage1_53[40],stage1_52[71],stage1_51[77]}
   );
   gpc606_5 gpc1015 (
      {stage0_51[189], stage0_51[190], stage0_51[191], stage0_51[192], stage0_51[193], stage0_51[194]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[17],stage1_53[41],stage1_52[72],stage1_51[78]}
   );
   gpc606_5 gpc1016 (
      {stage0_51[195], stage0_51[196], stage0_51[197], stage0_51[198], stage0_51[199], stage0_51[200]},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[18],stage1_53[42],stage1_52[73],stage1_51[79]}
   );
   gpc606_5 gpc1017 (
      {stage0_51[201], stage0_51[202], stage0_51[203], stage0_51[204], stage0_51[205], stage0_51[206]},
      {stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57], stage0_53[58], stage0_53[59]},
      {stage1_55[9],stage1_54[19],stage1_53[43],stage1_52[74],stage1_51[80]}
   );
   gpc606_5 gpc1018 (
      {stage0_51[207], stage0_51[208], stage0_51[209], stage0_51[210], stage0_51[211], stage0_51[212]},
      {stage0_53[60], stage0_53[61], stage0_53[62], stage0_53[63], stage0_53[64], stage0_53[65]},
      {stage1_55[10],stage1_54[20],stage1_53[44],stage1_52[75],stage1_51[81]}
   );
   gpc606_5 gpc1019 (
      {stage0_51[213], stage0_51[214], stage0_51[215], stage0_51[216], stage0_51[217], stage0_51[218]},
      {stage0_53[66], stage0_53[67], stage0_53[68], stage0_53[69], stage0_53[70], stage0_53[71]},
      {stage1_55[11],stage1_54[21],stage1_53[45],stage1_52[76],stage1_51[82]}
   );
   gpc606_5 gpc1020 (
      {stage0_51[219], stage0_51[220], stage0_51[221], stage0_51[222], stage0_51[223], stage0_51[224]},
      {stage0_53[72], stage0_53[73], stage0_53[74], stage0_53[75], stage0_53[76], stage0_53[77]},
      {stage1_55[12],stage1_54[22],stage1_53[46],stage1_52[77],stage1_51[83]}
   );
   gpc606_5 gpc1021 (
      {stage0_51[225], stage0_51[226], stage0_51[227], stage0_51[228], stage0_51[229], stage0_51[230]},
      {stage0_53[78], stage0_53[79], stage0_53[80], stage0_53[81], stage0_53[82], stage0_53[83]},
      {stage1_55[13],stage1_54[23],stage1_53[47],stage1_52[78],stage1_51[84]}
   );
   gpc615_5 gpc1022 (
      {stage0_51[231], stage0_51[232], stage0_51[233], stage0_51[234], stage0_51[235]},
      {stage0_52[60]},
      {stage0_53[84], stage0_53[85], stage0_53[86], stage0_53[87], stage0_53[88], stage0_53[89]},
      {stage1_55[14],stage1_54[24],stage1_53[48],stage1_52[79],stage1_51[85]}
   );
   gpc606_5 gpc1023 (
      {stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65], stage0_52[66]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[15],stage1_54[25],stage1_53[49],stage1_52[80]}
   );
   gpc606_5 gpc1024 (
      {stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71], stage0_52[72]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[16],stage1_54[26],stage1_53[50],stage1_52[81]}
   );
   gpc606_5 gpc1025 (
      {stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77], stage0_52[78]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[17],stage1_54[27],stage1_53[51],stage1_52[82]}
   );
   gpc606_5 gpc1026 (
      {stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83], stage0_52[84]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[18],stage1_54[28],stage1_53[52],stage1_52[83]}
   );
   gpc606_5 gpc1027 (
      {stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89], stage0_52[90]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[19],stage1_54[29],stage1_53[53],stage1_52[84]}
   );
   gpc606_5 gpc1028 (
      {stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95], stage0_52[96]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[20],stage1_54[30],stage1_53[54],stage1_52[85]}
   );
   gpc606_5 gpc1029 (
      {stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101], stage0_52[102]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[21],stage1_54[31],stage1_53[55],stage1_52[86]}
   );
   gpc606_5 gpc1030 (
      {stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107], stage0_52[108]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[22],stage1_54[32],stage1_53[56],stage1_52[87]}
   );
   gpc606_5 gpc1031 (
      {stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113], stage0_52[114]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[23],stage1_54[33],stage1_53[57],stage1_52[88]}
   );
   gpc606_5 gpc1032 (
      {stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119], stage0_52[120]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[24],stage1_54[34],stage1_53[58],stage1_52[89]}
   );
   gpc606_5 gpc1033 (
      {stage0_52[121], stage0_52[122], stage0_52[123], stage0_52[124], stage0_52[125], stage0_52[126]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[25],stage1_54[35],stage1_53[59],stage1_52[90]}
   );
   gpc606_5 gpc1034 (
      {stage0_52[127], stage0_52[128], stage0_52[129], stage0_52[130], stage0_52[131], stage0_52[132]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[26],stage1_54[36],stage1_53[60],stage1_52[91]}
   );
   gpc606_5 gpc1035 (
      {stage0_52[133], stage0_52[134], stage0_52[135], stage0_52[136], stage0_52[137], stage0_52[138]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[27],stage1_54[37],stage1_53[61],stage1_52[92]}
   );
   gpc606_5 gpc1036 (
      {stage0_52[139], stage0_52[140], stage0_52[141], stage0_52[142], stage0_52[143], stage0_52[144]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[28],stage1_54[38],stage1_53[62],stage1_52[93]}
   );
   gpc606_5 gpc1037 (
      {stage0_52[145], stage0_52[146], stage0_52[147], stage0_52[148], stage0_52[149], stage0_52[150]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87], stage0_54[88], stage0_54[89]},
      {stage1_56[14],stage1_55[29],stage1_54[39],stage1_53[63],stage1_52[94]}
   );
   gpc606_5 gpc1038 (
      {stage0_52[151], stage0_52[152], stage0_52[153], stage0_52[154], stage0_52[155], stage0_52[156]},
      {stage0_54[90], stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95]},
      {stage1_56[15],stage1_55[30],stage1_54[40],stage1_53[64],stage1_52[95]}
   );
   gpc606_5 gpc1039 (
      {stage0_52[157], stage0_52[158], stage0_52[159], stage0_52[160], stage0_52[161], stage0_52[162]},
      {stage0_54[96], stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101]},
      {stage1_56[16],stage1_55[31],stage1_54[41],stage1_53[65],stage1_52[96]}
   );
   gpc606_5 gpc1040 (
      {stage0_52[163], stage0_52[164], stage0_52[165], stage0_52[166], stage0_52[167], stage0_52[168]},
      {stage0_54[102], stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage1_56[17],stage1_55[32],stage1_54[42],stage1_53[66],stage1_52[97]}
   );
   gpc606_5 gpc1041 (
      {stage0_52[169], stage0_52[170], stage0_52[171], stage0_52[172], stage0_52[173], stage0_52[174]},
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112], stage0_54[113]},
      {stage1_56[18],stage1_55[33],stage1_54[43],stage1_53[67],stage1_52[98]}
   );
   gpc606_5 gpc1042 (
      {stage0_52[175], stage0_52[176], stage0_52[177], stage0_52[178], stage0_52[179], stage0_52[180]},
      {stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117], stage0_54[118], stage0_54[119]},
      {stage1_56[19],stage1_55[34],stage1_54[44],stage1_53[68],stage1_52[99]}
   );
   gpc606_5 gpc1043 (
      {stage0_52[181], stage0_52[182], stage0_52[183], stage0_52[184], stage0_52[185], stage0_52[186]},
      {stage0_54[120], stage0_54[121], stage0_54[122], stage0_54[123], stage0_54[124], stage0_54[125]},
      {stage1_56[20],stage1_55[35],stage1_54[45],stage1_53[69],stage1_52[100]}
   );
   gpc606_5 gpc1044 (
      {stage0_52[187], stage0_52[188], stage0_52[189], stage0_52[190], stage0_52[191], stage0_52[192]},
      {stage0_54[126], stage0_54[127], stage0_54[128], stage0_54[129], stage0_54[130], stage0_54[131]},
      {stage1_56[21],stage1_55[36],stage1_54[46],stage1_53[70],stage1_52[101]}
   );
   gpc606_5 gpc1045 (
      {stage0_52[193], stage0_52[194], stage0_52[195], stage0_52[196], stage0_52[197], stage0_52[198]},
      {stage0_54[132], stage0_54[133], stage0_54[134], stage0_54[135], stage0_54[136], stage0_54[137]},
      {stage1_56[22],stage1_55[37],stage1_54[47],stage1_53[71],stage1_52[102]}
   );
   gpc606_5 gpc1046 (
      {stage0_52[199], stage0_52[200], stage0_52[201], stage0_52[202], stage0_52[203], stage0_52[204]},
      {stage0_54[138], stage0_54[139], stage0_54[140], stage0_54[141], stage0_54[142], stage0_54[143]},
      {stage1_56[23],stage1_55[38],stage1_54[48],stage1_53[72],stage1_52[103]}
   );
   gpc606_5 gpc1047 (
      {stage0_52[205], stage0_52[206], stage0_52[207], stage0_52[208], stage0_52[209], stage0_52[210]},
      {stage0_54[144], stage0_54[145], stage0_54[146], stage0_54[147], stage0_54[148], stage0_54[149]},
      {stage1_56[24],stage1_55[39],stage1_54[49],stage1_53[73],stage1_52[104]}
   );
   gpc606_5 gpc1048 (
      {stage0_52[211], stage0_52[212], stage0_52[213], stage0_52[214], stage0_52[215], stage0_52[216]},
      {stage0_54[150], stage0_54[151], stage0_54[152], stage0_54[153], stage0_54[154], stage0_54[155]},
      {stage1_56[25],stage1_55[40],stage1_54[50],stage1_53[74],stage1_52[105]}
   );
   gpc606_5 gpc1049 (
      {stage0_52[217], stage0_52[218], stage0_52[219], stage0_52[220], stage0_52[221], stage0_52[222]},
      {stage0_54[156], stage0_54[157], stage0_54[158], stage0_54[159], stage0_54[160], stage0_54[161]},
      {stage1_56[26],stage1_55[41],stage1_54[51],stage1_53[75],stage1_52[106]}
   );
   gpc606_5 gpc1050 (
      {stage0_53[90], stage0_53[91], stage0_53[92], stage0_53[93], stage0_53[94], stage0_53[95]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[27],stage1_55[42],stage1_54[52],stage1_53[76]}
   );
   gpc606_5 gpc1051 (
      {stage0_53[96], stage0_53[97], stage0_53[98], stage0_53[99], stage0_53[100], stage0_53[101]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[28],stage1_55[43],stage1_54[53],stage1_53[77]}
   );
   gpc606_5 gpc1052 (
      {stage0_53[102], stage0_53[103], stage0_53[104], stage0_53[105], stage0_53[106], stage0_53[107]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[29],stage1_55[44],stage1_54[54],stage1_53[78]}
   );
   gpc606_5 gpc1053 (
      {stage0_53[108], stage0_53[109], stage0_53[110], stage0_53[111], stage0_53[112], stage0_53[113]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[30],stage1_55[45],stage1_54[55],stage1_53[79]}
   );
   gpc606_5 gpc1054 (
      {stage0_53[114], stage0_53[115], stage0_53[116], stage0_53[117], stage0_53[118], stage0_53[119]},
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage1_57[4],stage1_56[31],stage1_55[46],stage1_54[56],stage1_53[80]}
   );
   gpc606_5 gpc1055 (
      {stage0_53[120], stage0_53[121], stage0_53[122], stage0_53[123], stage0_53[124], stage0_53[125]},
      {stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33], stage0_55[34], stage0_55[35]},
      {stage1_57[5],stage1_56[32],stage1_55[47],stage1_54[57],stage1_53[81]}
   );
   gpc606_5 gpc1056 (
      {stage0_53[126], stage0_53[127], stage0_53[128], stage0_53[129], stage0_53[130], stage0_53[131]},
      {stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39], stage0_55[40], stage0_55[41]},
      {stage1_57[6],stage1_56[33],stage1_55[48],stage1_54[58],stage1_53[82]}
   );
   gpc606_5 gpc1057 (
      {stage0_53[132], stage0_53[133], stage0_53[134], stage0_53[135], stage0_53[136], stage0_53[137]},
      {stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45], stage0_55[46], stage0_55[47]},
      {stage1_57[7],stage1_56[34],stage1_55[49],stage1_54[59],stage1_53[83]}
   );
   gpc606_5 gpc1058 (
      {stage0_53[138], stage0_53[139], stage0_53[140], stage0_53[141], stage0_53[142], stage0_53[143]},
      {stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51], stage0_55[52], stage0_55[53]},
      {stage1_57[8],stage1_56[35],stage1_55[50],stage1_54[60],stage1_53[84]}
   );
   gpc606_5 gpc1059 (
      {stage0_53[144], stage0_53[145], stage0_53[146], stage0_53[147], stage0_53[148], stage0_53[149]},
      {stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57], stage0_55[58], stage0_55[59]},
      {stage1_57[9],stage1_56[36],stage1_55[51],stage1_54[61],stage1_53[85]}
   );
   gpc606_5 gpc1060 (
      {stage0_53[150], stage0_53[151], stage0_53[152], stage0_53[153], stage0_53[154], stage0_53[155]},
      {stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63], stage0_55[64], stage0_55[65]},
      {stage1_57[10],stage1_56[37],stage1_55[52],stage1_54[62],stage1_53[86]}
   );
   gpc606_5 gpc1061 (
      {stage0_53[156], stage0_53[157], stage0_53[158], stage0_53[159], stage0_53[160], stage0_53[161]},
      {stage0_55[66], stage0_55[67], stage0_55[68], stage0_55[69], stage0_55[70], stage0_55[71]},
      {stage1_57[11],stage1_56[38],stage1_55[53],stage1_54[63],stage1_53[87]}
   );
   gpc606_5 gpc1062 (
      {stage0_53[162], stage0_53[163], stage0_53[164], stage0_53[165], stage0_53[166], stage0_53[167]},
      {stage0_55[72], stage0_55[73], stage0_55[74], stage0_55[75], stage0_55[76], stage0_55[77]},
      {stage1_57[12],stage1_56[39],stage1_55[54],stage1_54[64],stage1_53[88]}
   );
   gpc606_5 gpc1063 (
      {stage0_53[168], stage0_53[169], stage0_53[170], stage0_53[171], stage0_53[172], stage0_53[173]},
      {stage0_55[78], stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83]},
      {stage1_57[13],stage1_56[40],stage1_55[55],stage1_54[65],stage1_53[89]}
   );
   gpc615_5 gpc1064 (
      {stage0_53[174], stage0_53[175], stage0_53[176], stage0_53[177], stage0_53[178]},
      {stage0_54[162]},
      {stage0_55[84], stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89]},
      {stage1_57[14],stage1_56[41],stage1_55[56],stage1_54[66],stage1_53[90]}
   );
   gpc615_5 gpc1065 (
      {stage0_53[179], stage0_53[180], stage0_53[181], stage0_53[182], stage0_53[183]},
      {stage0_54[163]},
      {stage0_55[90], stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95]},
      {stage1_57[15],stage1_56[42],stage1_55[57],stage1_54[67],stage1_53[91]}
   );
   gpc615_5 gpc1066 (
      {stage0_53[184], stage0_53[185], stage0_53[186], stage0_53[187], stage0_53[188]},
      {stage0_54[164]},
      {stage0_55[96], stage0_55[97], stage0_55[98], stage0_55[99], stage0_55[100], stage0_55[101]},
      {stage1_57[16],stage1_56[43],stage1_55[58],stage1_54[68],stage1_53[92]}
   );
   gpc615_5 gpc1067 (
      {stage0_53[189], stage0_53[190], stage0_53[191], stage0_53[192], stage0_53[193]},
      {stage0_54[165]},
      {stage0_55[102], stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106], stage0_55[107]},
      {stage1_57[17],stage1_56[44],stage1_55[59],stage1_54[69],stage1_53[93]}
   );
   gpc615_5 gpc1068 (
      {stage0_53[194], stage0_53[195], stage0_53[196], stage0_53[197], stage0_53[198]},
      {stage0_54[166]},
      {stage0_55[108], stage0_55[109], stage0_55[110], stage0_55[111], stage0_55[112], stage0_55[113]},
      {stage1_57[18],stage1_56[45],stage1_55[60],stage1_54[70],stage1_53[94]}
   );
   gpc615_5 gpc1069 (
      {stage0_53[199], stage0_53[200], stage0_53[201], stage0_53[202], stage0_53[203]},
      {stage0_54[167]},
      {stage0_55[114], stage0_55[115], stage0_55[116], stage0_55[117], stage0_55[118], stage0_55[119]},
      {stage1_57[19],stage1_56[46],stage1_55[61],stage1_54[71],stage1_53[95]}
   );
   gpc615_5 gpc1070 (
      {stage0_53[204], stage0_53[205], stage0_53[206], stage0_53[207], stage0_53[208]},
      {stage0_54[168]},
      {stage0_55[120], stage0_55[121], stage0_55[122], stage0_55[123], stage0_55[124], stage0_55[125]},
      {stage1_57[20],stage1_56[47],stage1_55[62],stage1_54[72],stage1_53[96]}
   );
   gpc615_5 gpc1071 (
      {stage0_53[209], stage0_53[210], stage0_53[211], stage0_53[212], stage0_53[213]},
      {stage0_54[169]},
      {stage0_55[126], stage0_55[127], stage0_55[128], stage0_55[129], stage0_55[130], stage0_55[131]},
      {stage1_57[21],stage1_56[48],stage1_55[63],stage1_54[73],stage1_53[97]}
   );
   gpc615_5 gpc1072 (
      {stage0_53[214], stage0_53[215], stage0_53[216], stage0_53[217], stage0_53[218]},
      {stage0_54[170]},
      {stage0_55[132], stage0_55[133], stage0_55[134], stage0_55[135], stage0_55[136], stage0_55[137]},
      {stage1_57[22],stage1_56[49],stage1_55[64],stage1_54[74],stage1_53[98]}
   );
   gpc615_5 gpc1073 (
      {stage0_53[219], stage0_53[220], stage0_53[221], stage0_53[222], stage0_53[223]},
      {stage0_54[171]},
      {stage0_55[138], stage0_55[139], stage0_55[140], stage0_55[141], stage0_55[142], stage0_55[143]},
      {stage1_57[23],stage1_56[50],stage1_55[65],stage1_54[75],stage1_53[99]}
   );
   gpc615_5 gpc1074 (
      {stage0_53[224], stage0_53[225], stage0_53[226], stage0_53[227], stage0_53[228]},
      {stage0_54[172]},
      {stage0_55[144], stage0_55[145], stage0_55[146], stage0_55[147], stage0_55[148], stage0_55[149]},
      {stage1_57[24],stage1_56[51],stage1_55[66],stage1_54[76],stage1_53[100]}
   );
   gpc615_5 gpc1075 (
      {stage0_53[229], stage0_53[230], stage0_53[231], stage0_53[232], stage0_53[233]},
      {stage0_54[173]},
      {stage0_55[150], stage0_55[151], stage0_55[152], stage0_55[153], stage0_55[154], stage0_55[155]},
      {stage1_57[25],stage1_56[52],stage1_55[67],stage1_54[77],stage1_53[101]}
   );
   gpc615_5 gpc1076 (
      {stage0_53[234], stage0_53[235], stage0_53[236], stage0_53[237], stage0_53[238]},
      {stage0_54[174]},
      {stage0_55[156], stage0_55[157], stage0_55[158], stage0_55[159], stage0_55[160], stage0_55[161]},
      {stage1_57[26],stage1_56[53],stage1_55[68],stage1_54[78],stage1_53[102]}
   );
   gpc615_5 gpc1077 (
      {stage0_53[239], stage0_53[240], stage0_53[241], stage0_53[242], stage0_53[243]},
      {stage0_54[175]},
      {stage0_55[162], stage0_55[163], stage0_55[164], stage0_55[165], stage0_55[166], stage0_55[167]},
      {stage1_57[27],stage1_56[54],stage1_55[69],stage1_54[79],stage1_53[103]}
   );
   gpc615_5 gpc1078 (
      {stage0_53[244], stage0_53[245], stage0_53[246], stage0_53[247], stage0_53[248]},
      {stage0_54[176]},
      {stage0_55[168], stage0_55[169], stage0_55[170], stage0_55[171], stage0_55[172], stage0_55[173]},
      {stage1_57[28],stage1_56[55],stage1_55[70],stage1_54[80],stage1_53[104]}
   );
   gpc615_5 gpc1079 (
      {stage0_53[249], stage0_53[250], stage0_53[251], stage0_53[252], stage0_53[253]},
      {stage0_54[177]},
      {stage0_55[174], stage0_55[175], stage0_55[176], stage0_55[177], stage0_55[178], stage0_55[179]},
      {stage1_57[29],stage1_56[56],stage1_55[71],stage1_54[81],stage1_53[105]}
   );
   gpc606_5 gpc1080 (
      {stage0_55[180], stage0_55[181], stage0_55[182], stage0_55[183], stage0_55[184], stage0_55[185]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[0],stage1_57[30],stage1_56[57],stage1_55[72]}
   );
   gpc606_5 gpc1081 (
      {stage0_55[186], stage0_55[187], stage0_55[188], stage0_55[189], stage0_55[190], stage0_55[191]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[1],stage1_57[31],stage1_56[58],stage1_55[73]}
   );
   gpc606_5 gpc1082 (
      {stage0_55[192], stage0_55[193], stage0_55[194], stage0_55[195], stage0_55[196], stage0_55[197]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[2],stage1_57[32],stage1_56[59],stage1_55[74]}
   );
   gpc606_5 gpc1083 (
      {stage0_55[198], stage0_55[199], stage0_55[200], stage0_55[201], stage0_55[202], stage0_55[203]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[3],stage1_57[33],stage1_56[60],stage1_55[75]}
   );
   gpc606_5 gpc1084 (
      {stage0_55[204], stage0_55[205], stage0_55[206], stage0_55[207], stage0_55[208], stage0_55[209]},
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage1_59[4],stage1_58[4],stage1_57[34],stage1_56[61],stage1_55[76]}
   );
   gpc606_5 gpc1085 (
      {stage0_55[210], stage0_55[211], stage0_55[212], stage0_55[213], stage0_55[214], stage0_55[215]},
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage1_59[5],stage1_58[5],stage1_57[35],stage1_56[62],stage1_55[77]}
   );
   gpc606_5 gpc1086 (
      {stage0_55[216], stage0_55[217], stage0_55[218], stage0_55[219], stage0_55[220], stage0_55[221]},
      {stage0_57[36], stage0_57[37], stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41]},
      {stage1_59[6],stage1_58[6],stage1_57[36],stage1_56[63],stage1_55[78]}
   );
   gpc606_5 gpc1087 (
      {stage0_55[222], stage0_55[223], stage0_55[224], stage0_55[225], stage0_55[226], stage0_55[227]},
      {stage0_57[42], stage0_57[43], stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47]},
      {stage1_59[7],stage1_58[7],stage1_57[37],stage1_56[64],stage1_55[79]}
   );
   gpc606_5 gpc1088 (
      {stage0_55[228], stage0_55[229], stage0_55[230], stage0_55[231], stage0_55[232], stage0_55[233]},
      {stage0_57[48], stage0_57[49], stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53]},
      {stage1_59[8],stage1_58[8],stage1_57[38],stage1_56[65],stage1_55[80]}
   );
   gpc606_5 gpc1089 (
      {stage0_55[234], stage0_55[235], stage0_55[236], stage0_55[237], stage0_55[238], stage0_55[239]},
      {stage0_57[54], stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage1_59[9],stage1_58[9],stage1_57[39],stage1_56[66],stage1_55[81]}
   );
   gpc615_5 gpc1090 (
      {stage0_55[240], stage0_55[241], stage0_55[242], stage0_55[243], stage0_55[244]},
      {stage0_56[0]},
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65]},
      {stage1_59[10],stage1_58[10],stage1_57[40],stage1_56[67],stage1_55[82]}
   );
   gpc615_5 gpc1091 (
      {stage0_55[245], stage0_55[246], stage0_55[247], stage0_55[248], stage0_55[249]},
      {stage0_56[1]},
      {stage0_57[66], stage0_57[67], stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71]},
      {stage1_59[11],stage1_58[11],stage1_57[41],stage1_56[68],stage1_55[83]}
   );
   gpc606_5 gpc1092 (
      {stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5], stage0_56[6], stage0_56[7]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[12],stage1_58[12],stage1_57[42],stage1_56[69]}
   );
   gpc606_5 gpc1093 (
      {stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11], stage0_56[12], stage0_56[13]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[13],stage1_58[13],stage1_57[43],stage1_56[70]}
   );
   gpc606_5 gpc1094 (
      {stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17], stage0_56[18], stage0_56[19]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[14],stage1_58[14],stage1_57[44],stage1_56[71]}
   );
   gpc606_5 gpc1095 (
      {stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23], stage0_56[24], stage0_56[25]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[15],stage1_58[15],stage1_57[45],stage1_56[72]}
   );
   gpc606_5 gpc1096 (
      {stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29], stage0_56[30], stage0_56[31]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[16],stage1_58[16],stage1_57[46],stage1_56[73]}
   );
   gpc606_5 gpc1097 (
      {stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35], stage0_56[36], stage0_56[37]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[17],stage1_58[17],stage1_57[47],stage1_56[74]}
   );
   gpc606_5 gpc1098 (
      {stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41], stage0_56[42], stage0_56[43]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[18],stage1_58[18],stage1_57[48],stage1_56[75]}
   );
   gpc606_5 gpc1099 (
      {stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47], stage0_56[48], stage0_56[49]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[19],stage1_58[19],stage1_57[49],stage1_56[76]}
   );
   gpc606_5 gpc1100 (
      {stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53], stage0_56[54], stage0_56[55]},
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage1_60[8],stage1_59[20],stage1_58[20],stage1_57[50],stage1_56[77]}
   );
   gpc606_5 gpc1101 (
      {stage0_56[56], stage0_56[57], stage0_56[58], stage0_56[59], stage0_56[60], stage0_56[61]},
      {stage0_58[54], stage0_58[55], stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59]},
      {stage1_60[9],stage1_59[21],stage1_58[21],stage1_57[51],stage1_56[78]}
   );
   gpc606_5 gpc1102 (
      {stage0_56[62], stage0_56[63], stage0_56[64], stage0_56[65], stage0_56[66], stage0_56[67]},
      {stage0_58[60], stage0_58[61], stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65]},
      {stage1_60[10],stage1_59[22],stage1_58[22],stage1_57[52],stage1_56[79]}
   );
   gpc606_5 gpc1103 (
      {stage0_56[68], stage0_56[69], stage0_56[70], stage0_56[71], stage0_56[72], stage0_56[73]},
      {stage0_58[66], stage0_58[67], stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71]},
      {stage1_60[11],stage1_59[23],stage1_58[23],stage1_57[53],stage1_56[80]}
   );
   gpc606_5 gpc1104 (
      {stage0_56[74], stage0_56[75], stage0_56[76], stage0_56[77], stage0_56[78], stage0_56[79]},
      {stage0_58[72], stage0_58[73], stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77]},
      {stage1_60[12],stage1_59[24],stage1_58[24],stage1_57[54],stage1_56[81]}
   );
   gpc606_5 gpc1105 (
      {stage0_56[80], stage0_56[81], stage0_56[82], stage0_56[83], stage0_56[84], stage0_56[85]},
      {stage0_58[78], stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage1_60[13],stage1_59[25],stage1_58[25],stage1_57[55],stage1_56[82]}
   );
   gpc606_5 gpc1106 (
      {stage0_56[86], stage0_56[87], stage0_56[88], stage0_56[89], stage0_56[90], stage0_56[91]},
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88], stage0_58[89]},
      {stage1_60[14],stage1_59[26],stage1_58[26],stage1_57[56],stage1_56[83]}
   );
   gpc606_5 gpc1107 (
      {stage0_56[92], stage0_56[93], stage0_56[94], stage0_56[95], stage0_56[96], stage0_56[97]},
      {stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93], stage0_58[94], stage0_58[95]},
      {stage1_60[15],stage1_59[27],stage1_58[27],stage1_57[57],stage1_56[84]}
   );
   gpc606_5 gpc1108 (
      {stage0_56[98], stage0_56[99], stage0_56[100], stage0_56[101], stage0_56[102], stage0_56[103]},
      {stage0_58[96], stage0_58[97], stage0_58[98], stage0_58[99], stage0_58[100], stage0_58[101]},
      {stage1_60[16],stage1_59[28],stage1_58[28],stage1_57[58],stage1_56[85]}
   );
   gpc606_5 gpc1109 (
      {stage0_56[104], stage0_56[105], stage0_56[106], stage0_56[107], stage0_56[108], stage0_56[109]},
      {stage0_58[102], stage0_58[103], stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107]},
      {stage1_60[17],stage1_59[29],stage1_58[29],stage1_57[59],stage1_56[86]}
   );
   gpc606_5 gpc1110 (
      {stage0_56[110], stage0_56[111], stage0_56[112], stage0_56[113], stage0_56[114], stage0_56[115]},
      {stage0_58[108], stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage1_60[18],stage1_59[30],stage1_58[30],stage1_57[60],stage1_56[87]}
   );
   gpc606_5 gpc1111 (
      {stage0_56[116], stage0_56[117], stage0_56[118], stage0_56[119], stage0_56[120], stage0_56[121]},
      {stage0_58[114], stage0_58[115], stage0_58[116], stage0_58[117], stage0_58[118], stage0_58[119]},
      {stage1_60[19],stage1_59[31],stage1_58[31],stage1_57[61],stage1_56[88]}
   );
   gpc606_5 gpc1112 (
      {stage0_56[122], stage0_56[123], stage0_56[124], stage0_56[125], stage0_56[126], stage0_56[127]},
      {stage0_58[120], stage0_58[121], stage0_58[122], stage0_58[123], stage0_58[124], stage0_58[125]},
      {stage1_60[20],stage1_59[32],stage1_58[32],stage1_57[62],stage1_56[89]}
   );
   gpc606_5 gpc1113 (
      {stage0_56[128], stage0_56[129], stage0_56[130], stage0_56[131], stage0_56[132], stage0_56[133]},
      {stage0_58[126], stage0_58[127], stage0_58[128], stage0_58[129], stage0_58[130], stage0_58[131]},
      {stage1_60[21],stage1_59[33],stage1_58[33],stage1_57[63],stage1_56[90]}
   );
   gpc606_5 gpc1114 (
      {stage0_56[134], stage0_56[135], stage0_56[136], stage0_56[137], stage0_56[138], stage0_56[139]},
      {stage0_58[132], stage0_58[133], stage0_58[134], stage0_58[135], stage0_58[136], stage0_58[137]},
      {stage1_60[22],stage1_59[34],stage1_58[34],stage1_57[64],stage1_56[91]}
   );
   gpc606_5 gpc1115 (
      {stage0_56[140], stage0_56[141], stage0_56[142], stage0_56[143], stage0_56[144], stage0_56[145]},
      {stage0_58[138], stage0_58[139], stage0_58[140], stage0_58[141], stage0_58[142], stage0_58[143]},
      {stage1_60[23],stage1_59[35],stage1_58[35],stage1_57[65],stage1_56[92]}
   );
   gpc606_5 gpc1116 (
      {stage0_56[146], stage0_56[147], stage0_56[148], stage0_56[149], stage0_56[150], stage0_56[151]},
      {stage0_58[144], stage0_58[145], stage0_58[146], stage0_58[147], stage0_58[148], stage0_58[149]},
      {stage1_60[24],stage1_59[36],stage1_58[36],stage1_57[66],stage1_56[93]}
   );
   gpc606_5 gpc1117 (
      {stage0_56[152], stage0_56[153], stage0_56[154], stage0_56[155], stage0_56[156], stage0_56[157]},
      {stage0_58[150], stage0_58[151], stage0_58[152], stage0_58[153], stage0_58[154], stage0_58[155]},
      {stage1_60[25],stage1_59[37],stage1_58[37],stage1_57[67],stage1_56[94]}
   );
   gpc606_5 gpc1118 (
      {stage0_56[158], stage0_56[159], stage0_56[160], stage0_56[161], stage0_56[162], stage0_56[163]},
      {stage0_58[156], stage0_58[157], stage0_58[158], stage0_58[159], stage0_58[160], stage0_58[161]},
      {stage1_60[26],stage1_59[38],stage1_58[38],stage1_57[68],stage1_56[95]}
   );
   gpc606_5 gpc1119 (
      {stage0_56[164], stage0_56[165], stage0_56[166], stage0_56[167], stage0_56[168], stage0_56[169]},
      {stage0_58[162], stage0_58[163], stage0_58[164], stage0_58[165], stage0_58[166], stage0_58[167]},
      {stage1_60[27],stage1_59[39],stage1_58[39],stage1_57[69],stage1_56[96]}
   );
   gpc606_5 gpc1120 (
      {stage0_56[170], stage0_56[171], stage0_56[172], stage0_56[173], stage0_56[174], stage0_56[175]},
      {stage0_58[168], stage0_58[169], stage0_58[170], stage0_58[171], stage0_58[172], stage0_58[173]},
      {stage1_60[28],stage1_59[40],stage1_58[40],stage1_57[70],stage1_56[97]}
   );
   gpc606_5 gpc1121 (
      {stage0_57[72], stage0_57[73], stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[29],stage1_59[41],stage1_58[41],stage1_57[71]}
   );
   gpc606_5 gpc1122 (
      {stage0_57[78], stage0_57[79], stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[30],stage1_59[42],stage1_58[42],stage1_57[72]}
   );
   gpc606_5 gpc1123 (
      {stage0_57[84], stage0_57[85], stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[31],stage1_59[43],stage1_58[43],stage1_57[73]}
   );
   gpc606_5 gpc1124 (
      {stage0_57[90], stage0_57[91], stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[32],stage1_59[44],stage1_58[44],stage1_57[74]}
   );
   gpc606_5 gpc1125 (
      {stage0_57[96], stage0_57[97], stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[33],stage1_59[45],stage1_58[45],stage1_57[75]}
   );
   gpc606_5 gpc1126 (
      {stage0_57[102], stage0_57[103], stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[34],stage1_59[46],stage1_58[46],stage1_57[76]}
   );
   gpc606_5 gpc1127 (
      {stage0_57[108], stage0_57[109], stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[35],stage1_59[47],stage1_58[47],stage1_57[77]}
   );
   gpc606_5 gpc1128 (
      {stage0_57[114], stage0_57[115], stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[36],stage1_59[48],stage1_58[48],stage1_57[78]}
   );
   gpc606_5 gpc1129 (
      {stage0_57[120], stage0_57[121], stage0_57[122], stage0_57[123], stage0_57[124], stage0_57[125]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[37],stage1_59[49],stage1_58[49],stage1_57[79]}
   );
   gpc606_5 gpc1130 (
      {stage0_57[126], stage0_57[127], stage0_57[128], stage0_57[129], stage0_57[130], stage0_57[131]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[38],stage1_59[50],stage1_58[50],stage1_57[80]}
   );
   gpc606_5 gpc1131 (
      {stage0_57[132], stage0_57[133], stage0_57[134], stage0_57[135], stage0_57[136], stage0_57[137]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[39],stage1_59[51],stage1_58[51],stage1_57[81]}
   );
   gpc606_5 gpc1132 (
      {stage0_57[138], stage0_57[139], stage0_57[140], stage0_57[141], stage0_57[142], stage0_57[143]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[40],stage1_59[52],stage1_58[52],stage1_57[82]}
   );
   gpc606_5 gpc1133 (
      {stage0_57[144], stage0_57[145], stage0_57[146], stage0_57[147], stage0_57[148], stage0_57[149]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[41],stage1_59[53],stage1_58[53],stage1_57[83]}
   );
   gpc606_5 gpc1134 (
      {stage0_57[150], stage0_57[151], stage0_57[152], stage0_57[153], stage0_57[154], stage0_57[155]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[42],stage1_59[54],stage1_58[54],stage1_57[84]}
   );
   gpc606_5 gpc1135 (
      {stage0_57[156], stage0_57[157], stage0_57[158], stage0_57[159], stage0_57[160], stage0_57[161]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[43],stage1_59[55],stage1_58[55],stage1_57[85]}
   );
   gpc606_5 gpc1136 (
      {stage0_57[162], stage0_57[163], stage0_57[164], stage0_57[165], stage0_57[166], stage0_57[167]},
      {stage0_59[90], stage0_59[91], stage0_59[92], stage0_59[93], stage0_59[94], stage0_59[95]},
      {stage1_61[15],stage1_60[44],stage1_59[56],stage1_58[56],stage1_57[86]}
   );
   gpc606_5 gpc1137 (
      {stage0_57[168], stage0_57[169], stage0_57[170], stage0_57[171], stage0_57[172], stage0_57[173]},
      {stage0_59[96], stage0_59[97], stage0_59[98], stage0_59[99], stage0_59[100], stage0_59[101]},
      {stage1_61[16],stage1_60[45],stage1_59[57],stage1_58[57],stage1_57[87]}
   );
   gpc606_5 gpc1138 (
      {stage0_57[174], stage0_57[175], stage0_57[176], stage0_57[177], stage0_57[178], stage0_57[179]},
      {stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105], stage0_59[106], stage0_59[107]},
      {stage1_61[17],stage1_60[46],stage1_59[58],stage1_58[58],stage1_57[88]}
   );
   gpc606_5 gpc1139 (
      {stage0_57[180], stage0_57[181], stage0_57[182], stage0_57[183], stage0_57[184], stage0_57[185]},
      {stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111], stage0_59[112], stage0_59[113]},
      {stage1_61[18],stage1_60[47],stage1_59[59],stage1_58[59],stage1_57[89]}
   );
   gpc606_5 gpc1140 (
      {stage0_57[186], stage0_57[187], stage0_57[188], stage0_57[189], stage0_57[190], stage0_57[191]},
      {stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117], stage0_59[118], stage0_59[119]},
      {stage1_61[19],stage1_60[48],stage1_59[60],stage1_58[60],stage1_57[90]}
   );
   gpc606_5 gpc1141 (
      {stage0_57[192], stage0_57[193], stage0_57[194], stage0_57[195], stage0_57[196], stage0_57[197]},
      {stage0_59[120], stage0_59[121], stage0_59[122], stage0_59[123], stage0_59[124], stage0_59[125]},
      {stage1_61[20],stage1_60[49],stage1_59[61],stage1_58[61],stage1_57[91]}
   );
   gpc606_5 gpc1142 (
      {stage0_57[198], stage0_57[199], stage0_57[200], stage0_57[201], stage0_57[202], stage0_57[203]},
      {stage0_59[126], stage0_59[127], stage0_59[128], stage0_59[129], stage0_59[130], stage0_59[131]},
      {stage1_61[21],stage1_60[50],stage1_59[62],stage1_58[62],stage1_57[92]}
   );
   gpc606_5 gpc1143 (
      {stage0_57[204], stage0_57[205], stage0_57[206], stage0_57[207], stage0_57[208], stage0_57[209]},
      {stage0_59[132], stage0_59[133], stage0_59[134], stage0_59[135], stage0_59[136], stage0_59[137]},
      {stage1_61[22],stage1_60[51],stage1_59[63],stage1_58[63],stage1_57[93]}
   );
   gpc606_5 gpc1144 (
      {stage0_57[210], stage0_57[211], stage0_57[212], stage0_57[213], stage0_57[214], stage0_57[215]},
      {stage0_59[138], stage0_59[139], stage0_59[140], stage0_59[141], stage0_59[142], stage0_59[143]},
      {stage1_61[23],stage1_60[52],stage1_59[64],stage1_58[64],stage1_57[94]}
   );
   gpc606_5 gpc1145 (
      {stage0_57[216], stage0_57[217], stage0_57[218], stage0_57[219], stage0_57[220], stage0_57[221]},
      {stage0_59[144], stage0_59[145], stage0_59[146], stage0_59[147], stage0_59[148], stage0_59[149]},
      {stage1_61[24],stage1_60[53],stage1_59[65],stage1_58[65],stage1_57[95]}
   );
   gpc606_5 gpc1146 (
      {stage0_57[222], stage0_57[223], stage0_57[224], stage0_57[225], stage0_57[226], stage0_57[227]},
      {stage0_59[150], stage0_59[151], stage0_59[152], stage0_59[153], stage0_59[154], stage0_59[155]},
      {stage1_61[25],stage1_60[54],stage1_59[66],stage1_58[66],stage1_57[96]}
   );
   gpc615_5 gpc1147 (
      {stage0_57[228], stage0_57[229], stage0_57[230], stage0_57[231], stage0_57[232]},
      {stage0_58[174]},
      {stage0_59[156], stage0_59[157], stage0_59[158], stage0_59[159], stage0_59[160], stage0_59[161]},
      {stage1_61[26],stage1_60[55],stage1_59[67],stage1_58[67],stage1_57[97]}
   );
   gpc615_5 gpc1148 (
      {stage0_57[233], stage0_57[234], stage0_57[235], stage0_57[236], stage0_57[237]},
      {stage0_58[175]},
      {stage0_59[162], stage0_59[163], stage0_59[164], stage0_59[165], stage0_59[166], stage0_59[167]},
      {stage1_61[27],stage1_60[56],stage1_59[68],stage1_58[68],stage1_57[98]}
   );
   gpc615_5 gpc1149 (
      {stage0_57[238], stage0_57[239], stage0_57[240], stage0_57[241], stage0_57[242]},
      {stage0_58[176]},
      {stage0_59[168], stage0_59[169], stage0_59[170], stage0_59[171], stage0_59[172], stage0_59[173]},
      {stage1_61[28],stage1_60[57],stage1_59[69],stage1_58[69],stage1_57[99]}
   );
   gpc615_5 gpc1150 (
      {stage0_57[243], stage0_57[244], stage0_57[245], stage0_57[246], stage0_57[247]},
      {stage0_58[177]},
      {stage0_59[174], stage0_59[175], stage0_59[176], stage0_59[177], stage0_59[178], stage0_59[179]},
      {stage1_61[29],stage1_60[58],stage1_59[70],stage1_58[70],stage1_57[100]}
   );
   gpc615_5 gpc1151 (
      {stage0_57[248], stage0_57[249], stage0_57[250], stage0_57[251], stage0_57[252]},
      {stage0_58[178]},
      {stage0_59[180], stage0_59[181], stage0_59[182], stage0_59[183], stage0_59[184], stage0_59[185]},
      {stage1_61[30],stage1_60[59],stage1_59[71],stage1_58[71],stage1_57[101]}
   );
   gpc606_5 gpc1152 (
      {stage0_58[179], stage0_58[180], stage0_58[181], stage0_58[182], stage0_58[183], stage0_58[184]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[31],stage1_60[60],stage1_59[72],stage1_58[72]}
   );
   gpc606_5 gpc1153 (
      {stage0_58[185], stage0_58[186], stage0_58[187], stage0_58[188], stage0_58[189], stage0_58[190]},
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage1_62[1],stage1_61[32],stage1_60[61],stage1_59[73],stage1_58[73]}
   );
   gpc606_5 gpc1154 (
      {stage0_58[191], stage0_58[192], stage0_58[193], stage0_58[194], stage0_58[195], stage0_58[196]},
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage1_62[2],stage1_61[33],stage1_60[62],stage1_59[74],stage1_58[74]}
   );
   gpc606_5 gpc1155 (
      {stage0_58[197], stage0_58[198], stage0_58[199], stage0_58[200], stage0_58[201], stage0_58[202]},
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage1_62[3],stage1_61[34],stage1_60[63],stage1_59[75],stage1_58[75]}
   );
   gpc606_5 gpc1156 (
      {stage0_58[203], stage0_58[204], stage0_58[205], stage0_58[206], stage0_58[207], stage0_58[208]},
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage1_62[4],stage1_61[35],stage1_60[64],stage1_59[76],stage1_58[76]}
   );
   gpc606_5 gpc1157 (
      {stage0_58[209], stage0_58[210], stage0_58[211], stage0_58[212], stage0_58[213], stage0_58[214]},
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage1_62[5],stage1_61[36],stage1_60[65],stage1_59[77],stage1_58[77]}
   );
   gpc606_5 gpc1158 (
      {stage0_58[215], stage0_58[216], stage0_58[217], stage0_58[218], stage0_58[219], stage0_58[220]},
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage1_62[6],stage1_61[37],stage1_60[66],stage1_59[78],stage1_58[78]}
   );
   gpc606_5 gpc1159 (
      {stage0_58[221], stage0_58[222], stage0_58[223], stage0_58[224], stage0_58[225], stage0_58[226]},
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage1_62[7],stage1_61[38],stage1_60[67],stage1_59[79],stage1_58[79]}
   );
   gpc606_5 gpc1160 (
      {stage0_58[227], stage0_58[228], stage0_58[229], stage0_58[230], stage0_58[231], stage0_58[232]},
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage1_62[8],stage1_61[39],stage1_60[68],stage1_59[80],stage1_58[80]}
   );
   gpc606_5 gpc1161 (
      {stage0_58[233], stage0_58[234], stage0_58[235], stage0_58[236], stage0_58[237], stage0_58[238]},
      {stage0_60[54], stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59]},
      {stage1_62[9],stage1_61[40],stage1_60[69],stage1_59[81],stage1_58[81]}
   );
   gpc606_5 gpc1162 (
      {stage0_58[239], stage0_58[240], stage0_58[241], stage0_58[242], stage0_58[243], stage0_58[244]},
      {stage0_60[60], stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65]},
      {stage1_62[10],stage1_61[41],stage1_60[70],stage1_59[82],stage1_58[82]}
   );
   gpc615_5 gpc1163 (
      {stage0_58[245], stage0_58[246], stage0_58[247], stage0_58[248], stage0_58[249]},
      {stage0_59[186]},
      {stage0_60[66], stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71]},
      {stage1_62[11],stage1_61[42],stage1_60[71],stage1_59[83],stage1_58[83]}
   );
   gpc615_5 gpc1164 (
      {stage0_58[250], stage0_58[251], stage0_58[252], stage0_58[253], stage0_58[254]},
      {stage0_59[187]},
      {stage0_60[72], stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77]},
      {stage1_62[12],stage1_61[43],stage1_60[72],stage1_59[84],stage1_58[84]}
   );
   gpc1406_5 gpc1165 (
      {stage0_59[188], stage0_59[189], stage0_59[190], stage0_59[191], stage0_59[192], stage0_59[193]},
      {stage0_61[0], stage0_61[1], stage0_61[2], stage0_61[3]},
      {stage0_62[0]},
      {stage1_63[0],stage1_62[13],stage1_61[44],stage1_60[73],stage1_59[85]}
   );
   gpc606_5 gpc1166 (
      {stage0_60[78], stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83]},
      {stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5], stage0_62[6]},
      {stage1_64[0],stage1_63[1],stage1_62[14],stage1_61[45],stage1_60[74]}
   );
   gpc606_5 gpc1167 (
      {stage0_60[84], stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89]},
      {stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11], stage0_62[12]},
      {stage1_64[1],stage1_63[2],stage1_62[15],stage1_61[46],stage1_60[75]}
   );
   gpc606_5 gpc1168 (
      {stage0_60[90], stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95]},
      {stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17], stage0_62[18]},
      {stage1_64[2],stage1_63[3],stage1_62[16],stage1_61[47],stage1_60[76]}
   );
   gpc606_5 gpc1169 (
      {stage0_60[96], stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101]},
      {stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23], stage0_62[24]},
      {stage1_64[3],stage1_63[4],stage1_62[17],stage1_61[48],stage1_60[77]}
   );
   gpc606_5 gpc1170 (
      {stage0_60[102], stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107]},
      {stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29], stage0_62[30]},
      {stage1_64[4],stage1_63[5],stage1_62[18],stage1_61[49],stage1_60[78]}
   );
   gpc606_5 gpc1171 (
      {stage0_60[108], stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113]},
      {stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35], stage0_62[36]},
      {stage1_64[5],stage1_63[6],stage1_62[19],stage1_61[50],stage1_60[79]}
   );
   gpc606_5 gpc1172 (
      {stage0_60[114], stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119]},
      {stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41], stage0_62[42]},
      {stage1_64[6],stage1_63[7],stage1_62[20],stage1_61[51],stage1_60[80]}
   );
   gpc606_5 gpc1173 (
      {stage0_60[120], stage0_60[121], stage0_60[122], stage0_60[123], stage0_60[124], stage0_60[125]},
      {stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47], stage0_62[48]},
      {stage1_64[7],stage1_63[8],stage1_62[21],stage1_61[52],stage1_60[81]}
   );
   gpc606_5 gpc1174 (
      {stage0_60[126], stage0_60[127], stage0_60[128], stage0_60[129], stage0_60[130], stage0_60[131]},
      {stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53], stage0_62[54]},
      {stage1_64[8],stage1_63[9],stage1_62[22],stage1_61[53],stage1_60[82]}
   );
   gpc606_5 gpc1175 (
      {stage0_60[132], stage0_60[133], stage0_60[134], stage0_60[135], stage0_60[136], stage0_60[137]},
      {stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59], stage0_62[60]},
      {stage1_64[9],stage1_63[10],stage1_62[23],stage1_61[54],stage1_60[83]}
   );
   gpc606_5 gpc1176 (
      {stage0_60[138], stage0_60[139], stage0_60[140], stage0_60[141], stage0_60[142], stage0_60[143]},
      {stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65], stage0_62[66]},
      {stage1_64[10],stage1_63[11],stage1_62[24],stage1_61[55],stage1_60[84]}
   );
   gpc606_5 gpc1177 (
      {stage0_60[144], stage0_60[145], stage0_60[146], stage0_60[147], stage0_60[148], stage0_60[149]},
      {stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71], stage0_62[72]},
      {stage1_64[11],stage1_63[12],stage1_62[25],stage1_61[56],stage1_60[85]}
   );
   gpc606_5 gpc1178 (
      {stage0_60[150], stage0_60[151], stage0_60[152], stage0_60[153], stage0_60[154], stage0_60[155]},
      {stage0_62[73], stage0_62[74], stage0_62[75], stage0_62[76], stage0_62[77], stage0_62[78]},
      {stage1_64[12],stage1_63[13],stage1_62[26],stage1_61[57],stage1_60[86]}
   );
   gpc606_5 gpc1179 (
      {stage0_60[156], stage0_60[157], stage0_60[158], stage0_60[159], stage0_60[160], stage0_60[161]},
      {stage0_62[79], stage0_62[80], stage0_62[81], stage0_62[82], stage0_62[83], stage0_62[84]},
      {stage1_64[13],stage1_63[14],stage1_62[27],stage1_61[58],stage1_60[87]}
   );
   gpc606_5 gpc1180 (
      {stage0_60[162], stage0_60[163], stage0_60[164], stage0_60[165], stage0_60[166], stage0_60[167]},
      {stage0_62[85], stage0_62[86], stage0_62[87], stage0_62[88], stage0_62[89], stage0_62[90]},
      {stage1_64[14],stage1_63[15],stage1_62[28],stage1_61[59],stage1_60[88]}
   );
   gpc606_5 gpc1181 (
      {stage0_60[168], stage0_60[169], stage0_60[170], stage0_60[171], stage0_60[172], stage0_60[173]},
      {stage0_62[91], stage0_62[92], stage0_62[93], stage0_62[94], stage0_62[95], stage0_62[96]},
      {stage1_64[15],stage1_63[16],stage1_62[29],stage1_61[60],stage1_60[89]}
   );
   gpc606_5 gpc1182 (
      {stage0_60[174], stage0_60[175], stage0_60[176], stage0_60[177], stage0_60[178], stage0_60[179]},
      {stage0_62[97], stage0_62[98], stage0_62[99], stage0_62[100], stage0_62[101], stage0_62[102]},
      {stage1_64[16],stage1_63[17],stage1_62[30],stage1_61[61],stage1_60[90]}
   );
   gpc606_5 gpc1183 (
      {stage0_60[180], stage0_60[181], stage0_60[182], stage0_60[183], stage0_60[184], stage0_60[185]},
      {stage0_62[103], stage0_62[104], stage0_62[105], stage0_62[106], stage0_62[107], stage0_62[108]},
      {stage1_64[17],stage1_63[18],stage1_62[31],stage1_61[62],stage1_60[91]}
   );
   gpc606_5 gpc1184 (
      {stage0_60[186], stage0_60[187], stage0_60[188], stage0_60[189], stage0_60[190], stage0_60[191]},
      {stage0_62[109], stage0_62[110], stage0_62[111], stage0_62[112], stage0_62[113], stage0_62[114]},
      {stage1_64[18],stage1_63[19],stage1_62[32],stage1_61[63],stage1_60[92]}
   );
   gpc606_5 gpc1185 (
      {stage0_60[192], stage0_60[193], stage0_60[194], stage0_60[195], stage0_60[196], stage0_60[197]},
      {stage0_62[115], stage0_62[116], stage0_62[117], stage0_62[118], stage0_62[119], stage0_62[120]},
      {stage1_64[19],stage1_63[20],stage1_62[33],stage1_61[64],stage1_60[93]}
   );
   gpc606_5 gpc1186 (
      {stage0_60[198], stage0_60[199], stage0_60[200], stage0_60[201], stage0_60[202], stage0_60[203]},
      {stage0_62[121], stage0_62[122], stage0_62[123], stage0_62[124], stage0_62[125], stage0_62[126]},
      {stage1_64[20],stage1_63[21],stage1_62[34],stage1_61[65],stage1_60[94]}
   );
   gpc606_5 gpc1187 (
      {stage0_60[204], stage0_60[205], stage0_60[206], stage0_60[207], stage0_60[208], stage0_60[209]},
      {stage0_62[127], stage0_62[128], stage0_62[129], stage0_62[130], stage0_62[131], stage0_62[132]},
      {stage1_64[21],stage1_63[22],stage1_62[35],stage1_61[66],stage1_60[95]}
   );
   gpc606_5 gpc1188 (
      {stage0_61[4], stage0_61[5], stage0_61[6], stage0_61[7], stage0_61[8], stage0_61[9]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[22],stage1_63[23],stage1_62[36],stage1_61[67]}
   );
   gpc606_5 gpc1189 (
      {stage0_61[10], stage0_61[11], stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[23],stage1_63[24],stage1_62[37],stage1_61[68]}
   );
   gpc606_5 gpc1190 (
      {stage0_61[16], stage0_61[17], stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[24],stage1_63[25],stage1_62[38],stage1_61[69]}
   );
   gpc606_5 gpc1191 (
      {stage0_61[22], stage0_61[23], stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[25],stage1_63[26],stage1_62[39],stage1_61[70]}
   );
   gpc606_5 gpc1192 (
      {stage0_61[28], stage0_61[29], stage0_61[30], stage0_61[31], stage0_61[32], stage0_61[33]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[26],stage1_63[27],stage1_62[40],stage1_61[71]}
   );
   gpc606_5 gpc1193 (
      {stage0_61[34], stage0_61[35], stage0_61[36], stage0_61[37], stage0_61[38], stage0_61[39]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[27],stage1_63[28],stage1_62[41],stage1_61[72]}
   );
   gpc606_5 gpc1194 (
      {stage0_61[40], stage0_61[41], stage0_61[42], stage0_61[43], stage0_61[44], stage0_61[45]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[28],stage1_63[29],stage1_62[42],stage1_61[73]}
   );
   gpc606_5 gpc1195 (
      {stage0_61[46], stage0_61[47], stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[29],stage1_63[30],stage1_62[43],stage1_61[74]}
   );
   gpc606_5 gpc1196 (
      {stage0_61[52], stage0_61[53], stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[30],stage1_63[31],stage1_62[44],stage1_61[75]}
   );
   gpc606_5 gpc1197 (
      {stage0_61[58], stage0_61[59], stage0_61[60], stage0_61[61], stage0_61[62], stage0_61[63]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[31],stage1_63[32],stage1_62[45],stage1_61[76]}
   );
   gpc606_5 gpc1198 (
      {stage0_61[64], stage0_61[65], stage0_61[66], stage0_61[67], stage0_61[68], stage0_61[69]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[32],stage1_63[33],stage1_62[46],stage1_61[77]}
   );
   gpc606_5 gpc1199 (
      {stage0_61[70], stage0_61[71], stage0_61[72], stage0_61[73], stage0_61[74], stage0_61[75]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[33],stage1_63[34],stage1_62[47],stage1_61[78]}
   );
   gpc606_5 gpc1200 (
      {stage0_61[76], stage0_61[77], stage0_61[78], stage0_61[79], stage0_61[80], stage0_61[81]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[34],stage1_63[35],stage1_62[48],stage1_61[79]}
   );
   gpc606_5 gpc1201 (
      {stage0_61[82], stage0_61[83], stage0_61[84], stage0_61[85], stage0_61[86], stage0_61[87]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[35],stage1_63[36],stage1_62[49],stage1_61[80]}
   );
   gpc606_5 gpc1202 (
      {stage0_61[88], stage0_61[89], stage0_61[90], stage0_61[91], stage0_61[92], stage0_61[93]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[36],stage1_63[37],stage1_62[50],stage1_61[81]}
   );
   gpc606_5 gpc1203 (
      {stage0_61[94], stage0_61[95], stage0_61[96], stage0_61[97], stage0_61[98], stage0_61[99]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[37],stage1_63[38],stage1_62[51],stage1_61[82]}
   );
   gpc606_5 gpc1204 (
      {stage0_61[100], stage0_61[101], stage0_61[102], stage0_61[103], stage0_61[104], stage0_61[105]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[38],stage1_63[39],stage1_62[52],stage1_61[83]}
   );
   gpc606_5 gpc1205 (
      {stage0_61[106], stage0_61[107], stage0_61[108], stage0_61[109], stage0_61[110], stage0_61[111]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[39],stage1_63[40],stage1_62[53],stage1_61[84]}
   );
   gpc606_5 gpc1206 (
      {stage0_61[112], stage0_61[113], stage0_61[114], stage0_61[115], stage0_61[116], stage0_61[117]},
      {stage0_63[108], stage0_63[109], stage0_63[110], stage0_63[111], stage0_63[112], stage0_63[113]},
      {stage1_65[18],stage1_64[40],stage1_63[41],stage1_62[54],stage1_61[85]}
   );
   gpc606_5 gpc1207 (
      {stage0_61[118], stage0_61[119], stage0_61[120], stage0_61[121], stage0_61[122], stage0_61[123]},
      {stage0_63[114], stage0_63[115], stage0_63[116], stage0_63[117], stage0_63[118], stage0_63[119]},
      {stage1_65[19],stage1_64[41],stage1_63[42],stage1_62[55],stage1_61[86]}
   );
   gpc606_5 gpc1208 (
      {stage0_61[124], stage0_61[125], stage0_61[126], stage0_61[127], stage0_61[128], stage0_61[129]},
      {stage0_63[120], stage0_63[121], stage0_63[122], stage0_63[123], stage0_63[124], stage0_63[125]},
      {stage1_65[20],stage1_64[42],stage1_63[43],stage1_62[56],stage1_61[87]}
   );
   gpc606_5 gpc1209 (
      {stage0_61[130], stage0_61[131], stage0_61[132], stage0_61[133], stage0_61[134], stage0_61[135]},
      {stage0_63[126], stage0_63[127], stage0_63[128], stage0_63[129], stage0_63[130], stage0_63[131]},
      {stage1_65[21],stage1_64[43],stage1_63[44],stage1_62[57],stage1_61[88]}
   );
   gpc606_5 gpc1210 (
      {stage0_61[136], stage0_61[137], stage0_61[138], stage0_61[139], stage0_61[140], stage0_61[141]},
      {stage0_63[132], stage0_63[133], stage0_63[134], stage0_63[135], stage0_63[136], stage0_63[137]},
      {stage1_65[22],stage1_64[44],stage1_63[45],stage1_62[58],stage1_61[89]}
   );
   gpc606_5 gpc1211 (
      {stage0_61[142], stage0_61[143], stage0_61[144], stage0_61[145], stage0_61[146], stage0_61[147]},
      {stage0_63[138], stage0_63[139], stage0_63[140], stage0_63[141], stage0_63[142], stage0_63[143]},
      {stage1_65[23],stage1_64[45],stage1_63[46],stage1_62[59],stage1_61[90]}
   );
   gpc606_5 gpc1212 (
      {stage0_61[148], stage0_61[149], stage0_61[150], stage0_61[151], stage0_61[152], stage0_61[153]},
      {stage0_63[144], stage0_63[145], stage0_63[146], stage0_63[147], stage0_63[148], stage0_63[149]},
      {stage1_65[24],stage1_64[46],stage1_63[47],stage1_62[60],stage1_61[91]}
   );
   gpc606_5 gpc1213 (
      {stage0_61[154], stage0_61[155], stage0_61[156], stage0_61[157], stage0_61[158], stage0_61[159]},
      {stage0_63[150], stage0_63[151], stage0_63[152], stage0_63[153], stage0_63[154], stage0_63[155]},
      {stage1_65[25],stage1_64[47],stage1_63[48],stage1_62[61],stage1_61[92]}
   );
   gpc606_5 gpc1214 (
      {stage0_61[160], stage0_61[161], stage0_61[162], stage0_61[163], stage0_61[164], stage0_61[165]},
      {stage0_63[156], stage0_63[157], stage0_63[158], stage0_63[159], stage0_63[160], stage0_63[161]},
      {stage1_65[26],stage1_64[48],stage1_63[49],stage1_62[62],stage1_61[93]}
   );
   gpc606_5 gpc1215 (
      {stage0_61[166], stage0_61[167], stage0_61[168], stage0_61[169], stage0_61[170], stage0_61[171]},
      {stage0_63[162], stage0_63[163], stage0_63[164], stage0_63[165], stage0_63[166], stage0_63[167]},
      {stage1_65[27],stage1_64[49],stage1_63[50],stage1_62[63],stage1_61[94]}
   );
   gpc606_5 gpc1216 (
      {stage0_61[172], stage0_61[173], stage0_61[174], stage0_61[175], stage0_61[176], stage0_61[177]},
      {stage0_63[168], stage0_63[169], stage0_63[170], stage0_63[171], stage0_63[172], stage0_63[173]},
      {stage1_65[28],stage1_64[50],stage1_63[51],stage1_62[64],stage1_61[95]}
   );
   gpc606_5 gpc1217 (
      {stage0_61[178], stage0_61[179], stage0_61[180], stage0_61[181], stage0_61[182], stage0_61[183]},
      {stage0_63[174], stage0_63[175], stage0_63[176], stage0_63[177], stage0_63[178], stage0_63[179]},
      {stage1_65[29],stage1_64[51],stage1_63[52],stage1_62[65],stage1_61[96]}
   );
   gpc606_5 gpc1218 (
      {stage0_61[184], stage0_61[185], stage0_61[186], stage0_61[187], stage0_61[188], stage0_61[189]},
      {stage0_63[180], stage0_63[181], stage0_63[182], stage0_63[183], stage0_63[184], stage0_63[185]},
      {stage1_65[30],stage1_64[52],stage1_63[53],stage1_62[66],stage1_61[97]}
   );
   gpc606_5 gpc1219 (
      {stage0_61[190], stage0_61[191], stage0_61[192], stage0_61[193], stage0_61[194], stage0_61[195]},
      {stage0_63[186], stage0_63[187], stage0_63[188], stage0_63[189], stage0_63[190], stage0_63[191]},
      {stage1_65[31],stage1_64[53],stage1_63[54],stage1_62[67],stage1_61[98]}
   );
   gpc606_5 gpc1220 (
      {stage0_61[196], stage0_61[197], stage0_61[198], stage0_61[199], stage0_61[200], stage0_61[201]},
      {stage0_63[192], stage0_63[193], stage0_63[194], stage0_63[195], stage0_63[196], stage0_63[197]},
      {stage1_65[32],stage1_64[54],stage1_63[55],stage1_62[68],stage1_61[99]}
   );
   gpc606_5 gpc1221 (
      {stage0_61[202], stage0_61[203], stage0_61[204], stage0_61[205], stage0_61[206], stage0_61[207]},
      {stage0_63[198], stage0_63[199], stage0_63[200], stage0_63[201], stage0_63[202], stage0_63[203]},
      {stage1_65[33],stage1_64[55],stage1_63[56],stage1_62[69],stage1_61[100]}
   );
   gpc606_5 gpc1222 (
      {stage0_61[208], stage0_61[209], stage0_61[210], stage0_61[211], stage0_61[212], stage0_61[213]},
      {stage0_63[204], stage0_63[205], stage0_63[206], stage0_63[207], stage0_63[208], stage0_63[209]},
      {stage1_65[34],stage1_64[56],stage1_63[57],stage1_62[70],stage1_61[101]}
   );
   gpc606_5 gpc1223 (
      {stage0_61[214], stage0_61[215], stage0_61[216], stage0_61[217], stage0_61[218], stage0_61[219]},
      {stage0_63[210], stage0_63[211], stage0_63[212], stage0_63[213], stage0_63[214], stage0_63[215]},
      {stage1_65[35],stage1_64[57],stage1_63[58],stage1_62[71],stage1_61[102]}
   );
   gpc606_5 gpc1224 (
      {stage0_61[220], stage0_61[221], stage0_61[222], stage0_61[223], stage0_61[224], stage0_61[225]},
      {stage0_63[216], stage0_63[217], stage0_63[218], stage0_63[219], stage0_63[220], stage0_63[221]},
      {stage1_65[36],stage1_64[58],stage1_63[59],stage1_62[72],stage1_61[103]}
   );
   gpc606_5 gpc1225 (
      {stage0_61[226], stage0_61[227], stage0_61[228], stage0_61[229], stage0_61[230], stage0_61[231]},
      {stage0_63[222], stage0_63[223], stage0_63[224], stage0_63[225], stage0_63[226], stage0_63[227]},
      {stage1_65[37],stage1_64[59],stage1_63[60],stage1_62[73],stage1_61[104]}
   );
   gpc606_5 gpc1226 (
      {stage0_61[232], stage0_61[233], stage0_61[234], stage0_61[235], stage0_61[236], stage0_61[237]},
      {stage0_63[228], stage0_63[229], stage0_63[230], stage0_63[231], stage0_63[232], stage0_63[233]},
      {stage1_65[38],stage1_64[60],stage1_63[61],stage1_62[74],stage1_61[105]}
   );
   gpc606_5 gpc1227 (
      {stage0_61[238], stage0_61[239], stage0_61[240], stage0_61[241], stage0_61[242], stage0_61[243]},
      {stage0_63[234], stage0_63[235], stage0_63[236], stage0_63[237], stage0_63[238], stage0_63[239]},
      {stage1_65[39],stage1_64[61],stage1_63[62],stage1_62[75],stage1_61[106]}
   );
   gpc606_5 gpc1228 (
      {stage0_61[244], stage0_61[245], stage0_61[246], stage0_61[247], stage0_61[248], stage0_61[249]},
      {stage0_63[240], stage0_63[241], stage0_63[242], stage0_63[243], stage0_63[244], stage0_63[245]},
      {stage1_65[40],stage1_64[62],stage1_63[63],stage1_62[76],stage1_61[107]}
   );
   gpc606_5 gpc1229 (
      {stage0_61[250], stage0_61[251], stage0_61[252], stage0_61[253], stage0_61[254], stage0_61[255]},
      {stage0_63[246], stage0_63[247], stage0_63[248], stage0_63[249], stage0_63[250], stage0_63[251]},
      {stage1_65[41],stage1_64[63],stage1_63[64],stage1_62[77],stage1_61[108]}
   );
   gpc1_1 gpc1230 (
      {stage0_0[212]},
      {stage1_0[47]}
   );
   gpc1_1 gpc1231 (
      {stage0_0[213]},
      {stage1_0[48]}
   );
   gpc1_1 gpc1232 (
      {stage0_0[214]},
      {stage1_0[49]}
   );
   gpc1_1 gpc1233 (
      {stage0_0[215]},
      {stage1_0[50]}
   );
   gpc1_1 gpc1234 (
      {stage0_0[216]},
      {stage1_0[51]}
   );
   gpc1_1 gpc1235 (
      {stage0_0[217]},
      {stage1_0[52]}
   );
   gpc1_1 gpc1236 (
      {stage0_0[218]},
      {stage1_0[53]}
   );
   gpc1_1 gpc1237 (
      {stage0_0[219]},
      {stage1_0[54]}
   );
   gpc1_1 gpc1238 (
      {stage0_0[220]},
      {stage1_0[55]}
   );
   gpc1_1 gpc1239 (
      {stage0_0[221]},
      {stage1_0[56]}
   );
   gpc1_1 gpc1240 (
      {stage0_0[222]},
      {stage1_0[57]}
   );
   gpc1_1 gpc1241 (
      {stage0_0[223]},
      {stage1_0[58]}
   );
   gpc1_1 gpc1242 (
      {stage0_0[224]},
      {stage1_0[59]}
   );
   gpc1_1 gpc1243 (
      {stage0_0[225]},
      {stage1_0[60]}
   );
   gpc1_1 gpc1244 (
      {stage0_0[226]},
      {stage1_0[61]}
   );
   gpc1_1 gpc1245 (
      {stage0_0[227]},
      {stage1_0[62]}
   );
   gpc1_1 gpc1246 (
      {stage0_0[228]},
      {stage1_0[63]}
   );
   gpc1_1 gpc1247 (
      {stage0_0[229]},
      {stage1_0[64]}
   );
   gpc1_1 gpc1248 (
      {stage0_0[230]},
      {stage1_0[65]}
   );
   gpc1_1 gpc1249 (
      {stage0_0[231]},
      {stage1_0[66]}
   );
   gpc1_1 gpc1250 (
      {stage0_0[232]},
      {stage1_0[67]}
   );
   gpc1_1 gpc1251 (
      {stage0_0[233]},
      {stage1_0[68]}
   );
   gpc1_1 gpc1252 (
      {stage0_0[234]},
      {stage1_0[69]}
   );
   gpc1_1 gpc1253 (
      {stage0_0[235]},
      {stage1_0[70]}
   );
   gpc1_1 gpc1254 (
      {stage0_0[236]},
      {stage1_0[71]}
   );
   gpc1_1 gpc1255 (
      {stage0_0[237]},
      {stage1_0[72]}
   );
   gpc1_1 gpc1256 (
      {stage0_0[238]},
      {stage1_0[73]}
   );
   gpc1_1 gpc1257 (
      {stage0_0[239]},
      {stage1_0[74]}
   );
   gpc1_1 gpc1258 (
      {stage0_0[240]},
      {stage1_0[75]}
   );
   gpc1_1 gpc1259 (
      {stage0_0[241]},
      {stage1_0[76]}
   );
   gpc1_1 gpc1260 (
      {stage0_0[242]},
      {stage1_0[77]}
   );
   gpc1_1 gpc1261 (
      {stage0_0[243]},
      {stage1_0[78]}
   );
   gpc1_1 gpc1262 (
      {stage0_0[244]},
      {stage1_0[79]}
   );
   gpc1_1 gpc1263 (
      {stage0_0[245]},
      {stage1_0[80]}
   );
   gpc1_1 gpc1264 (
      {stage0_0[246]},
      {stage1_0[81]}
   );
   gpc1_1 gpc1265 (
      {stage0_0[247]},
      {stage1_0[82]}
   );
   gpc1_1 gpc1266 (
      {stage0_0[248]},
      {stage1_0[83]}
   );
   gpc1_1 gpc1267 (
      {stage0_0[249]},
      {stage1_0[84]}
   );
   gpc1_1 gpc1268 (
      {stage0_0[250]},
      {stage1_0[85]}
   );
   gpc1_1 gpc1269 (
      {stage0_0[251]},
      {stage1_0[86]}
   );
   gpc1_1 gpc1270 (
      {stage0_0[252]},
      {stage1_0[87]}
   );
   gpc1_1 gpc1271 (
      {stage0_0[253]},
      {stage1_0[88]}
   );
   gpc1_1 gpc1272 (
      {stage0_0[254]},
      {stage1_0[89]}
   );
   gpc1_1 gpc1273 (
      {stage0_0[255]},
      {stage1_0[90]}
   );
   gpc1_1 gpc1274 (
      {stage0_1[234]},
      {stage1_1[61]}
   );
   gpc1_1 gpc1275 (
      {stage0_1[235]},
      {stage1_1[62]}
   );
   gpc1_1 gpc1276 (
      {stage0_1[236]},
      {stage1_1[63]}
   );
   gpc1_1 gpc1277 (
      {stage0_1[237]},
      {stage1_1[64]}
   );
   gpc1_1 gpc1278 (
      {stage0_1[238]},
      {stage1_1[65]}
   );
   gpc1_1 gpc1279 (
      {stage0_1[239]},
      {stage1_1[66]}
   );
   gpc1_1 gpc1280 (
      {stage0_1[240]},
      {stage1_1[67]}
   );
   gpc1_1 gpc1281 (
      {stage0_1[241]},
      {stage1_1[68]}
   );
   gpc1_1 gpc1282 (
      {stage0_1[242]},
      {stage1_1[69]}
   );
   gpc1_1 gpc1283 (
      {stage0_1[243]},
      {stage1_1[70]}
   );
   gpc1_1 gpc1284 (
      {stage0_1[244]},
      {stage1_1[71]}
   );
   gpc1_1 gpc1285 (
      {stage0_1[245]},
      {stage1_1[72]}
   );
   gpc1_1 gpc1286 (
      {stage0_1[246]},
      {stage1_1[73]}
   );
   gpc1_1 gpc1287 (
      {stage0_1[247]},
      {stage1_1[74]}
   );
   gpc1_1 gpc1288 (
      {stage0_1[248]},
      {stage1_1[75]}
   );
   gpc1_1 gpc1289 (
      {stage0_1[249]},
      {stage1_1[76]}
   );
   gpc1_1 gpc1290 (
      {stage0_1[250]},
      {stage1_1[77]}
   );
   gpc1_1 gpc1291 (
      {stage0_1[251]},
      {stage1_1[78]}
   );
   gpc1_1 gpc1292 (
      {stage0_1[252]},
      {stage1_1[79]}
   );
   gpc1_1 gpc1293 (
      {stage0_1[253]},
      {stage1_1[80]}
   );
   gpc1_1 gpc1294 (
      {stage0_1[254]},
      {stage1_1[81]}
   );
   gpc1_1 gpc1295 (
      {stage0_1[255]},
      {stage1_1[82]}
   );
   gpc1_1 gpc1296 (
      {stage0_2[199]},
      {stage1_2[74]}
   );
   gpc1_1 gpc1297 (
      {stage0_2[200]},
      {stage1_2[75]}
   );
   gpc1_1 gpc1298 (
      {stage0_2[201]},
      {stage1_2[76]}
   );
   gpc1_1 gpc1299 (
      {stage0_2[202]},
      {stage1_2[77]}
   );
   gpc1_1 gpc1300 (
      {stage0_2[203]},
      {stage1_2[78]}
   );
   gpc1_1 gpc1301 (
      {stage0_2[204]},
      {stage1_2[79]}
   );
   gpc1_1 gpc1302 (
      {stage0_2[205]},
      {stage1_2[80]}
   );
   gpc1_1 gpc1303 (
      {stage0_2[206]},
      {stage1_2[81]}
   );
   gpc1_1 gpc1304 (
      {stage0_2[207]},
      {stage1_2[82]}
   );
   gpc1_1 gpc1305 (
      {stage0_2[208]},
      {stage1_2[83]}
   );
   gpc1_1 gpc1306 (
      {stage0_2[209]},
      {stage1_2[84]}
   );
   gpc1_1 gpc1307 (
      {stage0_2[210]},
      {stage1_2[85]}
   );
   gpc1_1 gpc1308 (
      {stage0_2[211]},
      {stage1_2[86]}
   );
   gpc1_1 gpc1309 (
      {stage0_2[212]},
      {stage1_2[87]}
   );
   gpc1_1 gpc1310 (
      {stage0_2[213]},
      {stage1_2[88]}
   );
   gpc1_1 gpc1311 (
      {stage0_2[214]},
      {stage1_2[89]}
   );
   gpc1_1 gpc1312 (
      {stage0_2[215]},
      {stage1_2[90]}
   );
   gpc1_1 gpc1313 (
      {stage0_2[216]},
      {stage1_2[91]}
   );
   gpc1_1 gpc1314 (
      {stage0_2[217]},
      {stage1_2[92]}
   );
   gpc1_1 gpc1315 (
      {stage0_2[218]},
      {stage1_2[93]}
   );
   gpc1_1 gpc1316 (
      {stage0_2[219]},
      {stage1_2[94]}
   );
   gpc1_1 gpc1317 (
      {stage0_2[220]},
      {stage1_2[95]}
   );
   gpc1_1 gpc1318 (
      {stage0_2[221]},
      {stage1_2[96]}
   );
   gpc1_1 gpc1319 (
      {stage0_2[222]},
      {stage1_2[97]}
   );
   gpc1_1 gpc1320 (
      {stage0_2[223]},
      {stage1_2[98]}
   );
   gpc1_1 gpc1321 (
      {stage0_2[224]},
      {stage1_2[99]}
   );
   gpc1_1 gpc1322 (
      {stage0_2[225]},
      {stage1_2[100]}
   );
   gpc1_1 gpc1323 (
      {stage0_2[226]},
      {stage1_2[101]}
   );
   gpc1_1 gpc1324 (
      {stage0_2[227]},
      {stage1_2[102]}
   );
   gpc1_1 gpc1325 (
      {stage0_2[228]},
      {stage1_2[103]}
   );
   gpc1_1 gpc1326 (
      {stage0_2[229]},
      {stage1_2[104]}
   );
   gpc1_1 gpc1327 (
      {stage0_2[230]},
      {stage1_2[105]}
   );
   gpc1_1 gpc1328 (
      {stage0_2[231]},
      {stage1_2[106]}
   );
   gpc1_1 gpc1329 (
      {stage0_2[232]},
      {stage1_2[107]}
   );
   gpc1_1 gpc1330 (
      {stage0_2[233]},
      {stage1_2[108]}
   );
   gpc1_1 gpc1331 (
      {stage0_2[234]},
      {stage1_2[109]}
   );
   gpc1_1 gpc1332 (
      {stage0_2[235]},
      {stage1_2[110]}
   );
   gpc1_1 gpc1333 (
      {stage0_2[236]},
      {stage1_2[111]}
   );
   gpc1_1 gpc1334 (
      {stage0_2[237]},
      {stage1_2[112]}
   );
   gpc1_1 gpc1335 (
      {stage0_2[238]},
      {stage1_2[113]}
   );
   gpc1_1 gpc1336 (
      {stage0_2[239]},
      {stage1_2[114]}
   );
   gpc1_1 gpc1337 (
      {stage0_2[240]},
      {stage1_2[115]}
   );
   gpc1_1 gpc1338 (
      {stage0_2[241]},
      {stage1_2[116]}
   );
   gpc1_1 gpc1339 (
      {stage0_2[242]},
      {stage1_2[117]}
   );
   gpc1_1 gpc1340 (
      {stage0_2[243]},
      {stage1_2[118]}
   );
   gpc1_1 gpc1341 (
      {stage0_2[244]},
      {stage1_2[119]}
   );
   gpc1_1 gpc1342 (
      {stage0_2[245]},
      {stage1_2[120]}
   );
   gpc1_1 gpc1343 (
      {stage0_2[246]},
      {stage1_2[121]}
   );
   gpc1_1 gpc1344 (
      {stage0_2[247]},
      {stage1_2[122]}
   );
   gpc1_1 gpc1345 (
      {stage0_2[248]},
      {stage1_2[123]}
   );
   gpc1_1 gpc1346 (
      {stage0_2[249]},
      {stage1_2[124]}
   );
   gpc1_1 gpc1347 (
      {stage0_2[250]},
      {stage1_2[125]}
   );
   gpc1_1 gpc1348 (
      {stage0_2[251]},
      {stage1_2[126]}
   );
   gpc1_1 gpc1349 (
      {stage0_2[252]},
      {stage1_2[127]}
   );
   gpc1_1 gpc1350 (
      {stage0_2[253]},
      {stage1_2[128]}
   );
   gpc1_1 gpc1351 (
      {stage0_2[254]},
      {stage1_2[129]}
   );
   gpc1_1 gpc1352 (
      {stage0_2[255]},
      {stage1_2[130]}
   );
   gpc1_1 gpc1353 (
      {stage0_3[245]},
      {stage1_3[96]}
   );
   gpc1_1 gpc1354 (
      {stage0_3[246]},
      {stage1_3[97]}
   );
   gpc1_1 gpc1355 (
      {stage0_3[247]},
      {stage1_3[98]}
   );
   gpc1_1 gpc1356 (
      {stage0_3[248]},
      {stage1_3[99]}
   );
   gpc1_1 gpc1357 (
      {stage0_3[249]},
      {stage1_3[100]}
   );
   gpc1_1 gpc1358 (
      {stage0_3[250]},
      {stage1_3[101]}
   );
   gpc1_1 gpc1359 (
      {stage0_3[251]},
      {stage1_3[102]}
   );
   gpc1_1 gpc1360 (
      {stage0_3[252]},
      {stage1_3[103]}
   );
   gpc1_1 gpc1361 (
      {stage0_3[253]},
      {stage1_3[104]}
   );
   gpc1_1 gpc1362 (
      {stage0_3[254]},
      {stage1_3[105]}
   );
   gpc1_1 gpc1363 (
      {stage0_3[255]},
      {stage1_3[106]}
   );
   gpc1_1 gpc1364 (
      {stage0_6[236]},
      {stage1_6[96]}
   );
   gpc1_1 gpc1365 (
      {stage0_6[237]},
      {stage1_6[97]}
   );
   gpc1_1 gpc1366 (
      {stage0_6[238]},
      {stage1_6[98]}
   );
   gpc1_1 gpc1367 (
      {stage0_6[239]},
      {stage1_6[99]}
   );
   gpc1_1 gpc1368 (
      {stage0_6[240]},
      {stage1_6[100]}
   );
   gpc1_1 gpc1369 (
      {stage0_6[241]},
      {stage1_6[101]}
   );
   gpc1_1 gpc1370 (
      {stage0_6[242]},
      {stage1_6[102]}
   );
   gpc1_1 gpc1371 (
      {stage0_6[243]},
      {stage1_6[103]}
   );
   gpc1_1 gpc1372 (
      {stage0_6[244]},
      {stage1_6[104]}
   );
   gpc1_1 gpc1373 (
      {stage0_6[245]},
      {stage1_6[105]}
   );
   gpc1_1 gpc1374 (
      {stage0_6[246]},
      {stage1_6[106]}
   );
   gpc1_1 gpc1375 (
      {stage0_6[247]},
      {stage1_6[107]}
   );
   gpc1_1 gpc1376 (
      {stage0_6[248]},
      {stage1_6[108]}
   );
   gpc1_1 gpc1377 (
      {stage0_6[249]},
      {stage1_6[109]}
   );
   gpc1_1 gpc1378 (
      {stage0_6[250]},
      {stage1_6[110]}
   );
   gpc1_1 gpc1379 (
      {stage0_6[251]},
      {stage1_6[111]}
   );
   gpc1_1 gpc1380 (
      {stage0_6[252]},
      {stage1_6[112]}
   );
   gpc1_1 gpc1381 (
      {stage0_6[253]},
      {stage1_6[113]}
   );
   gpc1_1 gpc1382 (
      {stage0_6[254]},
      {stage1_6[114]}
   );
   gpc1_1 gpc1383 (
      {stage0_6[255]},
      {stage1_6[115]}
   );
   gpc1_1 gpc1384 (
      {stage0_7[251]},
      {stage1_7[105]}
   );
   gpc1_1 gpc1385 (
      {stage0_7[252]},
      {stage1_7[106]}
   );
   gpc1_1 gpc1386 (
      {stage0_7[253]},
      {stage1_7[107]}
   );
   gpc1_1 gpc1387 (
      {stage0_7[254]},
      {stage1_7[108]}
   );
   gpc1_1 gpc1388 (
      {stage0_7[255]},
      {stage1_7[109]}
   );
   gpc1_1 gpc1389 (
      {stage0_8[233]},
      {stage1_8[109]}
   );
   gpc1_1 gpc1390 (
      {stage0_8[234]},
      {stage1_8[110]}
   );
   gpc1_1 gpc1391 (
      {stage0_8[235]},
      {stage1_8[111]}
   );
   gpc1_1 gpc1392 (
      {stage0_8[236]},
      {stage1_8[112]}
   );
   gpc1_1 gpc1393 (
      {stage0_8[237]},
      {stage1_8[113]}
   );
   gpc1_1 gpc1394 (
      {stage0_8[238]},
      {stage1_8[114]}
   );
   gpc1_1 gpc1395 (
      {stage0_8[239]},
      {stage1_8[115]}
   );
   gpc1_1 gpc1396 (
      {stage0_8[240]},
      {stage1_8[116]}
   );
   gpc1_1 gpc1397 (
      {stage0_8[241]},
      {stage1_8[117]}
   );
   gpc1_1 gpc1398 (
      {stage0_8[242]},
      {stage1_8[118]}
   );
   gpc1_1 gpc1399 (
      {stage0_8[243]},
      {stage1_8[119]}
   );
   gpc1_1 gpc1400 (
      {stage0_8[244]},
      {stage1_8[120]}
   );
   gpc1_1 gpc1401 (
      {stage0_8[245]},
      {stage1_8[121]}
   );
   gpc1_1 gpc1402 (
      {stage0_8[246]},
      {stage1_8[122]}
   );
   gpc1_1 gpc1403 (
      {stage0_8[247]},
      {stage1_8[123]}
   );
   gpc1_1 gpc1404 (
      {stage0_8[248]},
      {stage1_8[124]}
   );
   gpc1_1 gpc1405 (
      {stage0_8[249]},
      {stage1_8[125]}
   );
   gpc1_1 gpc1406 (
      {stage0_8[250]},
      {stage1_8[126]}
   );
   gpc1_1 gpc1407 (
      {stage0_8[251]},
      {stage1_8[127]}
   );
   gpc1_1 gpc1408 (
      {stage0_8[252]},
      {stage1_8[128]}
   );
   gpc1_1 gpc1409 (
      {stage0_8[253]},
      {stage1_8[129]}
   );
   gpc1_1 gpc1410 (
      {stage0_8[254]},
      {stage1_8[130]}
   );
   gpc1_1 gpc1411 (
      {stage0_8[255]},
      {stage1_8[131]}
   );
   gpc1_1 gpc1412 (
      {stage0_9[235]},
      {stage1_9[99]}
   );
   gpc1_1 gpc1413 (
      {stage0_9[236]},
      {stage1_9[100]}
   );
   gpc1_1 gpc1414 (
      {stage0_9[237]},
      {stage1_9[101]}
   );
   gpc1_1 gpc1415 (
      {stage0_9[238]},
      {stage1_9[102]}
   );
   gpc1_1 gpc1416 (
      {stage0_9[239]},
      {stage1_9[103]}
   );
   gpc1_1 gpc1417 (
      {stage0_9[240]},
      {stage1_9[104]}
   );
   gpc1_1 gpc1418 (
      {stage0_9[241]},
      {stage1_9[105]}
   );
   gpc1_1 gpc1419 (
      {stage0_9[242]},
      {stage1_9[106]}
   );
   gpc1_1 gpc1420 (
      {stage0_9[243]},
      {stage1_9[107]}
   );
   gpc1_1 gpc1421 (
      {stage0_9[244]},
      {stage1_9[108]}
   );
   gpc1_1 gpc1422 (
      {stage0_9[245]},
      {stage1_9[109]}
   );
   gpc1_1 gpc1423 (
      {stage0_9[246]},
      {stage1_9[110]}
   );
   gpc1_1 gpc1424 (
      {stage0_9[247]},
      {stage1_9[111]}
   );
   gpc1_1 gpc1425 (
      {stage0_9[248]},
      {stage1_9[112]}
   );
   gpc1_1 gpc1426 (
      {stage0_9[249]},
      {stage1_9[113]}
   );
   gpc1_1 gpc1427 (
      {stage0_9[250]},
      {stage1_9[114]}
   );
   gpc1_1 gpc1428 (
      {stage0_9[251]},
      {stage1_9[115]}
   );
   gpc1_1 gpc1429 (
      {stage0_9[252]},
      {stage1_9[116]}
   );
   gpc1_1 gpc1430 (
      {stage0_9[253]},
      {stage1_9[117]}
   );
   gpc1_1 gpc1431 (
      {stage0_9[254]},
      {stage1_9[118]}
   );
   gpc1_1 gpc1432 (
      {stage0_9[255]},
      {stage1_9[119]}
   );
   gpc1_1 gpc1433 (
      {stage0_10[181]},
      {stage1_10[81]}
   );
   gpc1_1 gpc1434 (
      {stage0_10[182]},
      {stage1_10[82]}
   );
   gpc1_1 gpc1435 (
      {stage0_10[183]},
      {stage1_10[83]}
   );
   gpc1_1 gpc1436 (
      {stage0_10[184]},
      {stage1_10[84]}
   );
   gpc1_1 gpc1437 (
      {stage0_10[185]},
      {stage1_10[85]}
   );
   gpc1_1 gpc1438 (
      {stage0_10[186]},
      {stage1_10[86]}
   );
   gpc1_1 gpc1439 (
      {stage0_10[187]},
      {stage1_10[87]}
   );
   gpc1_1 gpc1440 (
      {stage0_10[188]},
      {stage1_10[88]}
   );
   gpc1_1 gpc1441 (
      {stage0_10[189]},
      {stage1_10[89]}
   );
   gpc1_1 gpc1442 (
      {stage0_10[190]},
      {stage1_10[90]}
   );
   gpc1_1 gpc1443 (
      {stage0_10[191]},
      {stage1_10[91]}
   );
   gpc1_1 gpc1444 (
      {stage0_10[192]},
      {stage1_10[92]}
   );
   gpc1_1 gpc1445 (
      {stage0_10[193]},
      {stage1_10[93]}
   );
   gpc1_1 gpc1446 (
      {stage0_10[194]},
      {stage1_10[94]}
   );
   gpc1_1 gpc1447 (
      {stage0_10[195]},
      {stage1_10[95]}
   );
   gpc1_1 gpc1448 (
      {stage0_10[196]},
      {stage1_10[96]}
   );
   gpc1_1 gpc1449 (
      {stage0_10[197]},
      {stage1_10[97]}
   );
   gpc1_1 gpc1450 (
      {stage0_10[198]},
      {stage1_10[98]}
   );
   gpc1_1 gpc1451 (
      {stage0_10[199]},
      {stage1_10[99]}
   );
   gpc1_1 gpc1452 (
      {stage0_10[200]},
      {stage1_10[100]}
   );
   gpc1_1 gpc1453 (
      {stage0_10[201]},
      {stage1_10[101]}
   );
   gpc1_1 gpc1454 (
      {stage0_10[202]},
      {stage1_10[102]}
   );
   gpc1_1 gpc1455 (
      {stage0_10[203]},
      {stage1_10[103]}
   );
   gpc1_1 gpc1456 (
      {stage0_10[204]},
      {stage1_10[104]}
   );
   gpc1_1 gpc1457 (
      {stage0_10[205]},
      {stage1_10[105]}
   );
   gpc1_1 gpc1458 (
      {stage0_10[206]},
      {stage1_10[106]}
   );
   gpc1_1 gpc1459 (
      {stage0_10[207]},
      {stage1_10[107]}
   );
   gpc1_1 gpc1460 (
      {stage0_10[208]},
      {stage1_10[108]}
   );
   gpc1_1 gpc1461 (
      {stage0_10[209]},
      {stage1_10[109]}
   );
   gpc1_1 gpc1462 (
      {stage0_10[210]},
      {stage1_10[110]}
   );
   gpc1_1 gpc1463 (
      {stage0_10[211]},
      {stage1_10[111]}
   );
   gpc1_1 gpc1464 (
      {stage0_10[212]},
      {stage1_10[112]}
   );
   gpc1_1 gpc1465 (
      {stage0_10[213]},
      {stage1_10[113]}
   );
   gpc1_1 gpc1466 (
      {stage0_10[214]},
      {stage1_10[114]}
   );
   gpc1_1 gpc1467 (
      {stage0_10[215]},
      {stage1_10[115]}
   );
   gpc1_1 gpc1468 (
      {stage0_10[216]},
      {stage1_10[116]}
   );
   gpc1_1 gpc1469 (
      {stage0_10[217]},
      {stage1_10[117]}
   );
   gpc1_1 gpc1470 (
      {stage0_10[218]},
      {stage1_10[118]}
   );
   gpc1_1 gpc1471 (
      {stage0_10[219]},
      {stage1_10[119]}
   );
   gpc1_1 gpc1472 (
      {stage0_10[220]},
      {stage1_10[120]}
   );
   gpc1_1 gpc1473 (
      {stage0_10[221]},
      {stage1_10[121]}
   );
   gpc1_1 gpc1474 (
      {stage0_10[222]},
      {stage1_10[122]}
   );
   gpc1_1 gpc1475 (
      {stage0_10[223]},
      {stage1_10[123]}
   );
   gpc1_1 gpc1476 (
      {stage0_10[224]},
      {stage1_10[124]}
   );
   gpc1_1 gpc1477 (
      {stage0_10[225]},
      {stage1_10[125]}
   );
   gpc1_1 gpc1478 (
      {stage0_10[226]},
      {stage1_10[126]}
   );
   gpc1_1 gpc1479 (
      {stage0_10[227]},
      {stage1_10[127]}
   );
   gpc1_1 gpc1480 (
      {stage0_10[228]},
      {stage1_10[128]}
   );
   gpc1_1 gpc1481 (
      {stage0_10[229]},
      {stage1_10[129]}
   );
   gpc1_1 gpc1482 (
      {stage0_10[230]},
      {stage1_10[130]}
   );
   gpc1_1 gpc1483 (
      {stage0_10[231]},
      {stage1_10[131]}
   );
   gpc1_1 gpc1484 (
      {stage0_10[232]},
      {stage1_10[132]}
   );
   gpc1_1 gpc1485 (
      {stage0_10[233]},
      {stage1_10[133]}
   );
   gpc1_1 gpc1486 (
      {stage0_10[234]},
      {stage1_10[134]}
   );
   gpc1_1 gpc1487 (
      {stage0_10[235]},
      {stage1_10[135]}
   );
   gpc1_1 gpc1488 (
      {stage0_10[236]},
      {stage1_10[136]}
   );
   gpc1_1 gpc1489 (
      {stage0_10[237]},
      {stage1_10[137]}
   );
   gpc1_1 gpc1490 (
      {stage0_10[238]},
      {stage1_10[138]}
   );
   gpc1_1 gpc1491 (
      {stage0_10[239]},
      {stage1_10[139]}
   );
   gpc1_1 gpc1492 (
      {stage0_10[240]},
      {stage1_10[140]}
   );
   gpc1_1 gpc1493 (
      {stage0_10[241]},
      {stage1_10[141]}
   );
   gpc1_1 gpc1494 (
      {stage0_10[242]},
      {stage1_10[142]}
   );
   gpc1_1 gpc1495 (
      {stage0_10[243]},
      {stage1_10[143]}
   );
   gpc1_1 gpc1496 (
      {stage0_10[244]},
      {stage1_10[144]}
   );
   gpc1_1 gpc1497 (
      {stage0_10[245]},
      {stage1_10[145]}
   );
   gpc1_1 gpc1498 (
      {stage0_10[246]},
      {stage1_10[146]}
   );
   gpc1_1 gpc1499 (
      {stage0_10[247]},
      {stage1_10[147]}
   );
   gpc1_1 gpc1500 (
      {stage0_10[248]},
      {stage1_10[148]}
   );
   gpc1_1 gpc1501 (
      {stage0_10[249]},
      {stage1_10[149]}
   );
   gpc1_1 gpc1502 (
      {stage0_10[250]},
      {stage1_10[150]}
   );
   gpc1_1 gpc1503 (
      {stage0_10[251]},
      {stage1_10[151]}
   );
   gpc1_1 gpc1504 (
      {stage0_10[252]},
      {stage1_10[152]}
   );
   gpc1_1 gpc1505 (
      {stage0_10[253]},
      {stage1_10[153]}
   );
   gpc1_1 gpc1506 (
      {stage0_10[254]},
      {stage1_10[154]}
   );
   gpc1_1 gpc1507 (
      {stage0_10[255]},
      {stage1_10[155]}
   );
   gpc1_1 gpc1508 (
      {stage0_11[183]},
      {stage1_11[81]}
   );
   gpc1_1 gpc1509 (
      {stage0_11[184]},
      {stage1_11[82]}
   );
   gpc1_1 gpc1510 (
      {stage0_11[185]},
      {stage1_11[83]}
   );
   gpc1_1 gpc1511 (
      {stage0_11[186]},
      {stage1_11[84]}
   );
   gpc1_1 gpc1512 (
      {stage0_11[187]},
      {stage1_11[85]}
   );
   gpc1_1 gpc1513 (
      {stage0_11[188]},
      {stage1_11[86]}
   );
   gpc1_1 gpc1514 (
      {stage0_11[189]},
      {stage1_11[87]}
   );
   gpc1_1 gpc1515 (
      {stage0_11[190]},
      {stage1_11[88]}
   );
   gpc1_1 gpc1516 (
      {stage0_11[191]},
      {stage1_11[89]}
   );
   gpc1_1 gpc1517 (
      {stage0_11[192]},
      {stage1_11[90]}
   );
   gpc1_1 gpc1518 (
      {stage0_11[193]},
      {stage1_11[91]}
   );
   gpc1_1 gpc1519 (
      {stage0_11[194]},
      {stage1_11[92]}
   );
   gpc1_1 gpc1520 (
      {stage0_11[195]},
      {stage1_11[93]}
   );
   gpc1_1 gpc1521 (
      {stage0_11[196]},
      {stage1_11[94]}
   );
   gpc1_1 gpc1522 (
      {stage0_11[197]},
      {stage1_11[95]}
   );
   gpc1_1 gpc1523 (
      {stage0_11[198]},
      {stage1_11[96]}
   );
   gpc1_1 gpc1524 (
      {stage0_11[199]},
      {stage1_11[97]}
   );
   gpc1_1 gpc1525 (
      {stage0_11[200]},
      {stage1_11[98]}
   );
   gpc1_1 gpc1526 (
      {stage0_11[201]},
      {stage1_11[99]}
   );
   gpc1_1 gpc1527 (
      {stage0_11[202]},
      {stage1_11[100]}
   );
   gpc1_1 gpc1528 (
      {stage0_11[203]},
      {stage1_11[101]}
   );
   gpc1_1 gpc1529 (
      {stage0_11[204]},
      {stage1_11[102]}
   );
   gpc1_1 gpc1530 (
      {stage0_11[205]},
      {stage1_11[103]}
   );
   gpc1_1 gpc1531 (
      {stage0_11[206]},
      {stage1_11[104]}
   );
   gpc1_1 gpc1532 (
      {stage0_11[207]},
      {stage1_11[105]}
   );
   gpc1_1 gpc1533 (
      {stage0_11[208]},
      {stage1_11[106]}
   );
   gpc1_1 gpc1534 (
      {stage0_11[209]},
      {stage1_11[107]}
   );
   gpc1_1 gpc1535 (
      {stage0_11[210]},
      {stage1_11[108]}
   );
   gpc1_1 gpc1536 (
      {stage0_11[211]},
      {stage1_11[109]}
   );
   gpc1_1 gpc1537 (
      {stage0_11[212]},
      {stage1_11[110]}
   );
   gpc1_1 gpc1538 (
      {stage0_11[213]},
      {stage1_11[111]}
   );
   gpc1_1 gpc1539 (
      {stage0_11[214]},
      {stage1_11[112]}
   );
   gpc1_1 gpc1540 (
      {stage0_11[215]},
      {stage1_11[113]}
   );
   gpc1_1 gpc1541 (
      {stage0_11[216]},
      {stage1_11[114]}
   );
   gpc1_1 gpc1542 (
      {stage0_11[217]},
      {stage1_11[115]}
   );
   gpc1_1 gpc1543 (
      {stage0_11[218]},
      {stage1_11[116]}
   );
   gpc1_1 gpc1544 (
      {stage0_11[219]},
      {stage1_11[117]}
   );
   gpc1_1 gpc1545 (
      {stage0_11[220]},
      {stage1_11[118]}
   );
   gpc1_1 gpc1546 (
      {stage0_11[221]},
      {stage1_11[119]}
   );
   gpc1_1 gpc1547 (
      {stage0_11[222]},
      {stage1_11[120]}
   );
   gpc1_1 gpc1548 (
      {stage0_11[223]},
      {stage1_11[121]}
   );
   gpc1_1 gpc1549 (
      {stage0_11[224]},
      {stage1_11[122]}
   );
   gpc1_1 gpc1550 (
      {stage0_11[225]},
      {stage1_11[123]}
   );
   gpc1_1 gpc1551 (
      {stage0_11[226]},
      {stage1_11[124]}
   );
   gpc1_1 gpc1552 (
      {stage0_11[227]},
      {stage1_11[125]}
   );
   gpc1_1 gpc1553 (
      {stage0_11[228]},
      {stage1_11[126]}
   );
   gpc1_1 gpc1554 (
      {stage0_11[229]},
      {stage1_11[127]}
   );
   gpc1_1 gpc1555 (
      {stage0_11[230]},
      {stage1_11[128]}
   );
   gpc1_1 gpc1556 (
      {stage0_11[231]},
      {stage1_11[129]}
   );
   gpc1_1 gpc1557 (
      {stage0_11[232]},
      {stage1_11[130]}
   );
   gpc1_1 gpc1558 (
      {stage0_11[233]},
      {stage1_11[131]}
   );
   gpc1_1 gpc1559 (
      {stage0_11[234]},
      {stage1_11[132]}
   );
   gpc1_1 gpc1560 (
      {stage0_11[235]},
      {stage1_11[133]}
   );
   gpc1_1 gpc1561 (
      {stage0_11[236]},
      {stage1_11[134]}
   );
   gpc1_1 gpc1562 (
      {stage0_11[237]},
      {stage1_11[135]}
   );
   gpc1_1 gpc1563 (
      {stage0_11[238]},
      {stage1_11[136]}
   );
   gpc1_1 gpc1564 (
      {stage0_11[239]},
      {stage1_11[137]}
   );
   gpc1_1 gpc1565 (
      {stage0_11[240]},
      {stage1_11[138]}
   );
   gpc1_1 gpc1566 (
      {stage0_11[241]},
      {stage1_11[139]}
   );
   gpc1_1 gpc1567 (
      {stage0_11[242]},
      {stage1_11[140]}
   );
   gpc1_1 gpc1568 (
      {stage0_11[243]},
      {stage1_11[141]}
   );
   gpc1_1 gpc1569 (
      {stage0_11[244]},
      {stage1_11[142]}
   );
   gpc1_1 gpc1570 (
      {stage0_11[245]},
      {stage1_11[143]}
   );
   gpc1_1 gpc1571 (
      {stage0_11[246]},
      {stage1_11[144]}
   );
   gpc1_1 gpc1572 (
      {stage0_11[247]},
      {stage1_11[145]}
   );
   gpc1_1 gpc1573 (
      {stage0_11[248]},
      {stage1_11[146]}
   );
   gpc1_1 gpc1574 (
      {stage0_11[249]},
      {stage1_11[147]}
   );
   gpc1_1 gpc1575 (
      {stage0_11[250]},
      {stage1_11[148]}
   );
   gpc1_1 gpc1576 (
      {stage0_11[251]},
      {stage1_11[149]}
   );
   gpc1_1 gpc1577 (
      {stage0_11[252]},
      {stage1_11[150]}
   );
   gpc1_1 gpc1578 (
      {stage0_11[253]},
      {stage1_11[151]}
   );
   gpc1_1 gpc1579 (
      {stage0_11[254]},
      {stage1_11[152]}
   );
   gpc1_1 gpc1580 (
      {stage0_11[255]},
      {stage1_11[153]}
   );
   gpc1_1 gpc1581 (
      {stage0_12[220]},
      {stage1_12[97]}
   );
   gpc1_1 gpc1582 (
      {stage0_12[221]},
      {stage1_12[98]}
   );
   gpc1_1 gpc1583 (
      {stage0_12[222]},
      {stage1_12[99]}
   );
   gpc1_1 gpc1584 (
      {stage0_12[223]},
      {stage1_12[100]}
   );
   gpc1_1 gpc1585 (
      {stage0_12[224]},
      {stage1_12[101]}
   );
   gpc1_1 gpc1586 (
      {stage0_12[225]},
      {stage1_12[102]}
   );
   gpc1_1 gpc1587 (
      {stage0_12[226]},
      {stage1_12[103]}
   );
   gpc1_1 gpc1588 (
      {stage0_12[227]},
      {stage1_12[104]}
   );
   gpc1_1 gpc1589 (
      {stage0_12[228]},
      {stage1_12[105]}
   );
   gpc1_1 gpc1590 (
      {stage0_12[229]},
      {stage1_12[106]}
   );
   gpc1_1 gpc1591 (
      {stage0_12[230]},
      {stage1_12[107]}
   );
   gpc1_1 gpc1592 (
      {stage0_12[231]},
      {stage1_12[108]}
   );
   gpc1_1 gpc1593 (
      {stage0_12[232]},
      {stage1_12[109]}
   );
   gpc1_1 gpc1594 (
      {stage0_12[233]},
      {stage1_12[110]}
   );
   gpc1_1 gpc1595 (
      {stage0_12[234]},
      {stage1_12[111]}
   );
   gpc1_1 gpc1596 (
      {stage0_12[235]},
      {stage1_12[112]}
   );
   gpc1_1 gpc1597 (
      {stage0_12[236]},
      {stage1_12[113]}
   );
   gpc1_1 gpc1598 (
      {stage0_12[237]},
      {stage1_12[114]}
   );
   gpc1_1 gpc1599 (
      {stage0_12[238]},
      {stage1_12[115]}
   );
   gpc1_1 gpc1600 (
      {stage0_12[239]},
      {stage1_12[116]}
   );
   gpc1_1 gpc1601 (
      {stage0_12[240]},
      {stage1_12[117]}
   );
   gpc1_1 gpc1602 (
      {stage0_12[241]},
      {stage1_12[118]}
   );
   gpc1_1 gpc1603 (
      {stage0_12[242]},
      {stage1_12[119]}
   );
   gpc1_1 gpc1604 (
      {stage0_12[243]},
      {stage1_12[120]}
   );
   gpc1_1 gpc1605 (
      {stage0_12[244]},
      {stage1_12[121]}
   );
   gpc1_1 gpc1606 (
      {stage0_12[245]},
      {stage1_12[122]}
   );
   gpc1_1 gpc1607 (
      {stage0_12[246]},
      {stage1_12[123]}
   );
   gpc1_1 gpc1608 (
      {stage0_12[247]},
      {stage1_12[124]}
   );
   gpc1_1 gpc1609 (
      {stage0_12[248]},
      {stage1_12[125]}
   );
   gpc1_1 gpc1610 (
      {stage0_12[249]},
      {stage1_12[126]}
   );
   gpc1_1 gpc1611 (
      {stage0_12[250]},
      {stage1_12[127]}
   );
   gpc1_1 gpc1612 (
      {stage0_12[251]},
      {stage1_12[128]}
   );
   gpc1_1 gpc1613 (
      {stage0_12[252]},
      {stage1_12[129]}
   );
   gpc1_1 gpc1614 (
      {stage0_12[253]},
      {stage1_12[130]}
   );
   gpc1_1 gpc1615 (
      {stage0_12[254]},
      {stage1_12[131]}
   );
   gpc1_1 gpc1616 (
      {stage0_12[255]},
      {stage1_12[132]}
   );
   gpc1_1 gpc1617 (
      {stage0_13[254]},
      {stage1_13[95]}
   );
   gpc1_1 gpc1618 (
      {stage0_13[255]},
      {stage1_13[96]}
   );
   gpc1_1 gpc1619 (
      {stage0_15[220]},
      {stage1_15[96]}
   );
   gpc1_1 gpc1620 (
      {stage0_15[221]},
      {stage1_15[97]}
   );
   gpc1_1 gpc1621 (
      {stage0_15[222]},
      {stage1_15[98]}
   );
   gpc1_1 gpc1622 (
      {stage0_15[223]},
      {stage1_15[99]}
   );
   gpc1_1 gpc1623 (
      {stage0_15[224]},
      {stage1_15[100]}
   );
   gpc1_1 gpc1624 (
      {stage0_15[225]},
      {stage1_15[101]}
   );
   gpc1_1 gpc1625 (
      {stage0_15[226]},
      {stage1_15[102]}
   );
   gpc1_1 gpc1626 (
      {stage0_15[227]},
      {stage1_15[103]}
   );
   gpc1_1 gpc1627 (
      {stage0_15[228]},
      {stage1_15[104]}
   );
   gpc1_1 gpc1628 (
      {stage0_15[229]},
      {stage1_15[105]}
   );
   gpc1_1 gpc1629 (
      {stage0_15[230]},
      {stage1_15[106]}
   );
   gpc1_1 gpc1630 (
      {stage0_15[231]},
      {stage1_15[107]}
   );
   gpc1_1 gpc1631 (
      {stage0_15[232]},
      {stage1_15[108]}
   );
   gpc1_1 gpc1632 (
      {stage0_15[233]},
      {stage1_15[109]}
   );
   gpc1_1 gpc1633 (
      {stage0_15[234]},
      {stage1_15[110]}
   );
   gpc1_1 gpc1634 (
      {stage0_15[235]},
      {stage1_15[111]}
   );
   gpc1_1 gpc1635 (
      {stage0_15[236]},
      {stage1_15[112]}
   );
   gpc1_1 gpc1636 (
      {stage0_15[237]},
      {stage1_15[113]}
   );
   gpc1_1 gpc1637 (
      {stage0_15[238]},
      {stage1_15[114]}
   );
   gpc1_1 gpc1638 (
      {stage0_15[239]},
      {stage1_15[115]}
   );
   gpc1_1 gpc1639 (
      {stage0_15[240]},
      {stage1_15[116]}
   );
   gpc1_1 gpc1640 (
      {stage0_15[241]},
      {stage1_15[117]}
   );
   gpc1_1 gpc1641 (
      {stage0_15[242]},
      {stage1_15[118]}
   );
   gpc1_1 gpc1642 (
      {stage0_15[243]},
      {stage1_15[119]}
   );
   gpc1_1 gpc1643 (
      {stage0_15[244]},
      {stage1_15[120]}
   );
   gpc1_1 gpc1644 (
      {stage0_15[245]},
      {stage1_15[121]}
   );
   gpc1_1 gpc1645 (
      {stage0_15[246]},
      {stage1_15[122]}
   );
   gpc1_1 gpc1646 (
      {stage0_15[247]},
      {stage1_15[123]}
   );
   gpc1_1 gpc1647 (
      {stage0_15[248]},
      {stage1_15[124]}
   );
   gpc1_1 gpc1648 (
      {stage0_15[249]},
      {stage1_15[125]}
   );
   gpc1_1 gpc1649 (
      {stage0_15[250]},
      {stage1_15[126]}
   );
   gpc1_1 gpc1650 (
      {stage0_15[251]},
      {stage1_15[127]}
   );
   gpc1_1 gpc1651 (
      {stage0_15[252]},
      {stage1_15[128]}
   );
   gpc1_1 gpc1652 (
      {stage0_15[253]},
      {stage1_15[129]}
   );
   gpc1_1 gpc1653 (
      {stage0_15[254]},
      {stage1_15[130]}
   );
   gpc1_1 gpc1654 (
      {stage0_15[255]},
      {stage1_15[131]}
   );
   gpc1_1 gpc1655 (
      {stage0_16[255]},
      {stage1_16[119]}
   );
   gpc1_1 gpc1656 (
      {stage0_17[251]},
      {stage1_17[106]}
   );
   gpc1_1 gpc1657 (
      {stage0_17[252]},
      {stage1_17[107]}
   );
   gpc1_1 gpc1658 (
      {stage0_17[253]},
      {stage1_17[108]}
   );
   gpc1_1 gpc1659 (
      {stage0_17[254]},
      {stage1_17[109]}
   );
   gpc1_1 gpc1660 (
      {stage0_17[255]},
      {stage1_17[110]}
   );
   gpc1_1 gpc1661 (
      {stage0_18[242]},
      {stage1_18[86]}
   );
   gpc1_1 gpc1662 (
      {stage0_18[243]},
      {stage1_18[87]}
   );
   gpc1_1 gpc1663 (
      {stage0_18[244]},
      {stage1_18[88]}
   );
   gpc1_1 gpc1664 (
      {stage0_18[245]},
      {stage1_18[89]}
   );
   gpc1_1 gpc1665 (
      {stage0_18[246]},
      {stage1_18[90]}
   );
   gpc1_1 gpc1666 (
      {stage0_18[247]},
      {stage1_18[91]}
   );
   gpc1_1 gpc1667 (
      {stage0_18[248]},
      {stage1_18[92]}
   );
   gpc1_1 gpc1668 (
      {stage0_18[249]},
      {stage1_18[93]}
   );
   gpc1_1 gpc1669 (
      {stage0_18[250]},
      {stage1_18[94]}
   );
   gpc1_1 gpc1670 (
      {stage0_18[251]},
      {stage1_18[95]}
   );
   gpc1_1 gpc1671 (
      {stage0_18[252]},
      {stage1_18[96]}
   );
   gpc1_1 gpc1672 (
      {stage0_18[253]},
      {stage1_18[97]}
   );
   gpc1_1 gpc1673 (
      {stage0_18[254]},
      {stage1_18[98]}
   );
   gpc1_1 gpc1674 (
      {stage0_18[255]},
      {stage1_18[99]}
   );
   gpc1_1 gpc1675 (
      {stage0_19[224]},
      {stage1_19[94]}
   );
   gpc1_1 gpc1676 (
      {stage0_19[225]},
      {stage1_19[95]}
   );
   gpc1_1 gpc1677 (
      {stage0_19[226]},
      {stage1_19[96]}
   );
   gpc1_1 gpc1678 (
      {stage0_19[227]},
      {stage1_19[97]}
   );
   gpc1_1 gpc1679 (
      {stage0_19[228]},
      {stage1_19[98]}
   );
   gpc1_1 gpc1680 (
      {stage0_19[229]},
      {stage1_19[99]}
   );
   gpc1_1 gpc1681 (
      {stage0_19[230]},
      {stage1_19[100]}
   );
   gpc1_1 gpc1682 (
      {stage0_19[231]},
      {stage1_19[101]}
   );
   gpc1_1 gpc1683 (
      {stage0_19[232]},
      {stage1_19[102]}
   );
   gpc1_1 gpc1684 (
      {stage0_19[233]},
      {stage1_19[103]}
   );
   gpc1_1 gpc1685 (
      {stage0_19[234]},
      {stage1_19[104]}
   );
   gpc1_1 gpc1686 (
      {stage0_19[235]},
      {stage1_19[105]}
   );
   gpc1_1 gpc1687 (
      {stage0_19[236]},
      {stage1_19[106]}
   );
   gpc1_1 gpc1688 (
      {stage0_19[237]},
      {stage1_19[107]}
   );
   gpc1_1 gpc1689 (
      {stage0_19[238]},
      {stage1_19[108]}
   );
   gpc1_1 gpc1690 (
      {stage0_19[239]},
      {stage1_19[109]}
   );
   gpc1_1 gpc1691 (
      {stage0_19[240]},
      {stage1_19[110]}
   );
   gpc1_1 gpc1692 (
      {stage0_19[241]},
      {stage1_19[111]}
   );
   gpc1_1 gpc1693 (
      {stage0_19[242]},
      {stage1_19[112]}
   );
   gpc1_1 gpc1694 (
      {stage0_19[243]},
      {stage1_19[113]}
   );
   gpc1_1 gpc1695 (
      {stage0_19[244]},
      {stage1_19[114]}
   );
   gpc1_1 gpc1696 (
      {stage0_19[245]},
      {stage1_19[115]}
   );
   gpc1_1 gpc1697 (
      {stage0_19[246]},
      {stage1_19[116]}
   );
   gpc1_1 gpc1698 (
      {stage0_19[247]},
      {stage1_19[117]}
   );
   gpc1_1 gpc1699 (
      {stage0_19[248]},
      {stage1_19[118]}
   );
   gpc1_1 gpc1700 (
      {stage0_19[249]},
      {stage1_19[119]}
   );
   gpc1_1 gpc1701 (
      {stage0_19[250]},
      {stage1_19[120]}
   );
   gpc1_1 gpc1702 (
      {stage0_19[251]},
      {stage1_19[121]}
   );
   gpc1_1 gpc1703 (
      {stage0_19[252]},
      {stage1_19[122]}
   );
   gpc1_1 gpc1704 (
      {stage0_19[253]},
      {stage1_19[123]}
   );
   gpc1_1 gpc1705 (
      {stage0_19[254]},
      {stage1_19[124]}
   );
   gpc1_1 gpc1706 (
      {stage0_19[255]},
      {stage1_19[125]}
   );
   gpc1_1 gpc1707 (
      {stage0_20[245]},
      {stage1_20[119]}
   );
   gpc1_1 gpc1708 (
      {stage0_20[246]},
      {stage1_20[120]}
   );
   gpc1_1 gpc1709 (
      {stage0_20[247]},
      {stage1_20[121]}
   );
   gpc1_1 gpc1710 (
      {stage0_20[248]},
      {stage1_20[122]}
   );
   gpc1_1 gpc1711 (
      {stage0_20[249]},
      {stage1_20[123]}
   );
   gpc1_1 gpc1712 (
      {stage0_20[250]},
      {stage1_20[124]}
   );
   gpc1_1 gpc1713 (
      {stage0_20[251]},
      {stage1_20[125]}
   );
   gpc1_1 gpc1714 (
      {stage0_20[252]},
      {stage1_20[126]}
   );
   gpc1_1 gpc1715 (
      {stage0_20[253]},
      {stage1_20[127]}
   );
   gpc1_1 gpc1716 (
      {stage0_20[254]},
      {stage1_20[128]}
   );
   gpc1_1 gpc1717 (
      {stage0_20[255]},
      {stage1_20[129]}
   );
   gpc1_1 gpc1718 (
      {stage0_21[252]},
      {stage1_21[104]}
   );
   gpc1_1 gpc1719 (
      {stage0_21[253]},
      {stage1_21[105]}
   );
   gpc1_1 gpc1720 (
      {stage0_21[254]},
      {stage1_21[106]}
   );
   gpc1_1 gpc1721 (
      {stage0_21[255]},
      {stage1_21[107]}
   );
   gpc1_1 gpc1722 (
      {stage0_22[252]},
      {stage1_22[88]}
   );
   gpc1_1 gpc1723 (
      {stage0_22[253]},
      {stage1_22[89]}
   );
   gpc1_1 gpc1724 (
      {stage0_22[254]},
      {stage1_22[90]}
   );
   gpc1_1 gpc1725 (
      {stage0_22[255]},
      {stage1_22[91]}
   );
   gpc1_1 gpc1726 (
      {stage0_23[226]},
      {stage1_23[99]}
   );
   gpc1_1 gpc1727 (
      {stage0_23[227]},
      {stage1_23[100]}
   );
   gpc1_1 gpc1728 (
      {stage0_23[228]},
      {stage1_23[101]}
   );
   gpc1_1 gpc1729 (
      {stage0_23[229]},
      {stage1_23[102]}
   );
   gpc1_1 gpc1730 (
      {stage0_23[230]},
      {stage1_23[103]}
   );
   gpc1_1 gpc1731 (
      {stage0_23[231]},
      {stage1_23[104]}
   );
   gpc1_1 gpc1732 (
      {stage0_23[232]},
      {stage1_23[105]}
   );
   gpc1_1 gpc1733 (
      {stage0_23[233]},
      {stage1_23[106]}
   );
   gpc1_1 gpc1734 (
      {stage0_23[234]},
      {stage1_23[107]}
   );
   gpc1_1 gpc1735 (
      {stage0_23[235]},
      {stage1_23[108]}
   );
   gpc1_1 gpc1736 (
      {stage0_23[236]},
      {stage1_23[109]}
   );
   gpc1_1 gpc1737 (
      {stage0_23[237]},
      {stage1_23[110]}
   );
   gpc1_1 gpc1738 (
      {stage0_23[238]},
      {stage1_23[111]}
   );
   gpc1_1 gpc1739 (
      {stage0_23[239]},
      {stage1_23[112]}
   );
   gpc1_1 gpc1740 (
      {stage0_23[240]},
      {stage1_23[113]}
   );
   gpc1_1 gpc1741 (
      {stage0_23[241]},
      {stage1_23[114]}
   );
   gpc1_1 gpc1742 (
      {stage0_23[242]},
      {stage1_23[115]}
   );
   gpc1_1 gpc1743 (
      {stage0_23[243]},
      {stage1_23[116]}
   );
   gpc1_1 gpc1744 (
      {stage0_23[244]},
      {stage1_23[117]}
   );
   gpc1_1 gpc1745 (
      {stage0_23[245]},
      {stage1_23[118]}
   );
   gpc1_1 gpc1746 (
      {stage0_23[246]},
      {stage1_23[119]}
   );
   gpc1_1 gpc1747 (
      {stage0_23[247]},
      {stage1_23[120]}
   );
   gpc1_1 gpc1748 (
      {stage0_23[248]},
      {stage1_23[121]}
   );
   gpc1_1 gpc1749 (
      {stage0_23[249]},
      {stage1_23[122]}
   );
   gpc1_1 gpc1750 (
      {stage0_23[250]},
      {stage1_23[123]}
   );
   gpc1_1 gpc1751 (
      {stage0_23[251]},
      {stage1_23[124]}
   );
   gpc1_1 gpc1752 (
      {stage0_23[252]},
      {stage1_23[125]}
   );
   gpc1_1 gpc1753 (
      {stage0_23[253]},
      {stage1_23[126]}
   );
   gpc1_1 gpc1754 (
      {stage0_23[254]},
      {stage1_23[127]}
   );
   gpc1_1 gpc1755 (
      {stage0_23[255]},
      {stage1_23[128]}
   );
   gpc1_1 gpc1756 (
      {stage0_24[231]},
      {stage1_24[115]}
   );
   gpc1_1 gpc1757 (
      {stage0_24[232]},
      {stage1_24[116]}
   );
   gpc1_1 gpc1758 (
      {stage0_24[233]},
      {stage1_24[117]}
   );
   gpc1_1 gpc1759 (
      {stage0_24[234]},
      {stage1_24[118]}
   );
   gpc1_1 gpc1760 (
      {stage0_24[235]},
      {stage1_24[119]}
   );
   gpc1_1 gpc1761 (
      {stage0_24[236]},
      {stage1_24[120]}
   );
   gpc1_1 gpc1762 (
      {stage0_24[237]},
      {stage1_24[121]}
   );
   gpc1_1 gpc1763 (
      {stage0_24[238]},
      {stage1_24[122]}
   );
   gpc1_1 gpc1764 (
      {stage0_24[239]},
      {stage1_24[123]}
   );
   gpc1_1 gpc1765 (
      {stage0_24[240]},
      {stage1_24[124]}
   );
   gpc1_1 gpc1766 (
      {stage0_24[241]},
      {stage1_24[125]}
   );
   gpc1_1 gpc1767 (
      {stage0_24[242]},
      {stage1_24[126]}
   );
   gpc1_1 gpc1768 (
      {stage0_24[243]},
      {stage1_24[127]}
   );
   gpc1_1 gpc1769 (
      {stage0_24[244]},
      {stage1_24[128]}
   );
   gpc1_1 gpc1770 (
      {stage0_24[245]},
      {stage1_24[129]}
   );
   gpc1_1 gpc1771 (
      {stage0_24[246]},
      {stage1_24[130]}
   );
   gpc1_1 gpc1772 (
      {stage0_24[247]},
      {stage1_24[131]}
   );
   gpc1_1 gpc1773 (
      {stage0_24[248]},
      {stage1_24[132]}
   );
   gpc1_1 gpc1774 (
      {stage0_24[249]},
      {stage1_24[133]}
   );
   gpc1_1 gpc1775 (
      {stage0_24[250]},
      {stage1_24[134]}
   );
   gpc1_1 gpc1776 (
      {stage0_24[251]},
      {stage1_24[135]}
   );
   gpc1_1 gpc1777 (
      {stage0_24[252]},
      {stage1_24[136]}
   );
   gpc1_1 gpc1778 (
      {stage0_24[253]},
      {stage1_24[137]}
   );
   gpc1_1 gpc1779 (
      {stage0_24[254]},
      {stage1_24[138]}
   );
   gpc1_1 gpc1780 (
      {stage0_24[255]},
      {stage1_24[139]}
   );
   gpc1_1 gpc1781 (
      {stage0_25[245]},
      {stage1_25[99]}
   );
   gpc1_1 gpc1782 (
      {stage0_25[246]},
      {stage1_25[100]}
   );
   gpc1_1 gpc1783 (
      {stage0_25[247]},
      {stage1_25[101]}
   );
   gpc1_1 gpc1784 (
      {stage0_25[248]},
      {stage1_25[102]}
   );
   gpc1_1 gpc1785 (
      {stage0_25[249]},
      {stage1_25[103]}
   );
   gpc1_1 gpc1786 (
      {stage0_25[250]},
      {stage1_25[104]}
   );
   gpc1_1 gpc1787 (
      {stage0_25[251]},
      {stage1_25[105]}
   );
   gpc1_1 gpc1788 (
      {stage0_25[252]},
      {stage1_25[106]}
   );
   gpc1_1 gpc1789 (
      {stage0_25[253]},
      {stage1_25[107]}
   );
   gpc1_1 gpc1790 (
      {stage0_25[254]},
      {stage1_25[108]}
   );
   gpc1_1 gpc1791 (
      {stage0_25[255]},
      {stage1_25[109]}
   );
   gpc1_1 gpc1792 (
      {stage0_26[195]},
      {stage1_26[80]}
   );
   gpc1_1 gpc1793 (
      {stage0_26[196]},
      {stage1_26[81]}
   );
   gpc1_1 gpc1794 (
      {stage0_26[197]},
      {stage1_26[82]}
   );
   gpc1_1 gpc1795 (
      {stage0_26[198]},
      {stage1_26[83]}
   );
   gpc1_1 gpc1796 (
      {stage0_26[199]},
      {stage1_26[84]}
   );
   gpc1_1 gpc1797 (
      {stage0_26[200]},
      {stage1_26[85]}
   );
   gpc1_1 gpc1798 (
      {stage0_26[201]},
      {stage1_26[86]}
   );
   gpc1_1 gpc1799 (
      {stage0_26[202]},
      {stage1_26[87]}
   );
   gpc1_1 gpc1800 (
      {stage0_26[203]},
      {stage1_26[88]}
   );
   gpc1_1 gpc1801 (
      {stage0_26[204]},
      {stage1_26[89]}
   );
   gpc1_1 gpc1802 (
      {stage0_26[205]},
      {stage1_26[90]}
   );
   gpc1_1 gpc1803 (
      {stage0_26[206]},
      {stage1_26[91]}
   );
   gpc1_1 gpc1804 (
      {stage0_26[207]},
      {stage1_26[92]}
   );
   gpc1_1 gpc1805 (
      {stage0_26[208]},
      {stage1_26[93]}
   );
   gpc1_1 gpc1806 (
      {stage0_26[209]},
      {stage1_26[94]}
   );
   gpc1_1 gpc1807 (
      {stage0_26[210]},
      {stage1_26[95]}
   );
   gpc1_1 gpc1808 (
      {stage0_26[211]},
      {stage1_26[96]}
   );
   gpc1_1 gpc1809 (
      {stage0_26[212]},
      {stage1_26[97]}
   );
   gpc1_1 gpc1810 (
      {stage0_26[213]},
      {stage1_26[98]}
   );
   gpc1_1 gpc1811 (
      {stage0_26[214]},
      {stage1_26[99]}
   );
   gpc1_1 gpc1812 (
      {stage0_26[215]},
      {stage1_26[100]}
   );
   gpc1_1 gpc1813 (
      {stage0_26[216]},
      {stage1_26[101]}
   );
   gpc1_1 gpc1814 (
      {stage0_26[217]},
      {stage1_26[102]}
   );
   gpc1_1 gpc1815 (
      {stage0_26[218]},
      {stage1_26[103]}
   );
   gpc1_1 gpc1816 (
      {stage0_26[219]},
      {stage1_26[104]}
   );
   gpc1_1 gpc1817 (
      {stage0_26[220]},
      {stage1_26[105]}
   );
   gpc1_1 gpc1818 (
      {stage0_26[221]},
      {stage1_26[106]}
   );
   gpc1_1 gpc1819 (
      {stage0_26[222]},
      {stage1_26[107]}
   );
   gpc1_1 gpc1820 (
      {stage0_26[223]},
      {stage1_26[108]}
   );
   gpc1_1 gpc1821 (
      {stage0_26[224]},
      {stage1_26[109]}
   );
   gpc1_1 gpc1822 (
      {stage0_26[225]},
      {stage1_26[110]}
   );
   gpc1_1 gpc1823 (
      {stage0_26[226]},
      {stage1_26[111]}
   );
   gpc1_1 gpc1824 (
      {stage0_26[227]},
      {stage1_26[112]}
   );
   gpc1_1 gpc1825 (
      {stage0_26[228]},
      {stage1_26[113]}
   );
   gpc1_1 gpc1826 (
      {stage0_26[229]},
      {stage1_26[114]}
   );
   gpc1_1 gpc1827 (
      {stage0_26[230]},
      {stage1_26[115]}
   );
   gpc1_1 gpc1828 (
      {stage0_26[231]},
      {stage1_26[116]}
   );
   gpc1_1 gpc1829 (
      {stage0_26[232]},
      {stage1_26[117]}
   );
   gpc1_1 gpc1830 (
      {stage0_26[233]},
      {stage1_26[118]}
   );
   gpc1_1 gpc1831 (
      {stage0_26[234]},
      {stage1_26[119]}
   );
   gpc1_1 gpc1832 (
      {stage0_26[235]},
      {stage1_26[120]}
   );
   gpc1_1 gpc1833 (
      {stage0_26[236]},
      {stage1_26[121]}
   );
   gpc1_1 gpc1834 (
      {stage0_26[237]},
      {stage1_26[122]}
   );
   gpc1_1 gpc1835 (
      {stage0_26[238]},
      {stage1_26[123]}
   );
   gpc1_1 gpc1836 (
      {stage0_26[239]},
      {stage1_26[124]}
   );
   gpc1_1 gpc1837 (
      {stage0_26[240]},
      {stage1_26[125]}
   );
   gpc1_1 gpc1838 (
      {stage0_26[241]},
      {stage1_26[126]}
   );
   gpc1_1 gpc1839 (
      {stage0_26[242]},
      {stage1_26[127]}
   );
   gpc1_1 gpc1840 (
      {stage0_26[243]},
      {stage1_26[128]}
   );
   gpc1_1 gpc1841 (
      {stage0_26[244]},
      {stage1_26[129]}
   );
   gpc1_1 gpc1842 (
      {stage0_26[245]},
      {stage1_26[130]}
   );
   gpc1_1 gpc1843 (
      {stage0_26[246]},
      {stage1_26[131]}
   );
   gpc1_1 gpc1844 (
      {stage0_26[247]},
      {stage1_26[132]}
   );
   gpc1_1 gpc1845 (
      {stage0_26[248]},
      {stage1_26[133]}
   );
   gpc1_1 gpc1846 (
      {stage0_26[249]},
      {stage1_26[134]}
   );
   gpc1_1 gpc1847 (
      {stage0_26[250]},
      {stage1_26[135]}
   );
   gpc1_1 gpc1848 (
      {stage0_26[251]},
      {stage1_26[136]}
   );
   gpc1_1 gpc1849 (
      {stage0_26[252]},
      {stage1_26[137]}
   );
   gpc1_1 gpc1850 (
      {stage0_26[253]},
      {stage1_26[138]}
   );
   gpc1_1 gpc1851 (
      {stage0_26[254]},
      {stage1_26[139]}
   );
   gpc1_1 gpc1852 (
      {stage0_26[255]},
      {stage1_26[140]}
   );
   gpc1_1 gpc1853 (
      {stage0_27[224]},
      {stage1_27[87]}
   );
   gpc1_1 gpc1854 (
      {stage0_27[225]},
      {stage1_27[88]}
   );
   gpc1_1 gpc1855 (
      {stage0_27[226]},
      {stage1_27[89]}
   );
   gpc1_1 gpc1856 (
      {stage0_27[227]},
      {stage1_27[90]}
   );
   gpc1_1 gpc1857 (
      {stage0_27[228]},
      {stage1_27[91]}
   );
   gpc1_1 gpc1858 (
      {stage0_27[229]},
      {stage1_27[92]}
   );
   gpc1_1 gpc1859 (
      {stage0_27[230]},
      {stage1_27[93]}
   );
   gpc1_1 gpc1860 (
      {stage0_27[231]},
      {stage1_27[94]}
   );
   gpc1_1 gpc1861 (
      {stage0_27[232]},
      {stage1_27[95]}
   );
   gpc1_1 gpc1862 (
      {stage0_27[233]},
      {stage1_27[96]}
   );
   gpc1_1 gpc1863 (
      {stage0_27[234]},
      {stage1_27[97]}
   );
   gpc1_1 gpc1864 (
      {stage0_27[235]},
      {stage1_27[98]}
   );
   gpc1_1 gpc1865 (
      {stage0_27[236]},
      {stage1_27[99]}
   );
   gpc1_1 gpc1866 (
      {stage0_27[237]},
      {stage1_27[100]}
   );
   gpc1_1 gpc1867 (
      {stage0_27[238]},
      {stage1_27[101]}
   );
   gpc1_1 gpc1868 (
      {stage0_27[239]},
      {stage1_27[102]}
   );
   gpc1_1 gpc1869 (
      {stage0_27[240]},
      {stage1_27[103]}
   );
   gpc1_1 gpc1870 (
      {stage0_27[241]},
      {stage1_27[104]}
   );
   gpc1_1 gpc1871 (
      {stage0_27[242]},
      {stage1_27[105]}
   );
   gpc1_1 gpc1872 (
      {stage0_27[243]},
      {stage1_27[106]}
   );
   gpc1_1 gpc1873 (
      {stage0_27[244]},
      {stage1_27[107]}
   );
   gpc1_1 gpc1874 (
      {stage0_27[245]},
      {stage1_27[108]}
   );
   gpc1_1 gpc1875 (
      {stage0_27[246]},
      {stage1_27[109]}
   );
   gpc1_1 gpc1876 (
      {stage0_27[247]},
      {stage1_27[110]}
   );
   gpc1_1 gpc1877 (
      {stage0_27[248]},
      {stage1_27[111]}
   );
   gpc1_1 gpc1878 (
      {stage0_27[249]},
      {stage1_27[112]}
   );
   gpc1_1 gpc1879 (
      {stage0_27[250]},
      {stage1_27[113]}
   );
   gpc1_1 gpc1880 (
      {stage0_27[251]},
      {stage1_27[114]}
   );
   gpc1_1 gpc1881 (
      {stage0_27[252]},
      {stage1_27[115]}
   );
   gpc1_1 gpc1882 (
      {stage0_27[253]},
      {stage1_27[116]}
   );
   gpc1_1 gpc1883 (
      {stage0_27[254]},
      {stage1_27[117]}
   );
   gpc1_1 gpc1884 (
      {stage0_27[255]},
      {stage1_27[118]}
   );
   gpc1_1 gpc1885 (
      {stage0_28[235]},
      {stage1_28[106]}
   );
   gpc1_1 gpc1886 (
      {stage0_28[236]},
      {stage1_28[107]}
   );
   gpc1_1 gpc1887 (
      {stage0_28[237]},
      {stage1_28[108]}
   );
   gpc1_1 gpc1888 (
      {stage0_28[238]},
      {stage1_28[109]}
   );
   gpc1_1 gpc1889 (
      {stage0_28[239]},
      {stage1_28[110]}
   );
   gpc1_1 gpc1890 (
      {stage0_28[240]},
      {stage1_28[111]}
   );
   gpc1_1 gpc1891 (
      {stage0_28[241]},
      {stage1_28[112]}
   );
   gpc1_1 gpc1892 (
      {stage0_28[242]},
      {stage1_28[113]}
   );
   gpc1_1 gpc1893 (
      {stage0_28[243]},
      {stage1_28[114]}
   );
   gpc1_1 gpc1894 (
      {stage0_28[244]},
      {stage1_28[115]}
   );
   gpc1_1 gpc1895 (
      {stage0_28[245]},
      {stage1_28[116]}
   );
   gpc1_1 gpc1896 (
      {stage0_28[246]},
      {stage1_28[117]}
   );
   gpc1_1 gpc1897 (
      {stage0_28[247]},
      {stage1_28[118]}
   );
   gpc1_1 gpc1898 (
      {stage0_28[248]},
      {stage1_28[119]}
   );
   gpc1_1 gpc1899 (
      {stage0_28[249]},
      {stage1_28[120]}
   );
   gpc1_1 gpc1900 (
      {stage0_28[250]},
      {stage1_28[121]}
   );
   gpc1_1 gpc1901 (
      {stage0_28[251]},
      {stage1_28[122]}
   );
   gpc1_1 gpc1902 (
      {stage0_28[252]},
      {stage1_28[123]}
   );
   gpc1_1 gpc1903 (
      {stage0_28[253]},
      {stage1_28[124]}
   );
   gpc1_1 gpc1904 (
      {stage0_28[254]},
      {stage1_28[125]}
   );
   gpc1_1 gpc1905 (
      {stage0_28[255]},
      {stage1_28[126]}
   );
   gpc1_1 gpc1906 (
      {stage0_29[247]},
      {stage1_29[101]}
   );
   gpc1_1 gpc1907 (
      {stage0_29[248]},
      {stage1_29[102]}
   );
   gpc1_1 gpc1908 (
      {stage0_29[249]},
      {stage1_29[103]}
   );
   gpc1_1 gpc1909 (
      {stage0_29[250]},
      {stage1_29[104]}
   );
   gpc1_1 gpc1910 (
      {stage0_29[251]},
      {stage1_29[105]}
   );
   gpc1_1 gpc1911 (
      {stage0_29[252]},
      {stage1_29[106]}
   );
   gpc1_1 gpc1912 (
      {stage0_29[253]},
      {stage1_29[107]}
   );
   gpc1_1 gpc1913 (
      {stage0_29[254]},
      {stage1_29[108]}
   );
   gpc1_1 gpc1914 (
      {stage0_29[255]},
      {stage1_29[109]}
   );
   gpc1_1 gpc1915 (
      {stage0_30[254]},
      {stage1_30[89]}
   );
   gpc1_1 gpc1916 (
      {stage0_30[255]},
      {stage1_30[90]}
   );
   gpc1_1 gpc1917 (
      {stage0_31[243]},
      {stage1_31[102]}
   );
   gpc1_1 gpc1918 (
      {stage0_31[244]},
      {stage1_31[103]}
   );
   gpc1_1 gpc1919 (
      {stage0_31[245]},
      {stage1_31[104]}
   );
   gpc1_1 gpc1920 (
      {stage0_31[246]},
      {stage1_31[105]}
   );
   gpc1_1 gpc1921 (
      {stage0_31[247]},
      {stage1_31[106]}
   );
   gpc1_1 gpc1922 (
      {stage0_31[248]},
      {stage1_31[107]}
   );
   gpc1_1 gpc1923 (
      {stage0_31[249]},
      {stage1_31[108]}
   );
   gpc1_1 gpc1924 (
      {stage0_31[250]},
      {stage1_31[109]}
   );
   gpc1_1 gpc1925 (
      {stage0_31[251]},
      {stage1_31[110]}
   );
   gpc1_1 gpc1926 (
      {stage0_31[252]},
      {stage1_31[111]}
   );
   gpc1_1 gpc1927 (
      {stage0_31[253]},
      {stage1_31[112]}
   );
   gpc1_1 gpc1928 (
      {stage0_31[254]},
      {stage1_31[113]}
   );
   gpc1_1 gpc1929 (
      {stage0_31[255]},
      {stage1_31[114]}
   );
   gpc1_1 gpc1930 (
      {stage0_33[252]},
      {stage1_33[107]}
   );
   gpc1_1 gpc1931 (
      {stage0_33[253]},
      {stage1_33[108]}
   );
   gpc1_1 gpc1932 (
      {stage0_33[254]},
      {stage1_33[109]}
   );
   gpc1_1 gpc1933 (
      {stage0_33[255]},
      {stage1_33[110]}
   );
   gpc1_1 gpc1934 (
      {stage0_34[249]},
      {stage1_34[97]}
   );
   gpc1_1 gpc1935 (
      {stage0_34[250]},
      {stage1_34[98]}
   );
   gpc1_1 gpc1936 (
      {stage0_34[251]},
      {stage1_34[99]}
   );
   gpc1_1 gpc1937 (
      {stage0_34[252]},
      {stage1_34[100]}
   );
   gpc1_1 gpc1938 (
      {stage0_34[253]},
      {stage1_34[101]}
   );
   gpc1_1 gpc1939 (
      {stage0_34[254]},
      {stage1_34[102]}
   );
   gpc1_1 gpc1940 (
      {stage0_34[255]},
      {stage1_34[103]}
   );
   gpc1_1 gpc1941 (
      {stage0_35[236]},
      {stage1_35[99]}
   );
   gpc1_1 gpc1942 (
      {stage0_35[237]},
      {stage1_35[100]}
   );
   gpc1_1 gpc1943 (
      {stage0_35[238]},
      {stage1_35[101]}
   );
   gpc1_1 gpc1944 (
      {stage0_35[239]},
      {stage1_35[102]}
   );
   gpc1_1 gpc1945 (
      {stage0_35[240]},
      {stage1_35[103]}
   );
   gpc1_1 gpc1946 (
      {stage0_35[241]},
      {stage1_35[104]}
   );
   gpc1_1 gpc1947 (
      {stage0_35[242]},
      {stage1_35[105]}
   );
   gpc1_1 gpc1948 (
      {stage0_35[243]},
      {stage1_35[106]}
   );
   gpc1_1 gpc1949 (
      {stage0_35[244]},
      {stage1_35[107]}
   );
   gpc1_1 gpc1950 (
      {stage0_35[245]},
      {stage1_35[108]}
   );
   gpc1_1 gpc1951 (
      {stage0_35[246]},
      {stage1_35[109]}
   );
   gpc1_1 gpc1952 (
      {stage0_35[247]},
      {stage1_35[110]}
   );
   gpc1_1 gpc1953 (
      {stage0_35[248]},
      {stage1_35[111]}
   );
   gpc1_1 gpc1954 (
      {stage0_35[249]},
      {stage1_35[112]}
   );
   gpc1_1 gpc1955 (
      {stage0_35[250]},
      {stage1_35[113]}
   );
   gpc1_1 gpc1956 (
      {stage0_35[251]},
      {stage1_35[114]}
   );
   gpc1_1 gpc1957 (
      {stage0_35[252]},
      {stage1_35[115]}
   );
   gpc1_1 gpc1958 (
      {stage0_35[253]},
      {stage1_35[116]}
   );
   gpc1_1 gpc1959 (
      {stage0_35[254]},
      {stage1_35[117]}
   );
   gpc1_1 gpc1960 (
      {stage0_35[255]},
      {stage1_35[118]}
   );
   gpc1_1 gpc1961 (
      {stage0_36[212]},
      {stage1_36[101]}
   );
   gpc1_1 gpc1962 (
      {stage0_36[213]},
      {stage1_36[102]}
   );
   gpc1_1 gpc1963 (
      {stage0_36[214]},
      {stage1_36[103]}
   );
   gpc1_1 gpc1964 (
      {stage0_36[215]},
      {stage1_36[104]}
   );
   gpc1_1 gpc1965 (
      {stage0_36[216]},
      {stage1_36[105]}
   );
   gpc1_1 gpc1966 (
      {stage0_36[217]},
      {stage1_36[106]}
   );
   gpc1_1 gpc1967 (
      {stage0_36[218]},
      {stage1_36[107]}
   );
   gpc1_1 gpc1968 (
      {stage0_36[219]},
      {stage1_36[108]}
   );
   gpc1_1 gpc1969 (
      {stage0_36[220]},
      {stage1_36[109]}
   );
   gpc1_1 gpc1970 (
      {stage0_36[221]},
      {stage1_36[110]}
   );
   gpc1_1 gpc1971 (
      {stage0_36[222]},
      {stage1_36[111]}
   );
   gpc1_1 gpc1972 (
      {stage0_36[223]},
      {stage1_36[112]}
   );
   gpc1_1 gpc1973 (
      {stage0_36[224]},
      {stage1_36[113]}
   );
   gpc1_1 gpc1974 (
      {stage0_36[225]},
      {stage1_36[114]}
   );
   gpc1_1 gpc1975 (
      {stage0_36[226]},
      {stage1_36[115]}
   );
   gpc1_1 gpc1976 (
      {stage0_36[227]},
      {stage1_36[116]}
   );
   gpc1_1 gpc1977 (
      {stage0_36[228]},
      {stage1_36[117]}
   );
   gpc1_1 gpc1978 (
      {stage0_36[229]},
      {stage1_36[118]}
   );
   gpc1_1 gpc1979 (
      {stage0_36[230]},
      {stage1_36[119]}
   );
   gpc1_1 gpc1980 (
      {stage0_36[231]},
      {stage1_36[120]}
   );
   gpc1_1 gpc1981 (
      {stage0_36[232]},
      {stage1_36[121]}
   );
   gpc1_1 gpc1982 (
      {stage0_36[233]},
      {stage1_36[122]}
   );
   gpc1_1 gpc1983 (
      {stage0_36[234]},
      {stage1_36[123]}
   );
   gpc1_1 gpc1984 (
      {stage0_36[235]},
      {stage1_36[124]}
   );
   gpc1_1 gpc1985 (
      {stage0_36[236]},
      {stage1_36[125]}
   );
   gpc1_1 gpc1986 (
      {stage0_36[237]},
      {stage1_36[126]}
   );
   gpc1_1 gpc1987 (
      {stage0_36[238]},
      {stage1_36[127]}
   );
   gpc1_1 gpc1988 (
      {stage0_36[239]},
      {stage1_36[128]}
   );
   gpc1_1 gpc1989 (
      {stage0_36[240]},
      {stage1_36[129]}
   );
   gpc1_1 gpc1990 (
      {stage0_36[241]},
      {stage1_36[130]}
   );
   gpc1_1 gpc1991 (
      {stage0_36[242]},
      {stage1_36[131]}
   );
   gpc1_1 gpc1992 (
      {stage0_36[243]},
      {stage1_36[132]}
   );
   gpc1_1 gpc1993 (
      {stage0_36[244]},
      {stage1_36[133]}
   );
   gpc1_1 gpc1994 (
      {stage0_36[245]},
      {stage1_36[134]}
   );
   gpc1_1 gpc1995 (
      {stage0_36[246]},
      {stage1_36[135]}
   );
   gpc1_1 gpc1996 (
      {stage0_36[247]},
      {stage1_36[136]}
   );
   gpc1_1 gpc1997 (
      {stage0_36[248]},
      {stage1_36[137]}
   );
   gpc1_1 gpc1998 (
      {stage0_36[249]},
      {stage1_36[138]}
   );
   gpc1_1 gpc1999 (
      {stage0_36[250]},
      {stage1_36[139]}
   );
   gpc1_1 gpc2000 (
      {stage0_36[251]},
      {stage1_36[140]}
   );
   gpc1_1 gpc2001 (
      {stage0_36[252]},
      {stage1_36[141]}
   );
   gpc1_1 gpc2002 (
      {stage0_36[253]},
      {stage1_36[142]}
   );
   gpc1_1 gpc2003 (
      {stage0_36[254]},
      {stage1_36[143]}
   );
   gpc1_1 gpc2004 (
      {stage0_36[255]},
      {stage1_36[144]}
   );
   gpc1_1 gpc2005 (
      {stage0_37[252]},
      {stage1_37[101]}
   );
   gpc1_1 gpc2006 (
      {stage0_37[253]},
      {stage1_37[102]}
   );
   gpc1_1 gpc2007 (
      {stage0_37[254]},
      {stage1_37[103]}
   );
   gpc1_1 gpc2008 (
      {stage0_37[255]},
      {stage1_37[104]}
   );
   gpc1_1 gpc2009 (
      {stage0_38[217]},
      {stage1_38[98]}
   );
   gpc1_1 gpc2010 (
      {stage0_38[218]},
      {stage1_38[99]}
   );
   gpc1_1 gpc2011 (
      {stage0_38[219]},
      {stage1_38[100]}
   );
   gpc1_1 gpc2012 (
      {stage0_38[220]},
      {stage1_38[101]}
   );
   gpc1_1 gpc2013 (
      {stage0_38[221]},
      {stage1_38[102]}
   );
   gpc1_1 gpc2014 (
      {stage0_38[222]},
      {stage1_38[103]}
   );
   gpc1_1 gpc2015 (
      {stage0_38[223]},
      {stage1_38[104]}
   );
   gpc1_1 gpc2016 (
      {stage0_38[224]},
      {stage1_38[105]}
   );
   gpc1_1 gpc2017 (
      {stage0_38[225]},
      {stage1_38[106]}
   );
   gpc1_1 gpc2018 (
      {stage0_38[226]},
      {stage1_38[107]}
   );
   gpc1_1 gpc2019 (
      {stage0_38[227]},
      {stage1_38[108]}
   );
   gpc1_1 gpc2020 (
      {stage0_38[228]},
      {stage1_38[109]}
   );
   gpc1_1 gpc2021 (
      {stage0_38[229]},
      {stage1_38[110]}
   );
   gpc1_1 gpc2022 (
      {stage0_38[230]},
      {stage1_38[111]}
   );
   gpc1_1 gpc2023 (
      {stage0_38[231]},
      {stage1_38[112]}
   );
   gpc1_1 gpc2024 (
      {stage0_38[232]},
      {stage1_38[113]}
   );
   gpc1_1 gpc2025 (
      {stage0_38[233]},
      {stage1_38[114]}
   );
   gpc1_1 gpc2026 (
      {stage0_38[234]},
      {stage1_38[115]}
   );
   gpc1_1 gpc2027 (
      {stage0_38[235]},
      {stage1_38[116]}
   );
   gpc1_1 gpc2028 (
      {stage0_38[236]},
      {stage1_38[117]}
   );
   gpc1_1 gpc2029 (
      {stage0_38[237]},
      {stage1_38[118]}
   );
   gpc1_1 gpc2030 (
      {stage0_38[238]},
      {stage1_38[119]}
   );
   gpc1_1 gpc2031 (
      {stage0_38[239]},
      {stage1_38[120]}
   );
   gpc1_1 gpc2032 (
      {stage0_38[240]},
      {stage1_38[121]}
   );
   gpc1_1 gpc2033 (
      {stage0_38[241]},
      {stage1_38[122]}
   );
   gpc1_1 gpc2034 (
      {stage0_38[242]},
      {stage1_38[123]}
   );
   gpc1_1 gpc2035 (
      {stage0_38[243]},
      {stage1_38[124]}
   );
   gpc1_1 gpc2036 (
      {stage0_38[244]},
      {stage1_38[125]}
   );
   gpc1_1 gpc2037 (
      {stage0_38[245]},
      {stage1_38[126]}
   );
   gpc1_1 gpc2038 (
      {stage0_38[246]},
      {stage1_38[127]}
   );
   gpc1_1 gpc2039 (
      {stage0_38[247]},
      {stage1_38[128]}
   );
   gpc1_1 gpc2040 (
      {stage0_38[248]},
      {stage1_38[129]}
   );
   gpc1_1 gpc2041 (
      {stage0_38[249]},
      {stage1_38[130]}
   );
   gpc1_1 gpc2042 (
      {stage0_38[250]},
      {stage1_38[131]}
   );
   gpc1_1 gpc2043 (
      {stage0_38[251]},
      {stage1_38[132]}
   );
   gpc1_1 gpc2044 (
      {stage0_38[252]},
      {stage1_38[133]}
   );
   gpc1_1 gpc2045 (
      {stage0_38[253]},
      {stage1_38[134]}
   );
   gpc1_1 gpc2046 (
      {stage0_38[254]},
      {stage1_38[135]}
   );
   gpc1_1 gpc2047 (
      {stage0_38[255]},
      {stage1_38[136]}
   );
   gpc1_1 gpc2048 (
      {stage0_39[218]},
      {stage1_39[87]}
   );
   gpc1_1 gpc2049 (
      {stage0_39[219]},
      {stage1_39[88]}
   );
   gpc1_1 gpc2050 (
      {stage0_39[220]},
      {stage1_39[89]}
   );
   gpc1_1 gpc2051 (
      {stage0_39[221]},
      {stage1_39[90]}
   );
   gpc1_1 gpc2052 (
      {stage0_39[222]},
      {stage1_39[91]}
   );
   gpc1_1 gpc2053 (
      {stage0_39[223]},
      {stage1_39[92]}
   );
   gpc1_1 gpc2054 (
      {stage0_39[224]},
      {stage1_39[93]}
   );
   gpc1_1 gpc2055 (
      {stage0_39[225]},
      {stage1_39[94]}
   );
   gpc1_1 gpc2056 (
      {stage0_39[226]},
      {stage1_39[95]}
   );
   gpc1_1 gpc2057 (
      {stage0_39[227]},
      {stage1_39[96]}
   );
   gpc1_1 gpc2058 (
      {stage0_39[228]},
      {stage1_39[97]}
   );
   gpc1_1 gpc2059 (
      {stage0_39[229]},
      {stage1_39[98]}
   );
   gpc1_1 gpc2060 (
      {stage0_39[230]},
      {stage1_39[99]}
   );
   gpc1_1 gpc2061 (
      {stage0_39[231]},
      {stage1_39[100]}
   );
   gpc1_1 gpc2062 (
      {stage0_39[232]},
      {stage1_39[101]}
   );
   gpc1_1 gpc2063 (
      {stage0_39[233]},
      {stage1_39[102]}
   );
   gpc1_1 gpc2064 (
      {stage0_39[234]},
      {stage1_39[103]}
   );
   gpc1_1 gpc2065 (
      {stage0_39[235]},
      {stage1_39[104]}
   );
   gpc1_1 gpc2066 (
      {stage0_39[236]},
      {stage1_39[105]}
   );
   gpc1_1 gpc2067 (
      {stage0_39[237]},
      {stage1_39[106]}
   );
   gpc1_1 gpc2068 (
      {stage0_39[238]},
      {stage1_39[107]}
   );
   gpc1_1 gpc2069 (
      {stage0_39[239]},
      {stage1_39[108]}
   );
   gpc1_1 gpc2070 (
      {stage0_39[240]},
      {stage1_39[109]}
   );
   gpc1_1 gpc2071 (
      {stage0_39[241]},
      {stage1_39[110]}
   );
   gpc1_1 gpc2072 (
      {stage0_39[242]},
      {stage1_39[111]}
   );
   gpc1_1 gpc2073 (
      {stage0_39[243]},
      {stage1_39[112]}
   );
   gpc1_1 gpc2074 (
      {stage0_39[244]},
      {stage1_39[113]}
   );
   gpc1_1 gpc2075 (
      {stage0_39[245]},
      {stage1_39[114]}
   );
   gpc1_1 gpc2076 (
      {stage0_39[246]},
      {stage1_39[115]}
   );
   gpc1_1 gpc2077 (
      {stage0_39[247]},
      {stage1_39[116]}
   );
   gpc1_1 gpc2078 (
      {stage0_39[248]},
      {stage1_39[117]}
   );
   gpc1_1 gpc2079 (
      {stage0_39[249]},
      {stage1_39[118]}
   );
   gpc1_1 gpc2080 (
      {stage0_39[250]},
      {stage1_39[119]}
   );
   gpc1_1 gpc2081 (
      {stage0_39[251]},
      {stage1_39[120]}
   );
   gpc1_1 gpc2082 (
      {stage0_39[252]},
      {stage1_39[121]}
   );
   gpc1_1 gpc2083 (
      {stage0_39[253]},
      {stage1_39[122]}
   );
   gpc1_1 gpc2084 (
      {stage0_39[254]},
      {stage1_39[123]}
   );
   gpc1_1 gpc2085 (
      {stage0_39[255]},
      {stage1_39[124]}
   );
   gpc1_1 gpc2086 (
      {stage0_41[224]},
      {stage1_41[111]}
   );
   gpc1_1 gpc2087 (
      {stage0_41[225]},
      {stage1_41[112]}
   );
   gpc1_1 gpc2088 (
      {stage0_41[226]},
      {stage1_41[113]}
   );
   gpc1_1 gpc2089 (
      {stage0_41[227]},
      {stage1_41[114]}
   );
   gpc1_1 gpc2090 (
      {stage0_41[228]},
      {stage1_41[115]}
   );
   gpc1_1 gpc2091 (
      {stage0_41[229]},
      {stage1_41[116]}
   );
   gpc1_1 gpc2092 (
      {stage0_41[230]},
      {stage1_41[117]}
   );
   gpc1_1 gpc2093 (
      {stage0_41[231]},
      {stage1_41[118]}
   );
   gpc1_1 gpc2094 (
      {stage0_41[232]},
      {stage1_41[119]}
   );
   gpc1_1 gpc2095 (
      {stage0_41[233]},
      {stage1_41[120]}
   );
   gpc1_1 gpc2096 (
      {stage0_41[234]},
      {stage1_41[121]}
   );
   gpc1_1 gpc2097 (
      {stage0_41[235]},
      {stage1_41[122]}
   );
   gpc1_1 gpc2098 (
      {stage0_41[236]},
      {stage1_41[123]}
   );
   gpc1_1 gpc2099 (
      {stage0_41[237]},
      {stage1_41[124]}
   );
   gpc1_1 gpc2100 (
      {stage0_41[238]},
      {stage1_41[125]}
   );
   gpc1_1 gpc2101 (
      {stage0_41[239]},
      {stage1_41[126]}
   );
   gpc1_1 gpc2102 (
      {stage0_41[240]},
      {stage1_41[127]}
   );
   gpc1_1 gpc2103 (
      {stage0_41[241]},
      {stage1_41[128]}
   );
   gpc1_1 gpc2104 (
      {stage0_41[242]},
      {stage1_41[129]}
   );
   gpc1_1 gpc2105 (
      {stage0_41[243]},
      {stage1_41[130]}
   );
   gpc1_1 gpc2106 (
      {stage0_41[244]},
      {stage1_41[131]}
   );
   gpc1_1 gpc2107 (
      {stage0_41[245]},
      {stage1_41[132]}
   );
   gpc1_1 gpc2108 (
      {stage0_41[246]},
      {stage1_41[133]}
   );
   gpc1_1 gpc2109 (
      {stage0_41[247]},
      {stage1_41[134]}
   );
   gpc1_1 gpc2110 (
      {stage0_41[248]},
      {stage1_41[135]}
   );
   gpc1_1 gpc2111 (
      {stage0_41[249]},
      {stage1_41[136]}
   );
   gpc1_1 gpc2112 (
      {stage0_41[250]},
      {stage1_41[137]}
   );
   gpc1_1 gpc2113 (
      {stage0_41[251]},
      {stage1_41[138]}
   );
   gpc1_1 gpc2114 (
      {stage0_41[252]},
      {stage1_41[139]}
   );
   gpc1_1 gpc2115 (
      {stage0_41[253]},
      {stage1_41[140]}
   );
   gpc1_1 gpc2116 (
      {stage0_41[254]},
      {stage1_41[141]}
   );
   gpc1_1 gpc2117 (
      {stage0_41[255]},
      {stage1_41[142]}
   );
   gpc1_1 gpc2118 (
      {stage0_42[175]},
      {stage1_42[91]}
   );
   gpc1_1 gpc2119 (
      {stage0_42[176]},
      {stage1_42[92]}
   );
   gpc1_1 gpc2120 (
      {stage0_42[177]},
      {stage1_42[93]}
   );
   gpc1_1 gpc2121 (
      {stage0_42[178]},
      {stage1_42[94]}
   );
   gpc1_1 gpc2122 (
      {stage0_42[179]},
      {stage1_42[95]}
   );
   gpc1_1 gpc2123 (
      {stage0_42[180]},
      {stage1_42[96]}
   );
   gpc1_1 gpc2124 (
      {stage0_42[181]},
      {stage1_42[97]}
   );
   gpc1_1 gpc2125 (
      {stage0_42[182]},
      {stage1_42[98]}
   );
   gpc1_1 gpc2126 (
      {stage0_42[183]},
      {stage1_42[99]}
   );
   gpc1_1 gpc2127 (
      {stage0_42[184]},
      {stage1_42[100]}
   );
   gpc1_1 gpc2128 (
      {stage0_42[185]},
      {stage1_42[101]}
   );
   gpc1_1 gpc2129 (
      {stage0_42[186]},
      {stage1_42[102]}
   );
   gpc1_1 gpc2130 (
      {stage0_42[187]},
      {stage1_42[103]}
   );
   gpc1_1 gpc2131 (
      {stage0_42[188]},
      {stage1_42[104]}
   );
   gpc1_1 gpc2132 (
      {stage0_42[189]},
      {stage1_42[105]}
   );
   gpc1_1 gpc2133 (
      {stage0_42[190]},
      {stage1_42[106]}
   );
   gpc1_1 gpc2134 (
      {stage0_42[191]},
      {stage1_42[107]}
   );
   gpc1_1 gpc2135 (
      {stage0_42[192]},
      {stage1_42[108]}
   );
   gpc1_1 gpc2136 (
      {stage0_42[193]},
      {stage1_42[109]}
   );
   gpc1_1 gpc2137 (
      {stage0_42[194]},
      {stage1_42[110]}
   );
   gpc1_1 gpc2138 (
      {stage0_42[195]},
      {stage1_42[111]}
   );
   gpc1_1 gpc2139 (
      {stage0_42[196]},
      {stage1_42[112]}
   );
   gpc1_1 gpc2140 (
      {stage0_42[197]},
      {stage1_42[113]}
   );
   gpc1_1 gpc2141 (
      {stage0_42[198]},
      {stage1_42[114]}
   );
   gpc1_1 gpc2142 (
      {stage0_42[199]},
      {stage1_42[115]}
   );
   gpc1_1 gpc2143 (
      {stage0_42[200]},
      {stage1_42[116]}
   );
   gpc1_1 gpc2144 (
      {stage0_42[201]},
      {stage1_42[117]}
   );
   gpc1_1 gpc2145 (
      {stage0_42[202]},
      {stage1_42[118]}
   );
   gpc1_1 gpc2146 (
      {stage0_42[203]},
      {stage1_42[119]}
   );
   gpc1_1 gpc2147 (
      {stage0_42[204]},
      {stage1_42[120]}
   );
   gpc1_1 gpc2148 (
      {stage0_42[205]},
      {stage1_42[121]}
   );
   gpc1_1 gpc2149 (
      {stage0_42[206]},
      {stage1_42[122]}
   );
   gpc1_1 gpc2150 (
      {stage0_42[207]},
      {stage1_42[123]}
   );
   gpc1_1 gpc2151 (
      {stage0_42[208]},
      {stage1_42[124]}
   );
   gpc1_1 gpc2152 (
      {stage0_42[209]},
      {stage1_42[125]}
   );
   gpc1_1 gpc2153 (
      {stage0_42[210]},
      {stage1_42[126]}
   );
   gpc1_1 gpc2154 (
      {stage0_42[211]},
      {stage1_42[127]}
   );
   gpc1_1 gpc2155 (
      {stage0_42[212]},
      {stage1_42[128]}
   );
   gpc1_1 gpc2156 (
      {stage0_42[213]},
      {stage1_42[129]}
   );
   gpc1_1 gpc2157 (
      {stage0_42[214]},
      {stage1_42[130]}
   );
   gpc1_1 gpc2158 (
      {stage0_42[215]},
      {stage1_42[131]}
   );
   gpc1_1 gpc2159 (
      {stage0_42[216]},
      {stage1_42[132]}
   );
   gpc1_1 gpc2160 (
      {stage0_42[217]},
      {stage1_42[133]}
   );
   gpc1_1 gpc2161 (
      {stage0_42[218]},
      {stage1_42[134]}
   );
   gpc1_1 gpc2162 (
      {stage0_42[219]},
      {stage1_42[135]}
   );
   gpc1_1 gpc2163 (
      {stage0_42[220]},
      {stage1_42[136]}
   );
   gpc1_1 gpc2164 (
      {stage0_42[221]},
      {stage1_42[137]}
   );
   gpc1_1 gpc2165 (
      {stage0_42[222]},
      {stage1_42[138]}
   );
   gpc1_1 gpc2166 (
      {stage0_42[223]},
      {stage1_42[139]}
   );
   gpc1_1 gpc2167 (
      {stage0_42[224]},
      {stage1_42[140]}
   );
   gpc1_1 gpc2168 (
      {stage0_42[225]},
      {stage1_42[141]}
   );
   gpc1_1 gpc2169 (
      {stage0_42[226]},
      {stage1_42[142]}
   );
   gpc1_1 gpc2170 (
      {stage0_42[227]},
      {stage1_42[143]}
   );
   gpc1_1 gpc2171 (
      {stage0_42[228]},
      {stage1_42[144]}
   );
   gpc1_1 gpc2172 (
      {stage0_42[229]},
      {stage1_42[145]}
   );
   gpc1_1 gpc2173 (
      {stage0_42[230]},
      {stage1_42[146]}
   );
   gpc1_1 gpc2174 (
      {stage0_42[231]},
      {stage1_42[147]}
   );
   gpc1_1 gpc2175 (
      {stage0_42[232]},
      {stage1_42[148]}
   );
   gpc1_1 gpc2176 (
      {stage0_42[233]},
      {stage1_42[149]}
   );
   gpc1_1 gpc2177 (
      {stage0_42[234]},
      {stage1_42[150]}
   );
   gpc1_1 gpc2178 (
      {stage0_42[235]},
      {stage1_42[151]}
   );
   gpc1_1 gpc2179 (
      {stage0_42[236]},
      {stage1_42[152]}
   );
   gpc1_1 gpc2180 (
      {stage0_42[237]},
      {stage1_42[153]}
   );
   gpc1_1 gpc2181 (
      {stage0_42[238]},
      {stage1_42[154]}
   );
   gpc1_1 gpc2182 (
      {stage0_42[239]},
      {stage1_42[155]}
   );
   gpc1_1 gpc2183 (
      {stage0_42[240]},
      {stage1_42[156]}
   );
   gpc1_1 gpc2184 (
      {stage0_42[241]},
      {stage1_42[157]}
   );
   gpc1_1 gpc2185 (
      {stage0_42[242]},
      {stage1_42[158]}
   );
   gpc1_1 gpc2186 (
      {stage0_42[243]},
      {stage1_42[159]}
   );
   gpc1_1 gpc2187 (
      {stage0_42[244]},
      {stage1_42[160]}
   );
   gpc1_1 gpc2188 (
      {stage0_42[245]},
      {stage1_42[161]}
   );
   gpc1_1 gpc2189 (
      {stage0_42[246]},
      {stage1_42[162]}
   );
   gpc1_1 gpc2190 (
      {stage0_42[247]},
      {stage1_42[163]}
   );
   gpc1_1 gpc2191 (
      {stage0_42[248]},
      {stage1_42[164]}
   );
   gpc1_1 gpc2192 (
      {stage0_42[249]},
      {stage1_42[165]}
   );
   gpc1_1 gpc2193 (
      {stage0_42[250]},
      {stage1_42[166]}
   );
   gpc1_1 gpc2194 (
      {stage0_42[251]},
      {stage1_42[167]}
   );
   gpc1_1 gpc2195 (
      {stage0_42[252]},
      {stage1_42[168]}
   );
   gpc1_1 gpc2196 (
      {stage0_42[253]},
      {stage1_42[169]}
   );
   gpc1_1 gpc2197 (
      {stage0_42[254]},
      {stage1_42[170]}
   );
   gpc1_1 gpc2198 (
      {stage0_42[255]},
      {stage1_42[171]}
   );
   gpc1_1 gpc2199 (
      {stage0_43[250]},
      {stage1_43[73]}
   );
   gpc1_1 gpc2200 (
      {stage0_43[251]},
      {stage1_43[74]}
   );
   gpc1_1 gpc2201 (
      {stage0_43[252]},
      {stage1_43[75]}
   );
   gpc1_1 gpc2202 (
      {stage0_43[253]},
      {stage1_43[76]}
   );
   gpc1_1 gpc2203 (
      {stage0_43[254]},
      {stage1_43[77]}
   );
   gpc1_1 gpc2204 (
      {stage0_43[255]},
      {stage1_43[78]}
   );
   gpc1_1 gpc2205 (
      {stage0_44[203]},
      {stage1_44[93]}
   );
   gpc1_1 gpc2206 (
      {stage0_44[204]},
      {stage1_44[94]}
   );
   gpc1_1 gpc2207 (
      {stage0_44[205]},
      {stage1_44[95]}
   );
   gpc1_1 gpc2208 (
      {stage0_44[206]},
      {stage1_44[96]}
   );
   gpc1_1 gpc2209 (
      {stage0_44[207]},
      {stage1_44[97]}
   );
   gpc1_1 gpc2210 (
      {stage0_44[208]},
      {stage1_44[98]}
   );
   gpc1_1 gpc2211 (
      {stage0_44[209]},
      {stage1_44[99]}
   );
   gpc1_1 gpc2212 (
      {stage0_44[210]},
      {stage1_44[100]}
   );
   gpc1_1 gpc2213 (
      {stage0_44[211]},
      {stage1_44[101]}
   );
   gpc1_1 gpc2214 (
      {stage0_44[212]},
      {stage1_44[102]}
   );
   gpc1_1 gpc2215 (
      {stage0_44[213]},
      {stage1_44[103]}
   );
   gpc1_1 gpc2216 (
      {stage0_44[214]},
      {stage1_44[104]}
   );
   gpc1_1 gpc2217 (
      {stage0_44[215]},
      {stage1_44[105]}
   );
   gpc1_1 gpc2218 (
      {stage0_44[216]},
      {stage1_44[106]}
   );
   gpc1_1 gpc2219 (
      {stage0_44[217]},
      {stage1_44[107]}
   );
   gpc1_1 gpc2220 (
      {stage0_44[218]},
      {stage1_44[108]}
   );
   gpc1_1 gpc2221 (
      {stage0_44[219]},
      {stage1_44[109]}
   );
   gpc1_1 gpc2222 (
      {stage0_44[220]},
      {stage1_44[110]}
   );
   gpc1_1 gpc2223 (
      {stage0_44[221]},
      {stage1_44[111]}
   );
   gpc1_1 gpc2224 (
      {stage0_44[222]},
      {stage1_44[112]}
   );
   gpc1_1 gpc2225 (
      {stage0_44[223]},
      {stage1_44[113]}
   );
   gpc1_1 gpc2226 (
      {stage0_44[224]},
      {stage1_44[114]}
   );
   gpc1_1 gpc2227 (
      {stage0_44[225]},
      {stage1_44[115]}
   );
   gpc1_1 gpc2228 (
      {stage0_44[226]},
      {stage1_44[116]}
   );
   gpc1_1 gpc2229 (
      {stage0_44[227]},
      {stage1_44[117]}
   );
   gpc1_1 gpc2230 (
      {stage0_44[228]},
      {stage1_44[118]}
   );
   gpc1_1 gpc2231 (
      {stage0_44[229]},
      {stage1_44[119]}
   );
   gpc1_1 gpc2232 (
      {stage0_44[230]},
      {stage1_44[120]}
   );
   gpc1_1 gpc2233 (
      {stage0_44[231]},
      {stage1_44[121]}
   );
   gpc1_1 gpc2234 (
      {stage0_44[232]},
      {stage1_44[122]}
   );
   gpc1_1 gpc2235 (
      {stage0_44[233]},
      {stage1_44[123]}
   );
   gpc1_1 gpc2236 (
      {stage0_44[234]},
      {stage1_44[124]}
   );
   gpc1_1 gpc2237 (
      {stage0_44[235]},
      {stage1_44[125]}
   );
   gpc1_1 gpc2238 (
      {stage0_44[236]},
      {stage1_44[126]}
   );
   gpc1_1 gpc2239 (
      {stage0_44[237]},
      {stage1_44[127]}
   );
   gpc1_1 gpc2240 (
      {stage0_44[238]},
      {stage1_44[128]}
   );
   gpc1_1 gpc2241 (
      {stage0_44[239]},
      {stage1_44[129]}
   );
   gpc1_1 gpc2242 (
      {stage0_44[240]},
      {stage1_44[130]}
   );
   gpc1_1 gpc2243 (
      {stage0_44[241]},
      {stage1_44[131]}
   );
   gpc1_1 gpc2244 (
      {stage0_44[242]},
      {stage1_44[132]}
   );
   gpc1_1 gpc2245 (
      {stage0_44[243]},
      {stage1_44[133]}
   );
   gpc1_1 gpc2246 (
      {stage0_44[244]},
      {stage1_44[134]}
   );
   gpc1_1 gpc2247 (
      {stage0_44[245]},
      {stage1_44[135]}
   );
   gpc1_1 gpc2248 (
      {stage0_44[246]},
      {stage1_44[136]}
   );
   gpc1_1 gpc2249 (
      {stage0_44[247]},
      {stage1_44[137]}
   );
   gpc1_1 gpc2250 (
      {stage0_44[248]},
      {stage1_44[138]}
   );
   gpc1_1 gpc2251 (
      {stage0_44[249]},
      {stage1_44[139]}
   );
   gpc1_1 gpc2252 (
      {stage0_44[250]},
      {stage1_44[140]}
   );
   gpc1_1 gpc2253 (
      {stage0_44[251]},
      {stage1_44[141]}
   );
   gpc1_1 gpc2254 (
      {stage0_44[252]},
      {stage1_44[142]}
   );
   gpc1_1 gpc2255 (
      {stage0_44[253]},
      {stage1_44[143]}
   );
   gpc1_1 gpc2256 (
      {stage0_44[254]},
      {stage1_44[144]}
   );
   gpc1_1 gpc2257 (
      {stage0_44[255]},
      {stage1_44[145]}
   );
   gpc1_1 gpc2258 (
      {stage0_45[200]},
      {stage1_45[103]}
   );
   gpc1_1 gpc2259 (
      {stage0_45[201]},
      {stage1_45[104]}
   );
   gpc1_1 gpc2260 (
      {stage0_45[202]},
      {stage1_45[105]}
   );
   gpc1_1 gpc2261 (
      {stage0_45[203]},
      {stage1_45[106]}
   );
   gpc1_1 gpc2262 (
      {stage0_45[204]},
      {stage1_45[107]}
   );
   gpc1_1 gpc2263 (
      {stage0_45[205]},
      {stage1_45[108]}
   );
   gpc1_1 gpc2264 (
      {stage0_45[206]},
      {stage1_45[109]}
   );
   gpc1_1 gpc2265 (
      {stage0_45[207]},
      {stage1_45[110]}
   );
   gpc1_1 gpc2266 (
      {stage0_45[208]},
      {stage1_45[111]}
   );
   gpc1_1 gpc2267 (
      {stage0_45[209]},
      {stage1_45[112]}
   );
   gpc1_1 gpc2268 (
      {stage0_45[210]},
      {stage1_45[113]}
   );
   gpc1_1 gpc2269 (
      {stage0_45[211]},
      {stage1_45[114]}
   );
   gpc1_1 gpc2270 (
      {stage0_45[212]},
      {stage1_45[115]}
   );
   gpc1_1 gpc2271 (
      {stage0_45[213]},
      {stage1_45[116]}
   );
   gpc1_1 gpc2272 (
      {stage0_45[214]},
      {stage1_45[117]}
   );
   gpc1_1 gpc2273 (
      {stage0_45[215]},
      {stage1_45[118]}
   );
   gpc1_1 gpc2274 (
      {stage0_45[216]},
      {stage1_45[119]}
   );
   gpc1_1 gpc2275 (
      {stage0_45[217]},
      {stage1_45[120]}
   );
   gpc1_1 gpc2276 (
      {stage0_45[218]},
      {stage1_45[121]}
   );
   gpc1_1 gpc2277 (
      {stage0_45[219]},
      {stage1_45[122]}
   );
   gpc1_1 gpc2278 (
      {stage0_45[220]},
      {stage1_45[123]}
   );
   gpc1_1 gpc2279 (
      {stage0_45[221]},
      {stage1_45[124]}
   );
   gpc1_1 gpc2280 (
      {stage0_45[222]},
      {stage1_45[125]}
   );
   gpc1_1 gpc2281 (
      {stage0_45[223]},
      {stage1_45[126]}
   );
   gpc1_1 gpc2282 (
      {stage0_45[224]},
      {stage1_45[127]}
   );
   gpc1_1 gpc2283 (
      {stage0_45[225]},
      {stage1_45[128]}
   );
   gpc1_1 gpc2284 (
      {stage0_45[226]},
      {stage1_45[129]}
   );
   gpc1_1 gpc2285 (
      {stage0_45[227]},
      {stage1_45[130]}
   );
   gpc1_1 gpc2286 (
      {stage0_45[228]},
      {stage1_45[131]}
   );
   gpc1_1 gpc2287 (
      {stage0_45[229]},
      {stage1_45[132]}
   );
   gpc1_1 gpc2288 (
      {stage0_45[230]},
      {stage1_45[133]}
   );
   gpc1_1 gpc2289 (
      {stage0_45[231]},
      {stage1_45[134]}
   );
   gpc1_1 gpc2290 (
      {stage0_45[232]},
      {stage1_45[135]}
   );
   gpc1_1 gpc2291 (
      {stage0_45[233]},
      {stage1_45[136]}
   );
   gpc1_1 gpc2292 (
      {stage0_45[234]},
      {stage1_45[137]}
   );
   gpc1_1 gpc2293 (
      {stage0_45[235]},
      {stage1_45[138]}
   );
   gpc1_1 gpc2294 (
      {stage0_45[236]},
      {stage1_45[139]}
   );
   gpc1_1 gpc2295 (
      {stage0_45[237]},
      {stage1_45[140]}
   );
   gpc1_1 gpc2296 (
      {stage0_45[238]},
      {stage1_45[141]}
   );
   gpc1_1 gpc2297 (
      {stage0_45[239]},
      {stage1_45[142]}
   );
   gpc1_1 gpc2298 (
      {stage0_45[240]},
      {stage1_45[143]}
   );
   gpc1_1 gpc2299 (
      {stage0_45[241]},
      {stage1_45[144]}
   );
   gpc1_1 gpc2300 (
      {stage0_45[242]},
      {stage1_45[145]}
   );
   gpc1_1 gpc2301 (
      {stage0_45[243]},
      {stage1_45[146]}
   );
   gpc1_1 gpc2302 (
      {stage0_45[244]},
      {stage1_45[147]}
   );
   gpc1_1 gpc2303 (
      {stage0_45[245]},
      {stage1_45[148]}
   );
   gpc1_1 gpc2304 (
      {stage0_45[246]},
      {stage1_45[149]}
   );
   gpc1_1 gpc2305 (
      {stage0_45[247]},
      {stage1_45[150]}
   );
   gpc1_1 gpc2306 (
      {stage0_45[248]},
      {stage1_45[151]}
   );
   gpc1_1 gpc2307 (
      {stage0_45[249]},
      {stage1_45[152]}
   );
   gpc1_1 gpc2308 (
      {stage0_45[250]},
      {stage1_45[153]}
   );
   gpc1_1 gpc2309 (
      {stage0_45[251]},
      {stage1_45[154]}
   );
   gpc1_1 gpc2310 (
      {stage0_45[252]},
      {stage1_45[155]}
   );
   gpc1_1 gpc2311 (
      {stage0_45[253]},
      {stage1_45[156]}
   );
   gpc1_1 gpc2312 (
      {stage0_45[254]},
      {stage1_45[157]}
   );
   gpc1_1 gpc2313 (
      {stage0_45[255]},
      {stage1_45[158]}
   );
   gpc1_1 gpc2314 (
      {stage0_46[237]},
      {stage1_46[82]}
   );
   gpc1_1 gpc2315 (
      {stage0_46[238]},
      {stage1_46[83]}
   );
   gpc1_1 gpc2316 (
      {stage0_46[239]},
      {stage1_46[84]}
   );
   gpc1_1 gpc2317 (
      {stage0_46[240]},
      {stage1_46[85]}
   );
   gpc1_1 gpc2318 (
      {stage0_46[241]},
      {stage1_46[86]}
   );
   gpc1_1 gpc2319 (
      {stage0_46[242]},
      {stage1_46[87]}
   );
   gpc1_1 gpc2320 (
      {stage0_46[243]},
      {stage1_46[88]}
   );
   gpc1_1 gpc2321 (
      {stage0_46[244]},
      {stage1_46[89]}
   );
   gpc1_1 gpc2322 (
      {stage0_46[245]},
      {stage1_46[90]}
   );
   gpc1_1 gpc2323 (
      {stage0_46[246]},
      {stage1_46[91]}
   );
   gpc1_1 gpc2324 (
      {stage0_46[247]},
      {stage1_46[92]}
   );
   gpc1_1 gpc2325 (
      {stage0_46[248]},
      {stage1_46[93]}
   );
   gpc1_1 gpc2326 (
      {stage0_46[249]},
      {stage1_46[94]}
   );
   gpc1_1 gpc2327 (
      {stage0_46[250]},
      {stage1_46[95]}
   );
   gpc1_1 gpc2328 (
      {stage0_46[251]},
      {stage1_46[96]}
   );
   gpc1_1 gpc2329 (
      {stage0_46[252]},
      {stage1_46[97]}
   );
   gpc1_1 gpc2330 (
      {stage0_46[253]},
      {stage1_46[98]}
   );
   gpc1_1 gpc2331 (
      {stage0_46[254]},
      {stage1_46[99]}
   );
   gpc1_1 gpc2332 (
      {stage0_46[255]},
      {stage1_46[100]}
   );
   gpc1_1 gpc2333 (
      {stage0_47[205]},
      {stage1_47[79]}
   );
   gpc1_1 gpc2334 (
      {stage0_47[206]},
      {stage1_47[80]}
   );
   gpc1_1 gpc2335 (
      {stage0_47[207]},
      {stage1_47[81]}
   );
   gpc1_1 gpc2336 (
      {stage0_47[208]},
      {stage1_47[82]}
   );
   gpc1_1 gpc2337 (
      {stage0_47[209]},
      {stage1_47[83]}
   );
   gpc1_1 gpc2338 (
      {stage0_47[210]},
      {stage1_47[84]}
   );
   gpc1_1 gpc2339 (
      {stage0_47[211]},
      {stage1_47[85]}
   );
   gpc1_1 gpc2340 (
      {stage0_47[212]},
      {stage1_47[86]}
   );
   gpc1_1 gpc2341 (
      {stage0_47[213]},
      {stage1_47[87]}
   );
   gpc1_1 gpc2342 (
      {stage0_47[214]},
      {stage1_47[88]}
   );
   gpc1_1 gpc2343 (
      {stage0_47[215]},
      {stage1_47[89]}
   );
   gpc1_1 gpc2344 (
      {stage0_47[216]},
      {stage1_47[90]}
   );
   gpc1_1 gpc2345 (
      {stage0_47[217]},
      {stage1_47[91]}
   );
   gpc1_1 gpc2346 (
      {stage0_47[218]},
      {stage1_47[92]}
   );
   gpc1_1 gpc2347 (
      {stage0_47[219]},
      {stage1_47[93]}
   );
   gpc1_1 gpc2348 (
      {stage0_47[220]},
      {stage1_47[94]}
   );
   gpc1_1 gpc2349 (
      {stage0_47[221]},
      {stage1_47[95]}
   );
   gpc1_1 gpc2350 (
      {stage0_47[222]},
      {stage1_47[96]}
   );
   gpc1_1 gpc2351 (
      {stage0_47[223]},
      {stage1_47[97]}
   );
   gpc1_1 gpc2352 (
      {stage0_47[224]},
      {stage1_47[98]}
   );
   gpc1_1 gpc2353 (
      {stage0_47[225]},
      {stage1_47[99]}
   );
   gpc1_1 gpc2354 (
      {stage0_47[226]},
      {stage1_47[100]}
   );
   gpc1_1 gpc2355 (
      {stage0_47[227]},
      {stage1_47[101]}
   );
   gpc1_1 gpc2356 (
      {stage0_47[228]},
      {stage1_47[102]}
   );
   gpc1_1 gpc2357 (
      {stage0_47[229]},
      {stage1_47[103]}
   );
   gpc1_1 gpc2358 (
      {stage0_47[230]},
      {stage1_47[104]}
   );
   gpc1_1 gpc2359 (
      {stage0_47[231]},
      {stage1_47[105]}
   );
   gpc1_1 gpc2360 (
      {stage0_47[232]},
      {stage1_47[106]}
   );
   gpc1_1 gpc2361 (
      {stage0_47[233]},
      {stage1_47[107]}
   );
   gpc1_1 gpc2362 (
      {stage0_47[234]},
      {stage1_47[108]}
   );
   gpc1_1 gpc2363 (
      {stage0_47[235]},
      {stage1_47[109]}
   );
   gpc1_1 gpc2364 (
      {stage0_47[236]},
      {stage1_47[110]}
   );
   gpc1_1 gpc2365 (
      {stage0_47[237]},
      {stage1_47[111]}
   );
   gpc1_1 gpc2366 (
      {stage0_47[238]},
      {stage1_47[112]}
   );
   gpc1_1 gpc2367 (
      {stage0_47[239]},
      {stage1_47[113]}
   );
   gpc1_1 gpc2368 (
      {stage0_47[240]},
      {stage1_47[114]}
   );
   gpc1_1 gpc2369 (
      {stage0_47[241]},
      {stage1_47[115]}
   );
   gpc1_1 gpc2370 (
      {stage0_47[242]},
      {stage1_47[116]}
   );
   gpc1_1 gpc2371 (
      {stage0_47[243]},
      {stage1_47[117]}
   );
   gpc1_1 gpc2372 (
      {stage0_47[244]},
      {stage1_47[118]}
   );
   gpc1_1 gpc2373 (
      {stage0_47[245]},
      {stage1_47[119]}
   );
   gpc1_1 gpc2374 (
      {stage0_47[246]},
      {stage1_47[120]}
   );
   gpc1_1 gpc2375 (
      {stage0_47[247]},
      {stage1_47[121]}
   );
   gpc1_1 gpc2376 (
      {stage0_47[248]},
      {stage1_47[122]}
   );
   gpc1_1 gpc2377 (
      {stage0_47[249]},
      {stage1_47[123]}
   );
   gpc1_1 gpc2378 (
      {stage0_47[250]},
      {stage1_47[124]}
   );
   gpc1_1 gpc2379 (
      {stage0_47[251]},
      {stage1_47[125]}
   );
   gpc1_1 gpc2380 (
      {stage0_47[252]},
      {stage1_47[126]}
   );
   gpc1_1 gpc2381 (
      {stage0_47[253]},
      {stage1_47[127]}
   );
   gpc1_1 gpc2382 (
      {stage0_47[254]},
      {stage1_47[128]}
   );
   gpc1_1 gpc2383 (
      {stage0_47[255]},
      {stage1_47[129]}
   );
   gpc1_1 gpc2384 (
      {stage0_48[253]},
      {stage1_48[105]}
   );
   gpc1_1 gpc2385 (
      {stage0_48[254]},
      {stage1_48[106]}
   );
   gpc1_1 gpc2386 (
      {stage0_48[255]},
      {stage1_48[107]}
   );
   gpc1_1 gpc2387 (
      {stage0_49[209]},
      {stage1_49[105]}
   );
   gpc1_1 gpc2388 (
      {stage0_49[210]},
      {stage1_49[106]}
   );
   gpc1_1 gpc2389 (
      {stage0_49[211]},
      {stage1_49[107]}
   );
   gpc1_1 gpc2390 (
      {stage0_49[212]},
      {stage1_49[108]}
   );
   gpc1_1 gpc2391 (
      {stage0_49[213]},
      {stage1_49[109]}
   );
   gpc1_1 gpc2392 (
      {stage0_49[214]},
      {stage1_49[110]}
   );
   gpc1_1 gpc2393 (
      {stage0_49[215]},
      {stage1_49[111]}
   );
   gpc1_1 gpc2394 (
      {stage0_49[216]},
      {stage1_49[112]}
   );
   gpc1_1 gpc2395 (
      {stage0_49[217]},
      {stage1_49[113]}
   );
   gpc1_1 gpc2396 (
      {stage0_49[218]},
      {stage1_49[114]}
   );
   gpc1_1 gpc2397 (
      {stage0_49[219]},
      {stage1_49[115]}
   );
   gpc1_1 gpc2398 (
      {stage0_49[220]},
      {stage1_49[116]}
   );
   gpc1_1 gpc2399 (
      {stage0_49[221]},
      {stage1_49[117]}
   );
   gpc1_1 gpc2400 (
      {stage0_49[222]},
      {stage1_49[118]}
   );
   gpc1_1 gpc2401 (
      {stage0_49[223]},
      {stage1_49[119]}
   );
   gpc1_1 gpc2402 (
      {stage0_49[224]},
      {stage1_49[120]}
   );
   gpc1_1 gpc2403 (
      {stage0_49[225]},
      {stage1_49[121]}
   );
   gpc1_1 gpc2404 (
      {stage0_49[226]},
      {stage1_49[122]}
   );
   gpc1_1 gpc2405 (
      {stage0_49[227]},
      {stage1_49[123]}
   );
   gpc1_1 gpc2406 (
      {stage0_49[228]},
      {stage1_49[124]}
   );
   gpc1_1 gpc2407 (
      {stage0_49[229]},
      {stage1_49[125]}
   );
   gpc1_1 gpc2408 (
      {stage0_49[230]},
      {stage1_49[126]}
   );
   gpc1_1 gpc2409 (
      {stage0_49[231]},
      {stage1_49[127]}
   );
   gpc1_1 gpc2410 (
      {stage0_49[232]},
      {stage1_49[128]}
   );
   gpc1_1 gpc2411 (
      {stage0_49[233]},
      {stage1_49[129]}
   );
   gpc1_1 gpc2412 (
      {stage0_49[234]},
      {stage1_49[130]}
   );
   gpc1_1 gpc2413 (
      {stage0_49[235]},
      {stage1_49[131]}
   );
   gpc1_1 gpc2414 (
      {stage0_49[236]},
      {stage1_49[132]}
   );
   gpc1_1 gpc2415 (
      {stage0_49[237]},
      {stage1_49[133]}
   );
   gpc1_1 gpc2416 (
      {stage0_49[238]},
      {stage1_49[134]}
   );
   gpc1_1 gpc2417 (
      {stage0_49[239]},
      {stage1_49[135]}
   );
   gpc1_1 gpc2418 (
      {stage0_49[240]},
      {stage1_49[136]}
   );
   gpc1_1 gpc2419 (
      {stage0_49[241]},
      {stage1_49[137]}
   );
   gpc1_1 gpc2420 (
      {stage0_49[242]},
      {stage1_49[138]}
   );
   gpc1_1 gpc2421 (
      {stage0_49[243]},
      {stage1_49[139]}
   );
   gpc1_1 gpc2422 (
      {stage0_49[244]},
      {stage1_49[140]}
   );
   gpc1_1 gpc2423 (
      {stage0_49[245]},
      {stage1_49[141]}
   );
   gpc1_1 gpc2424 (
      {stage0_49[246]},
      {stage1_49[142]}
   );
   gpc1_1 gpc2425 (
      {stage0_49[247]},
      {stage1_49[143]}
   );
   gpc1_1 gpc2426 (
      {stage0_49[248]},
      {stage1_49[144]}
   );
   gpc1_1 gpc2427 (
      {stage0_49[249]},
      {stage1_49[145]}
   );
   gpc1_1 gpc2428 (
      {stage0_49[250]},
      {stage1_49[146]}
   );
   gpc1_1 gpc2429 (
      {stage0_49[251]},
      {stage1_49[147]}
   );
   gpc1_1 gpc2430 (
      {stage0_49[252]},
      {stage1_49[148]}
   );
   gpc1_1 gpc2431 (
      {stage0_49[253]},
      {stage1_49[149]}
   );
   gpc1_1 gpc2432 (
      {stage0_49[254]},
      {stage1_49[150]}
   );
   gpc1_1 gpc2433 (
      {stage0_49[255]},
      {stage1_49[151]}
   );
   gpc1_1 gpc2434 (
      {stage0_50[243]},
      {stage1_50[86]}
   );
   gpc1_1 gpc2435 (
      {stage0_50[244]},
      {stage1_50[87]}
   );
   gpc1_1 gpc2436 (
      {stage0_50[245]},
      {stage1_50[88]}
   );
   gpc1_1 gpc2437 (
      {stage0_50[246]},
      {stage1_50[89]}
   );
   gpc1_1 gpc2438 (
      {stage0_50[247]},
      {stage1_50[90]}
   );
   gpc1_1 gpc2439 (
      {stage0_50[248]},
      {stage1_50[91]}
   );
   gpc1_1 gpc2440 (
      {stage0_50[249]},
      {stage1_50[92]}
   );
   gpc1_1 gpc2441 (
      {stage0_50[250]},
      {stage1_50[93]}
   );
   gpc1_1 gpc2442 (
      {stage0_50[251]},
      {stage1_50[94]}
   );
   gpc1_1 gpc2443 (
      {stage0_50[252]},
      {stage1_50[95]}
   );
   gpc1_1 gpc2444 (
      {stage0_50[253]},
      {stage1_50[96]}
   );
   gpc1_1 gpc2445 (
      {stage0_50[254]},
      {stage1_50[97]}
   );
   gpc1_1 gpc2446 (
      {stage0_50[255]},
      {stage1_50[98]}
   );
   gpc1_1 gpc2447 (
      {stage0_51[236]},
      {stage1_51[86]}
   );
   gpc1_1 gpc2448 (
      {stage0_51[237]},
      {stage1_51[87]}
   );
   gpc1_1 gpc2449 (
      {stage0_51[238]},
      {stage1_51[88]}
   );
   gpc1_1 gpc2450 (
      {stage0_51[239]},
      {stage1_51[89]}
   );
   gpc1_1 gpc2451 (
      {stage0_51[240]},
      {stage1_51[90]}
   );
   gpc1_1 gpc2452 (
      {stage0_51[241]},
      {stage1_51[91]}
   );
   gpc1_1 gpc2453 (
      {stage0_51[242]},
      {stage1_51[92]}
   );
   gpc1_1 gpc2454 (
      {stage0_51[243]},
      {stage1_51[93]}
   );
   gpc1_1 gpc2455 (
      {stage0_51[244]},
      {stage1_51[94]}
   );
   gpc1_1 gpc2456 (
      {stage0_51[245]},
      {stage1_51[95]}
   );
   gpc1_1 gpc2457 (
      {stage0_51[246]},
      {stage1_51[96]}
   );
   gpc1_1 gpc2458 (
      {stage0_51[247]},
      {stage1_51[97]}
   );
   gpc1_1 gpc2459 (
      {stage0_51[248]},
      {stage1_51[98]}
   );
   gpc1_1 gpc2460 (
      {stage0_51[249]},
      {stage1_51[99]}
   );
   gpc1_1 gpc2461 (
      {stage0_51[250]},
      {stage1_51[100]}
   );
   gpc1_1 gpc2462 (
      {stage0_51[251]},
      {stage1_51[101]}
   );
   gpc1_1 gpc2463 (
      {stage0_51[252]},
      {stage1_51[102]}
   );
   gpc1_1 gpc2464 (
      {stage0_51[253]},
      {stage1_51[103]}
   );
   gpc1_1 gpc2465 (
      {stage0_51[254]},
      {stage1_51[104]}
   );
   gpc1_1 gpc2466 (
      {stage0_51[255]},
      {stage1_51[105]}
   );
   gpc1_1 gpc2467 (
      {stage0_52[223]},
      {stage1_52[107]}
   );
   gpc1_1 gpc2468 (
      {stage0_52[224]},
      {stage1_52[108]}
   );
   gpc1_1 gpc2469 (
      {stage0_52[225]},
      {stage1_52[109]}
   );
   gpc1_1 gpc2470 (
      {stage0_52[226]},
      {stage1_52[110]}
   );
   gpc1_1 gpc2471 (
      {stage0_52[227]},
      {stage1_52[111]}
   );
   gpc1_1 gpc2472 (
      {stage0_52[228]},
      {stage1_52[112]}
   );
   gpc1_1 gpc2473 (
      {stage0_52[229]},
      {stage1_52[113]}
   );
   gpc1_1 gpc2474 (
      {stage0_52[230]},
      {stage1_52[114]}
   );
   gpc1_1 gpc2475 (
      {stage0_52[231]},
      {stage1_52[115]}
   );
   gpc1_1 gpc2476 (
      {stage0_52[232]},
      {stage1_52[116]}
   );
   gpc1_1 gpc2477 (
      {stage0_52[233]},
      {stage1_52[117]}
   );
   gpc1_1 gpc2478 (
      {stage0_52[234]},
      {stage1_52[118]}
   );
   gpc1_1 gpc2479 (
      {stage0_52[235]},
      {stage1_52[119]}
   );
   gpc1_1 gpc2480 (
      {stage0_52[236]},
      {stage1_52[120]}
   );
   gpc1_1 gpc2481 (
      {stage0_52[237]},
      {stage1_52[121]}
   );
   gpc1_1 gpc2482 (
      {stage0_52[238]},
      {stage1_52[122]}
   );
   gpc1_1 gpc2483 (
      {stage0_52[239]},
      {stage1_52[123]}
   );
   gpc1_1 gpc2484 (
      {stage0_52[240]},
      {stage1_52[124]}
   );
   gpc1_1 gpc2485 (
      {stage0_52[241]},
      {stage1_52[125]}
   );
   gpc1_1 gpc2486 (
      {stage0_52[242]},
      {stage1_52[126]}
   );
   gpc1_1 gpc2487 (
      {stage0_52[243]},
      {stage1_52[127]}
   );
   gpc1_1 gpc2488 (
      {stage0_52[244]},
      {stage1_52[128]}
   );
   gpc1_1 gpc2489 (
      {stage0_52[245]},
      {stage1_52[129]}
   );
   gpc1_1 gpc2490 (
      {stage0_52[246]},
      {stage1_52[130]}
   );
   gpc1_1 gpc2491 (
      {stage0_52[247]},
      {stage1_52[131]}
   );
   gpc1_1 gpc2492 (
      {stage0_52[248]},
      {stage1_52[132]}
   );
   gpc1_1 gpc2493 (
      {stage0_52[249]},
      {stage1_52[133]}
   );
   gpc1_1 gpc2494 (
      {stage0_52[250]},
      {stage1_52[134]}
   );
   gpc1_1 gpc2495 (
      {stage0_52[251]},
      {stage1_52[135]}
   );
   gpc1_1 gpc2496 (
      {stage0_52[252]},
      {stage1_52[136]}
   );
   gpc1_1 gpc2497 (
      {stage0_52[253]},
      {stage1_52[137]}
   );
   gpc1_1 gpc2498 (
      {stage0_52[254]},
      {stage1_52[138]}
   );
   gpc1_1 gpc2499 (
      {stage0_52[255]},
      {stage1_52[139]}
   );
   gpc1_1 gpc2500 (
      {stage0_53[254]},
      {stage1_53[106]}
   );
   gpc1_1 gpc2501 (
      {stage0_53[255]},
      {stage1_53[107]}
   );
   gpc1_1 gpc2502 (
      {stage0_54[178]},
      {stage1_54[82]}
   );
   gpc1_1 gpc2503 (
      {stage0_54[179]},
      {stage1_54[83]}
   );
   gpc1_1 gpc2504 (
      {stage0_54[180]},
      {stage1_54[84]}
   );
   gpc1_1 gpc2505 (
      {stage0_54[181]},
      {stage1_54[85]}
   );
   gpc1_1 gpc2506 (
      {stage0_54[182]},
      {stage1_54[86]}
   );
   gpc1_1 gpc2507 (
      {stage0_54[183]},
      {stage1_54[87]}
   );
   gpc1_1 gpc2508 (
      {stage0_54[184]},
      {stage1_54[88]}
   );
   gpc1_1 gpc2509 (
      {stage0_54[185]},
      {stage1_54[89]}
   );
   gpc1_1 gpc2510 (
      {stage0_54[186]},
      {stage1_54[90]}
   );
   gpc1_1 gpc2511 (
      {stage0_54[187]},
      {stage1_54[91]}
   );
   gpc1_1 gpc2512 (
      {stage0_54[188]},
      {stage1_54[92]}
   );
   gpc1_1 gpc2513 (
      {stage0_54[189]},
      {stage1_54[93]}
   );
   gpc1_1 gpc2514 (
      {stage0_54[190]},
      {stage1_54[94]}
   );
   gpc1_1 gpc2515 (
      {stage0_54[191]},
      {stage1_54[95]}
   );
   gpc1_1 gpc2516 (
      {stage0_54[192]},
      {stage1_54[96]}
   );
   gpc1_1 gpc2517 (
      {stage0_54[193]},
      {stage1_54[97]}
   );
   gpc1_1 gpc2518 (
      {stage0_54[194]},
      {stage1_54[98]}
   );
   gpc1_1 gpc2519 (
      {stage0_54[195]},
      {stage1_54[99]}
   );
   gpc1_1 gpc2520 (
      {stage0_54[196]},
      {stage1_54[100]}
   );
   gpc1_1 gpc2521 (
      {stage0_54[197]},
      {stage1_54[101]}
   );
   gpc1_1 gpc2522 (
      {stage0_54[198]},
      {stage1_54[102]}
   );
   gpc1_1 gpc2523 (
      {stage0_54[199]},
      {stage1_54[103]}
   );
   gpc1_1 gpc2524 (
      {stage0_54[200]},
      {stage1_54[104]}
   );
   gpc1_1 gpc2525 (
      {stage0_54[201]},
      {stage1_54[105]}
   );
   gpc1_1 gpc2526 (
      {stage0_54[202]},
      {stage1_54[106]}
   );
   gpc1_1 gpc2527 (
      {stage0_54[203]},
      {stage1_54[107]}
   );
   gpc1_1 gpc2528 (
      {stage0_54[204]},
      {stage1_54[108]}
   );
   gpc1_1 gpc2529 (
      {stage0_54[205]},
      {stage1_54[109]}
   );
   gpc1_1 gpc2530 (
      {stage0_54[206]},
      {stage1_54[110]}
   );
   gpc1_1 gpc2531 (
      {stage0_54[207]},
      {stage1_54[111]}
   );
   gpc1_1 gpc2532 (
      {stage0_54[208]},
      {stage1_54[112]}
   );
   gpc1_1 gpc2533 (
      {stage0_54[209]},
      {stage1_54[113]}
   );
   gpc1_1 gpc2534 (
      {stage0_54[210]},
      {stage1_54[114]}
   );
   gpc1_1 gpc2535 (
      {stage0_54[211]},
      {stage1_54[115]}
   );
   gpc1_1 gpc2536 (
      {stage0_54[212]},
      {stage1_54[116]}
   );
   gpc1_1 gpc2537 (
      {stage0_54[213]},
      {stage1_54[117]}
   );
   gpc1_1 gpc2538 (
      {stage0_54[214]},
      {stage1_54[118]}
   );
   gpc1_1 gpc2539 (
      {stage0_54[215]},
      {stage1_54[119]}
   );
   gpc1_1 gpc2540 (
      {stage0_54[216]},
      {stage1_54[120]}
   );
   gpc1_1 gpc2541 (
      {stage0_54[217]},
      {stage1_54[121]}
   );
   gpc1_1 gpc2542 (
      {stage0_54[218]},
      {stage1_54[122]}
   );
   gpc1_1 gpc2543 (
      {stage0_54[219]},
      {stage1_54[123]}
   );
   gpc1_1 gpc2544 (
      {stage0_54[220]},
      {stage1_54[124]}
   );
   gpc1_1 gpc2545 (
      {stage0_54[221]},
      {stage1_54[125]}
   );
   gpc1_1 gpc2546 (
      {stage0_54[222]},
      {stage1_54[126]}
   );
   gpc1_1 gpc2547 (
      {stage0_54[223]},
      {stage1_54[127]}
   );
   gpc1_1 gpc2548 (
      {stage0_54[224]},
      {stage1_54[128]}
   );
   gpc1_1 gpc2549 (
      {stage0_54[225]},
      {stage1_54[129]}
   );
   gpc1_1 gpc2550 (
      {stage0_54[226]},
      {stage1_54[130]}
   );
   gpc1_1 gpc2551 (
      {stage0_54[227]},
      {stage1_54[131]}
   );
   gpc1_1 gpc2552 (
      {stage0_54[228]},
      {stage1_54[132]}
   );
   gpc1_1 gpc2553 (
      {stage0_54[229]},
      {stage1_54[133]}
   );
   gpc1_1 gpc2554 (
      {stage0_54[230]},
      {stage1_54[134]}
   );
   gpc1_1 gpc2555 (
      {stage0_54[231]},
      {stage1_54[135]}
   );
   gpc1_1 gpc2556 (
      {stage0_54[232]},
      {stage1_54[136]}
   );
   gpc1_1 gpc2557 (
      {stage0_54[233]},
      {stage1_54[137]}
   );
   gpc1_1 gpc2558 (
      {stage0_54[234]},
      {stage1_54[138]}
   );
   gpc1_1 gpc2559 (
      {stage0_54[235]},
      {stage1_54[139]}
   );
   gpc1_1 gpc2560 (
      {stage0_54[236]},
      {stage1_54[140]}
   );
   gpc1_1 gpc2561 (
      {stage0_54[237]},
      {stage1_54[141]}
   );
   gpc1_1 gpc2562 (
      {stage0_54[238]},
      {stage1_54[142]}
   );
   gpc1_1 gpc2563 (
      {stage0_54[239]},
      {stage1_54[143]}
   );
   gpc1_1 gpc2564 (
      {stage0_54[240]},
      {stage1_54[144]}
   );
   gpc1_1 gpc2565 (
      {stage0_54[241]},
      {stage1_54[145]}
   );
   gpc1_1 gpc2566 (
      {stage0_54[242]},
      {stage1_54[146]}
   );
   gpc1_1 gpc2567 (
      {stage0_54[243]},
      {stage1_54[147]}
   );
   gpc1_1 gpc2568 (
      {stage0_54[244]},
      {stage1_54[148]}
   );
   gpc1_1 gpc2569 (
      {stage0_54[245]},
      {stage1_54[149]}
   );
   gpc1_1 gpc2570 (
      {stage0_54[246]},
      {stage1_54[150]}
   );
   gpc1_1 gpc2571 (
      {stage0_54[247]},
      {stage1_54[151]}
   );
   gpc1_1 gpc2572 (
      {stage0_54[248]},
      {stage1_54[152]}
   );
   gpc1_1 gpc2573 (
      {stage0_54[249]},
      {stage1_54[153]}
   );
   gpc1_1 gpc2574 (
      {stage0_54[250]},
      {stage1_54[154]}
   );
   gpc1_1 gpc2575 (
      {stage0_54[251]},
      {stage1_54[155]}
   );
   gpc1_1 gpc2576 (
      {stage0_54[252]},
      {stage1_54[156]}
   );
   gpc1_1 gpc2577 (
      {stage0_54[253]},
      {stage1_54[157]}
   );
   gpc1_1 gpc2578 (
      {stage0_54[254]},
      {stage1_54[158]}
   );
   gpc1_1 gpc2579 (
      {stage0_54[255]},
      {stage1_54[159]}
   );
   gpc1_1 gpc2580 (
      {stage0_55[250]},
      {stage1_55[84]}
   );
   gpc1_1 gpc2581 (
      {stage0_55[251]},
      {stage1_55[85]}
   );
   gpc1_1 gpc2582 (
      {stage0_55[252]},
      {stage1_55[86]}
   );
   gpc1_1 gpc2583 (
      {stage0_55[253]},
      {stage1_55[87]}
   );
   gpc1_1 gpc2584 (
      {stage0_55[254]},
      {stage1_55[88]}
   );
   gpc1_1 gpc2585 (
      {stage0_55[255]},
      {stage1_55[89]}
   );
   gpc1_1 gpc2586 (
      {stage0_56[176]},
      {stage1_56[98]}
   );
   gpc1_1 gpc2587 (
      {stage0_56[177]},
      {stage1_56[99]}
   );
   gpc1_1 gpc2588 (
      {stage0_56[178]},
      {stage1_56[100]}
   );
   gpc1_1 gpc2589 (
      {stage0_56[179]},
      {stage1_56[101]}
   );
   gpc1_1 gpc2590 (
      {stage0_56[180]},
      {stage1_56[102]}
   );
   gpc1_1 gpc2591 (
      {stage0_56[181]},
      {stage1_56[103]}
   );
   gpc1_1 gpc2592 (
      {stage0_56[182]},
      {stage1_56[104]}
   );
   gpc1_1 gpc2593 (
      {stage0_56[183]},
      {stage1_56[105]}
   );
   gpc1_1 gpc2594 (
      {stage0_56[184]},
      {stage1_56[106]}
   );
   gpc1_1 gpc2595 (
      {stage0_56[185]},
      {stage1_56[107]}
   );
   gpc1_1 gpc2596 (
      {stage0_56[186]},
      {stage1_56[108]}
   );
   gpc1_1 gpc2597 (
      {stage0_56[187]},
      {stage1_56[109]}
   );
   gpc1_1 gpc2598 (
      {stage0_56[188]},
      {stage1_56[110]}
   );
   gpc1_1 gpc2599 (
      {stage0_56[189]},
      {stage1_56[111]}
   );
   gpc1_1 gpc2600 (
      {stage0_56[190]},
      {stage1_56[112]}
   );
   gpc1_1 gpc2601 (
      {stage0_56[191]},
      {stage1_56[113]}
   );
   gpc1_1 gpc2602 (
      {stage0_56[192]},
      {stage1_56[114]}
   );
   gpc1_1 gpc2603 (
      {stage0_56[193]},
      {stage1_56[115]}
   );
   gpc1_1 gpc2604 (
      {stage0_56[194]},
      {stage1_56[116]}
   );
   gpc1_1 gpc2605 (
      {stage0_56[195]},
      {stage1_56[117]}
   );
   gpc1_1 gpc2606 (
      {stage0_56[196]},
      {stage1_56[118]}
   );
   gpc1_1 gpc2607 (
      {stage0_56[197]},
      {stage1_56[119]}
   );
   gpc1_1 gpc2608 (
      {stage0_56[198]},
      {stage1_56[120]}
   );
   gpc1_1 gpc2609 (
      {stage0_56[199]},
      {stage1_56[121]}
   );
   gpc1_1 gpc2610 (
      {stage0_56[200]},
      {stage1_56[122]}
   );
   gpc1_1 gpc2611 (
      {stage0_56[201]},
      {stage1_56[123]}
   );
   gpc1_1 gpc2612 (
      {stage0_56[202]},
      {stage1_56[124]}
   );
   gpc1_1 gpc2613 (
      {stage0_56[203]},
      {stage1_56[125]}
   );
   gpc1_1 gpc2614 (
      {stage0_56[204]},
      {stage1_56[126]}
   );
   gpc1_1 gpc2615 (
      {stage0_56[205]},
      {stage1_56[127]}
   );
   gpc1_1 gpc2616 (
      {stage0_56[206]},
      {stage1_56[128]}
   );
   gpc1_1 gpc2617 (
      {stage0_56[207]},
      {stage1_56[129]}
   );
   gpc1_1 gpc2618 (
      {stage0_56[208]},
      {stage1_56[130]}
   );
   gpc1_1 gpc2619 (
      {stage0_56[209]},
      {stage1_56[131]}
   );
   gpc1_1 gpc2620 (
      {stage0_56[210]},
      {stage1_56[132]}
   );
   gpc1_1 gpc2621 (
      {stage0_56[211]},
      {stage1_56[133]}
   );
   gpc1_1 gpc2622 (
      {stage0_56[212]},
      {stage1_56[134]}
   );
   gpc1_1 gpc2623 (
      {stage0_56[213]},
      {stage1_56[135]}
   );
   gpc1_1 gpc2624 (
      {stage0_56[214]},
      {stage1_56[136]}
   );
   gpc1_1 gpc2625 (
      {stage0_56[215]},
      {stage1_56[137]}
   );
   gpc1_1 gpc2626 (
      {stage0_56[216]},
      {stage1_56[138]}
   );
   gpc1_1 gpc2627 (
      {stage0_56[217]},
      {stage1_56[139]}
   );
   gpc1_1 gpc2628 (
      {stage0_56[218]},
      {stage1_56[140]}
   );
   gpc1_1 gpc2629 (
      {stage0_56[219]},
      {stage1_56[141]}
   );
   gpc1_1 gpc2630 (
      {stage0_56[220]},
      {stage1_56[142]}
   );
   gpc1_1 gpc2631 (
      {stage0_56[221]},
      {stage1_56[143]}
   );
   gpc1_1 gpc2632 (
      {stage0_56[222]},
      {stage1_56[144]}
   );
   gpc1_1 gpc2633 (
      {stage0_56[223]},
      {stage1_56[145]}
   );
   gpc1_1 gpc2634 (
      {stage0_56[224]},
      {stage1_56[146]}
   );
   gpc1_1 gpc2635 (
      {stage0_56[225]},
      {stage1_56[147]}
   );
   gpc1_1 gpc2636 (
      {stage0_56[226]},
      {stage1_56[148]}
   );
   gpc1_1 gpc2637 (
      {stage0_56[227]},
      {stage1_56[149]}
   );
   gpc1_1 gpc2638 (
      {stage0_56[228]},
      {stage1_56[150]}
   );
   gpc1_1 gpc2639 (
      {stage0_56[229]},
      {stage1_56[151]}
   );
   gpc1_1 gpc2640 (
      {stage0_56[230]},
      {stage1_56[152]}
   );
   gpc1_1 gpc2641 (
      {stage0_56[231]},
      {stage1_56[153]}
   );
   gpc1_1 gpc2642 (
      {stage0_56[232]},
      {stage1_56[154]}
   );
   gpc1_1 gpc2643 (
      {stage0_56[233]},
      {stage1_56[155]}
   );
   gpc1_1 gpc2644 (
      {stage0_56[234]},
      {stage1_56[156]}
   );
   gpc1_1 gpc2645 (
      {stage0_56[235]},
      {stage1_56[157]}
   );
   gpc1_1 gpc2646 (
      {stage0_56[236]},
      {stage1_56[158]}
   );
   gpc1_1 gpc2647 (
      {stage0_56[237]},
      {stage1_56[159]}
   );
   gpc1_1 gpc2648 (
      {stage0_56[238]},
      {stage1_56[160]}
   );
   gpc1_1 gpc2649 (
      {stage0_56[239]},
      {stage1_56[161]}
   );
   gpc1_1 gpc2650 (
      {stage0_56[240]},
      {stage1_56[162]}
   );
   gpc1_1 gpc2651 (
      {stage0_56[241]},
      {stage1_56[163]}
   );
   gpc1_1 gpc2652 (
      {stage0_56[242]},
      {stage1_56[164]}
   );
   gpc1_1 gpc2653 (
      {stage0_56[243]},
      {stage1_56[165]}
   );
   gpc1_1 gpc2654 (
      {stage0_56[244]},
      {stage1_56[166]}
   );
   gpc1_1 gpc2655 (
      {stage0_56[245]},
      {stage1_56[167]}
   );
   gpc1_1 gpc2656 (
      {stage0_56[246]},
      {stage1_56[168]}
   );
   gpc1_1 gpc2657 (
      {stage0_56[247]},
      {stage1_56[169]}
   );
   gpc1_1 gpc2658 (
      {stage0_56[248]},
      {stage1_56[170]}
   );
   gpc1_1 gpc2659 (
      {stage0_56[249]},
      {stage1_56[171]}
   );
   gpc1_1 gpc2660 (
      {stage0_56[250]},
      {stage1_56[172]}
   );
   gpc1_1 gpc2661 (
      {stage0_56[251]},
      {stage1_56[173]}
   );
   gpc1_1 gpc2662 (
      {stage0_56[252]},
      {stage1_56[174]}
   );
   gpc1_1 gpc2663 (
      {stage0_56[253]},
      {stage1_56[175]}
   );
   gpc1_1 gpc2664 (
      {stage0_56[254]},
      {stage1_56[176]}
   );
   gpc1_1 gpc2665 (
      {stage0_56[255]},
      {stage1_56[177]}
   );
   gpc1_1 gpc2666 (
      {stage0_57[253]},
      {stage1_57[102]}
   );
   gpc1_1 gpc2667 (
      {stage0_57[254]},
      {stage1_57[103]}
   );
   gpc1_1 gpc2668 (
      {stage0_57[255]},
      {stage1_57[104]}
   );
   gpc1_1 gpc2669 (
      {stage0_58[255]},
      {stage1_58[85]}
   );
   gpc1_1 gpc2670 (
      {stage0_59[194]},
      {stage1_59[86]}
   );
   gpc1_1 gpc2671 (
      {stage0_59[195]},
      {stage1_59[87]}
   );
   gpc1_1 gpc2672 (
      {stage0_59[196]},
      {stage1_59[88]}
   );
   gpc1_1 gpc2673 (
      {stage0_59[197]},
      {stage1_59[89]}
   );
   gpc1_1 gpc2674 (
      {stage0_59[198]},
      {stage1_59[90]}
   );
   gpc1_1 gpc2675 (
      {stage0_59[199]},
      {stage1_59[91]}
   );
   gpc1_1 gpc2676 (
      {stage0_59[200]},
      {stage1_59[92]}
   );
   gpc1_1 gpc2677 (
      {stage0_59[201]},
      {stage1_59[93]}
   );
   gpc1_1 gpc2678 (
      {stage0_59[202]},
      {stage1_59[94]}
   );
   gpc1_1 gpc2679 (
      {stage0_59[203]},
      {stage1_59[95]}
   );
   gpc1_1 gpc2680 (
      {stage0_59[204]},
      {stage1_59[96]}
   );
   gpc1_1 gpc2681 (
      {stage0_59[205]},
      {stage1_59[97]}
   );
   gpc1_1 gpc2682 (
      {stage0_59[206]},
      {stage1_59[98]}
   );
   gpc1_1 gpc2683 (
      {stage0_59[207]},
      {stage1_59[99]}
   );
   gpc1_1 gpc2684 (
      {stage0_59[208]},
      {stage1_59[100]}
   );
   gpc1_1 gpc2685 (
      {stage0_59[209]},
      {stage1_59[101]}
   );
   gpc1_1 gpc2686 (
      {stage0_59[210]},
      {stage1_59[102]}
   );
   gpc1_1 gpc2687 (
      {stage0_59[211]},
      {stage1_59[103]}
   );
   gpc1_1 gpc2688 (
      {stage0_59[212]},
      {stage1_59[104]}
   );
   gpc1_1 gpc2689 (
      {stage0_59[213]},
      {stage1_59[105]}
   );
   gpc1_1 gpc2690 (
      {stage0_59[214]},
      {stage1_59[106]}
   );
   gpc1_1 gpc2691 (
      {stage0_59[215]},
      {stage1_59[107]}
   );
   gpc1_1 gpc2692 (
      {stage0_59[216]},
      {stage1_59[108]}
   );
   gpc1_1 gpc2693 (
      {stage0_59[217]},
      {stage1_59[109]}
   );
   gpc1_1 gpc2694 (
      {stage0_59[218]},
      {stage1_59[110]}
   );
   gpc1_1 gpc2695 (
      {stage0_59[219]},
      {stage1_59[111]}
   );
   gpc1_1 gpc2696 (
      {stage0_59[220]},
      {stage1_59[112]}
   );
   gpc1_1 gpc2697 (
      {stage0_59[221]},
      {stage1_59[113]}
   );
   gpc1_1 gpc2698 (
      {stage0_59[222]},
      {stage1_59[114]}
   );
   gpc1_1 gpc2699 (
      {stage0_59[223]},
      {stage1_59[115]}
   );
   gpc1_1 gpc2700 (
      {stage0_59[224]},
      {stage1_59[116]}
   );
   gpc1_1 gpc2701 (
      {stage0_59[225]},
      {stage1_59[117]}
   );
   gpc1_1 gpc2702 (
      {stage0_59[226]},
      {stage1_59[118]}
   );
   gpc1_1 gpc2703 (
      {stage0_59[227]},
      {stage1_59[119]}
   );
   gpc1_1 gpc2704 (
      {stage0_59[228]},
      {stage1_59[120]}
   );
   gpc1_1 gpc2705 (
      {stage0_59[229]},
      {stage1_59[121]}
   );
   gpc1_1 gpc2706 (
      {stage0_59[230]},
      {stage1_59[122]}
   );
   gpc1_1 gpc2707 (
      {stage0_59[231]},
      {stage1_59[123]}
   );
   gpc1_1 gpc2708 (
      {stage0_59[232]},
      {stage1_59[124]}
   );
   gpc1_1 gpc2709 (
      {stage0_59[233]},
      {stage1_59[125]}
   );
   gpc1_1 gpc2710 (
      {stage0_59[234]},
      {stage1_59[126]}
   );
   gpc1_1 gpc2711 (
      {stage0_59[235]},
      {stage1_59[127]}
   );
   gpc1_1 gpc2712 (
      {stage0_59[236]},
      {stage1_59[128]}
   );
   gpc1_1 gpc2713 (
      {stage0_59[237]},
      {stage1_59[129]}
   );
   gpc1_1 gpc2714 (
      {stage0_59[238]},
      {stage1_59[130]}
   );
   gpc1_1 gpc2715 (
      {stage0_59[239]},
      {stage1_59[131]}
   );
   gpc1_1 gpc2716 (
      {stage0_59[240]},
      {stage1_59[132]}
   );
   gpc1_1 gpc2717 (
      {stage0_59[241]},
      {stage1_59[133]}
   );
   gpc1_1 gpc2718 (
      {stage0_59[242]},
      {stage1_59[134]}
   );
   gpc1_1 gpc2719 (
      {stage0_59[243]},
      {stage1_59[135]}
   );
   gpc1_1 gpc2720 (
      {stage0_59[244]},
      {stage1_59[136]}
   );
   gpc1_1 gpc2721 (
      {stage0_59[245]},
      {stage1_59[137]}
   );
   gpc1_1 gpc2722 (
      {stage0_59[246]},
      {stage1_59[138]}
   );
   gpc1_1 gpc2723 (
      {stage0_59[247]},
      {stage1_59[139]}
   );
   gpc1_1 gpc2724 (
      {stage0_59[248]},
      {stage1_59[140]}
   );
   gpc1_1 gpc2725 (
      {stage0_59[249]},
      {stage1_59[141]}
   );
   gpc1_1 gpc2726 (
      {stage0_59[250]},
      {stage1_59[142]}
   );
   gpc1_1 gpc2727 (
      {stage0_59[251]},
      {stage1_59[143]}
   );
   gpc1_1 gpc2728 (
      {stage0_59[252]},
      {stage1_59[144]}
   );
   gpc1_1 gpc2729 (
      {stage0_59[253]},
      {stage1_59[145]}
   );
   gpc1_1 gpc2730 (
      {stage0_59[254]},
      {stage1_59[146]}
   );
   gpc1_1 gpc2731 (
      {stage0_59[255]},
      {stage1_59[147]}
   );
   gpc1_1 gpc2732 (
      {stage0_60[210]},
      {stage1_60[96]}
   );
   gpc1_1 gpc2733 (
      {stage0_60[211]},
      {stage1_60[97]}
   );
   gpc1_1 gpc2734 (
      {stage0_60[212]},
      {stage1_60[98]}
   );
   gpc1_1 gpc2735 (
      {stage0_60[213]},
      {stage1_60[99]}
   );
   gpc1_1 gpc2736 (
      {stage0_60[214]},
      {stage1_60[100]}
   );
   gpc1_1 gpc2737 (
      {stage0_60[215]},
      {stage1_60[101]}
   );
   gpc1_1 gpc2738 (
      {stage0_60[216]},
      {stage1_60[102]}
   );
   gpc1_1 gpc2739 (
      {stage0_60[217]},
      {stage1_60[103]}
   );
   gpc1_1 gpc2740 (
      {stage0_60[218]},
      {stage1_60[104]}
   );
   gpc1_1 gpc2741 (
      {stage0_60[219]},
      {stage1_60[105]}
   );
   gpc1_1 gpc2742 (
      {stage0_60[220]},
      {stage1_60[106]}
   );
   gpc1_1 gpc2743 (
      {stage0_60[221]},
      {stage1_60[107]}
   );
   gpc1_1 gpc2744 (
      {stage0_60[222]},
      {stage1_60[108]}
   );
   gpc1_1 gpc2745 (
      {stage0_60[223]},
      {stage1_60[109]}
   );
   gpc1_1 gpc2746 (
      {stage0_60[224]},
      {stage1_60[110]}
   );
   gpc1_1 gpc2747 (
      {stage0_60[225]},
      {stage1_60[111]}
   );
   gpc1_1 gpc2748 (
      {stage0_60[226]},
      {stage1_60[112]}
   );
   gpc1_1 gpc2749 (
      {stage0_60[227]},
      {stage1_60[113]}
   );
   gpc1_1 gpc2750 (
      {stage0_60[228]},
      {stage1_60[114]}
   );
   gpc1_1 gpc2751 (
      {stage0_60[229]},
      {stage1_60[115]}
   );
   gpc1_1 gpc2752 (
      {stage0_60[230]},
      {stage1_60[116]}
   );
   gpc1_1 gpc2753 (
      {stage0_60[231]},
      {stage1_60[117]}
   );
   gpc1_1 gpc2754 (
      {stage0_60[232]},
      {stage1_60[118]}
   );
   gpc1_1 gpc2755 (
      {stage0_60[233]},
      {stage1_60[119]}
   );
   gpc1_1 gpc2756 (
      {stage0_60[234]},
      {stage1_60[120]}
   );
   gpc1_1 gpc2757 (
      {stage0_60[235]},
      {stage1_60[121]}
   );
   gpc1_1 gpc2758 (
      {stage0_60[236]},
      {stage1_60[122]}
   );
   gpc1_1 gpc2759 (
      {stage0_60[237]},
      {stage1_60[123]}
   );
   gpc1_1 gpc2760 (
      {stage0_60[238]},
      {stage1_60[124]}
   );
   gpc1_1 gpc2761 (
      {stage0_60[239]},
      {stage1_60[125]}
   );
   gpc1_1 gpc2762 (
      {stage0_60[240]},
      {stage1_60[126]}
   );
   gpc1_1 gpc2763 (
      {stage0_60[241]},
      {stage1_60[127]}
   );
   gpc1_1 gpc2764 (
      {stage0_60[242]},
      {stage1_60[128]}
   );
   gpc1_1 gpc2765 (
      {stage0_60[243]},
      {stage1_60[129]}
   );
   gpc1_1 gpc2766 (
      {stage0_60[244]},
      {stage1_60[130]}
   );
   gpc1_1 gpc2767 (
      {stage0_60[245]},
      {stage1_60[131]}
   );
   gpc1_1 gpc2768 (
      {stage0_60[246]},
      {stage1_60[132]}
   );
   gpc1_1 gpc2769 (
      {stage0_60[247]},
      {stage1_60[133]}
   );
   gpc1_1 gpc2770 (
      {stage0_60[248]},
      {stage1_60[134]}
   );
   gpc1_1 gpc2771 (
      {stage0_60[249]},
      {stage1_60[135]}
   );
   gpc1_1 gpc2772 (
      {stage0_60[250]},
      {stage1_60[136]}
   );
   gpc1_1 gpc2773 (
      {stage0_60[251]},
      {stage1_60[137]}
   );
   gpc1_1 gpc2774 (
      {stage0_60[252]},
      {stage1_60[138]}
   );
   gpc1_1 gpc2775 (
      {stage0_60[253]},
      {stage1_60[139]}
   );
   gpc1_1 gpc2776 (
      {stage0_60[254]},
      {stage1_60[140]}
   );
   gpc1_1 gpc2777 (
      {stage0_60[255]},
      {stage1_60[141]}
   );
   gpc1_1 gpc2778 (
      {stage0_62[133]},
      {stage1_62[78]}
   );
   gpc1_1 gpc2779 (
      {stage0_62[134]},
      {stage1_62[79]}
   );
   gpc1_1 gpc2780 (
      {stage0_62[135]},
      {stage1_62[80]}
   );
   gpc1_1 gpc2781 (
      {stage0_62[136]},
      {stage1_62[81]}
   );
   gpc1_1 gpc2782 (
      {stage0_62[137]},
      {stage1_62[82]}
   );
   gpc1_1 gpc2783 (
      {stage0_62[138]},
      {stage1_62[83]}
   );
   gpc1_1 gpc2784 (
      {stage0_62[139]},
      {stage1_62[84]}
   );
   gpc1_1 gpc2785 (
      {stage0_62[140]},
      {stage1_62[85]}
   );
   gpc1_1 gpc2786 (
      {stage0_62[141]},
      {stage1_62[86]}
   );
   gpc1_1 gpc2787 (
      {stage0_62[142]},
      {stage1_62[87]}
   );
   gpc1_1 gpc2788 (
      {stage0_62[143]},
      {stage1_62[88]}
   );
   gpc1_1 gpc2789 (
      {stage0_62[144]},
      {stage1_62[89]}
   );
   gpc1_1 gpc2790 (
      {stage0_62[145]},
      {stage1_62[90]}
   );
   gpc1_1 gpc2791 (
      {stage0_62[146]},
      {stage1_62[91]}
   );
   gpc1_1 gpc2792 (
      {stage0_62[147]},
      {stage1_62[92]}
   );
   gpc1_1 gpc2793 (
      {stage0_62[148]},
      {stage1_62[93]}
   );
   gpc1_1 gpc2794 (
      {stage0_62[149]},
      {stage1_62[94]}
   );
   gpc1_1 gpc2795 (
      {stage0_62[150]},
      {stage1_62[95]}
   );
   gpc1_1 gpc2796 (
      {stage0_62[151]},
      {stage1_62[96]}
   );
   gpc1_1 gpc2797 (
      {stage0_62[152]},
      {stage1_62[97]}
   );
   gpc1_1 gpc2798 (
      {stage0_62[153]},
      {stage1_62[98]}
   );
   gpc1_1 gpc2799 (
      {stage0_62[154]},
      {stage1_62[99]}
   );
   gpc1_1 gpc2800 (
      {stage0_62[155]},
      {stage1_62[100]}
   );
   gpc1_1 gpc2801 (
      {stage0_62[156]},
      {stage1_62[101]}
   );
   gpc1_1 gpc2802 (
      {stage0_62[157]},
      {stage1_62[102]}
   );
   gpc1_1 gpc2803 (
      {stage0_62[158]},
      {stage1_62[103]}
   );
   gpc1_1 gpc2804 (
      {stage0_62[159]},
      {stage1_62[104]}
   );
   gpc1_1 gpc2805 (
      {stage0_62[160]},
      {stage1_62[105]}
   );
   gpc1_1 gpc2806 (
      {stage0_62[161]},
      {stage1_62[106]}
   );
   gpc1_1 gpc2807 (
      {stage0_62[162]},
      {stage1_62[107]}
   );
   gpc1_1 gpc2808 (
      {stage0_62[163]},
      {stage1_62[108]}
   );
   gpc1_1 gpc2809 (
      {stage0_62[164]},
      {stage1_62[109]}
   );
   gpc1_1 gpc2810 (
      {stage0_62[165]},
      {stage1_62[110]}
   );
   gpc1_1 gpc2811 (
      {stage0_62[166]},
      {stage1_62[111]}
   );
   gpc1_1 gpc2812 (
      {stage0_62[167]},
      {stage1_62[112]}
   );
   gpc1_1 gpc2813 (
      {stage0_62[168]},
      {stage1_62[113]}
   );
   gpc1_1 gpc2814 (
      {stage0_62[169]},
      {stage1_62[114]}
   );
   gpc1_1 gpc2815 (
      {stage0_62[170]},
      {stage1_62[115]}
   );
   gpc1_1 gpc2816 (
      {stage0_62[171]},
      {stage1_62[116]}
   );
   gpc1_1 gpc2817 (
      {stage0_62[172]},
      {stage1_62[117]}
   );
   gpc1_1 gpc2818 (
      {stage0_62[173]},
      {stage1_62[118]}
   );
   gpc1_1 gpc2819 (
      {stage0_62[174]},
      {stage1_62[119]}
   );
   gpc1_1 gpc2820 (
      {stage0_62[175]},
      {stage1_62[120]}
   );
   gpc1_1 gpc2821 (
      {stage0_62[176]},
      {stage1_62[121]}
   );
   gpc1_1 gpc2822 (
      {stage0_62[177]},
      {stage1_62[122]}
   );
   gpc1_1 gpc2823 (
      {stage0_62[178]},
      {stage1_62[123]}
   );
   gpc1_1 gpc2824 (
      {stage0_62[179]},
      {stage1_62[124]}
   );
   gpc1_1 gpc2825 (
      {stage0_62[180]},
      {stage1_62[125]}
   );
   gpc1_1 gpc2826 (
      {stage0_62[181]},
      {stage1_62[126]}
   );
   gpc1_1 gpc2827 (
      {stage0_62[182]},
      {stage1_62[127]}
   );
   gpc1_1 gpc2828 (
      {stage0_62[183]},
      {stage1_62[128]}
   );
   gpc1_1 gpc2829 (
      {stage0_62[184]},
      {stage1_62[129]}
   );
   gpc1_1 gpc2830 (
      {stage0_62[185]},
      {stage1_62[130]}
   );
   gpc1_1 gpc2831 (
      {stage0_62[186]},
      {stage1_62[131]}
   );
   gpc1_1 gpc2832 (
      {stage0_62[187]},
      {stage1_62[132]}
   );
   gpc1_1 gpc2833 (
      {stage0_62[188]},
      {stage1_62[133]}
   );
   gpc1_1 gpc2834 (
      {stage0_62[189]},
      {stage1_62[134]}
   );
   gpc1_1 gpc2835 (
      {stage0_62[190]},
      {stage1_62[135]}
   );
   gpc1_1 gpc2836 (
      {stage0_62[191]},
      {stage1_62[136]}
   );
   gpc1_1 gpc2837 (
      {stage0_62[192]},
      {stage1_62[137]}
   );
   gpc1_1 gpc2838 (
      {stage0_62[193]},
      {stage1_62[138]}
   );
   gpc1_1 gpc2839 (
      {stage0_62[194]},
      {stage1_62[139]}
   );
   gpc1_1 gpc2840 (
      {stage0_62[195]},
      {stage1_62[140]}
   );
   gpc1_1 gpc2841 (
      {stage0_62[196]},
      {stage1_62[141]}
   );
   gpc1_1 gpc2842 (
      {stage0_62[197]},
      {stage1_62[142]}
   );
   gpc1_1 gpc2843 (
      {stage0_62[198]},
      {stage1_62[143]}
   );
   gpc1_1 gpc2844 (
      {stage0_62[199]},
      {stage1_62[144]}
   );
   gpc1_1 gpc2845 (
      {stage0_62[200]},
      {stage1_62[145]}
   );
   gpc1_1 gpc2846 (
      {stage0_62[201]},
      {stage1_62[146]}
   );
   gpc1_1 gpc2847 (
      {stage0_62[202]},
      {stage1_62[147]}
   );
   gpc1_1 gpc2848 (
      {stage0_62[203]},
      {stage1_62[148]}
   );
   gpc1_1 gpc2849 (
      {stage0_62[204]},
      {stage1_62[149]}
   );
   gpc1_1 gpc2850 (
      {stage0_62[205]},
      {stage1_62[150]}
   );
   gpc1_1 gpc2851 (
      {stage0_62[206]},
      {stage1_62[151]}
   );
   gpc1_1 gpc2852 (
      {stage0_62[207]},
      {stage1_62[152]}
   );
   gpc1_1 gpc2853 (
      {stage0_62[208]},
      {stage1_62[153]}
   );
   gpc1_1 gpc2854 (
      {stage0_62[209]},
      {stage1_62[154]}
   );
   gpc1_1 gpc2855 (
      {stage0_62[210]},
      {stage1_62[155]}
   );
   gpc1_1 gpc2856 (
      {stage0_62[211]},
      {stage1_62[156]}
   );
   gpc1_1 gpc2857 (
      {stage0_62[212]},
      {stage1_62[157]}
   );
   gpc1_1 gpc2858 (
      {stage0_62[213]},
      {stage1_62[158]}
   );
   gpc1_1 gpc2859 (
      {stage0_62[214]},
      {stage1_62[159]}
   );
   gpc1_1 gpc2860 (
      {stage0_62[215]},
      {stage1_62[160]}
   );
   gpc1_1 gpc2861 (
      {stage0_62[216]},
      {stage1_62[161]}
   );
   gpc1_1 gpc2862 (
      {stage0_62[217]},
      {stage1_62[162]}
   );
   gpc1_1 gpc2863 (
      {stage0_62[218]},
      {stage1_62[163]}
   );
   gpc1_1 gpc2864 (
      {stage0_62[219]},
      {stage1_62[164]}
   );
   gpc1_1 gpc2865 (
      {stage0_62[220]},
      {stage1_62[165]}
   );
   gpc1_1 gpc2866 (
      {stage0_62[221]},
      {stage1_62[166]}
   );
   gpc1_1 gpc2867 (
      {stage0_62[222]},
      {stage1_62[167]}
   );
   gpc1_1 gpc2868 (
      {stage0_62[223]},
      {stage1_62[168]}
   );
   gpc1_1 gpc2869 (
      {stage0_62[224]},
      {stage1_62[169]}
   );
   gpc1_1 gpc2870 (
      {stage0_62[225]},
      {stage1_62[170]}
   );
   gpc1_1 gpc2871 (
      {stage0_62[226]},
      {stage1_62[171]}
   );
   gpc1_1 gpc2872 (
      {stage0_62[227]},
      {stage1_62[172]}
   );
   gpc1_1 gpc2873 (
      {stage0_62[228]},
      {stage1_62[173]}
   );
   gpc1_1 gpc2874 (
      {stage0_62[229]},
      {stage1_62[174]}
   );
   gpc1_1 gpc2875 (
      {stage0_62[230]},
      {stage1_62[175]}
   );
   gpc1_1 gpc2876 (
      {stage0_62[231]},
      {stage1_62[176]}
   );
   gpc1_1 gpc2877 (
      {stage0_62[232]},
      {stage1_62[177]}
   );
   gpc1_1 gpc2878 (
      {stage0_62[233]},
      {stage1_62[178]}
   );
   gpc1_1 gpc2879 (
      {stage0_62[234]},
      {stage1_62[179]}
   );
   gpc1_1 gpc2880 (
      {stage0_62[235]},
      {stage1_62[180]}
   );
   gpc1_1 gpc2881 (
      {stage0_62[236]},
      {stage1_62[181]}
   );
   gpc1_1 gpc2882 (
      {stage0_62[237]},
      {stage1_62[182]}
   );
   gpc1_1 gpc2883 (
      {stage0_62[238]},
      {stage1_62[183]}
   );
   gpc1_1 gpc2884 (
      {stage0_62[239]},
      {stage1_62[184]}
   );
   gpc1_1 gpc2885 (
      {stage0_62[240]},
      {stage1_62[185]}
   );
   gpc1_1 gpc2886 (
      {stage0_62[241]},
      {stage1_62[186]}
   );
   gpc1_1 gpc2887 (
      {stage0_62[242]},
      {stage1_62[187]}
   );
   gpc1_1 gpc2888 (
      {stage0_62[243]},
      {stage1_62[188]}
   );
   gpc1_1 gpc2889 (
      {stage0_62[244]},
      {stage1_62[189]}
   );
   gpc1_1 gpc2890 (
      {stage0_62[245]},
      {stage1_62[190]}
   );
   gpc1_1 gpc2891 (
      {stage0_62[246]},
      {stage1_62[191]}
   );
   gpc1_1 gpc2892 (
      {stage0_62[247]},
      {stage1_62[192]}
   );
   gpc1_1 gpc2893 (
      {stage0_62[248]},
      {stage1_62[193]}
   );
   gpc1_1 gpc2894 (
      {stage0_62[249]},
      {stage1_62[194]}
   );
   gpc1_1 gpc2895 (
      {stage0_62[250]},
      {stage1_62[195]}
   );
   gpc1_1 gpc2896 (
      {stage0_62[251]},
      {stage1_62[196]}
   );
   gpc1_1 gpc2897 (
      {stage0_62[252]},
      {stage1_62[197]}
   );
   gpc1_1 gpc2898 (
      {stage0_62[253]},
      {stage1_62[198]}
   );
   gpc1_1 gpc2899 (
      {stage0_62[254]},
      {stage1_62[199]}
   );
   gpc1_1 gpc2900 (
      {stage0_62[255]},
      {stage1_62[200]}
   );
   gpc1_1 gpc2901 (
      {stage0_63[252]},
      {stage1_63[65]}
   );
   gpc1_1 gpc2902 (
      {stage0_63[253]},
      {stage1_63[66]}
   );
   gpc1_1 gpc2903 (
      {stage0_63[254]},
      {stage1_63[67]}
   );
   gpc1_1 gpc2904 (
      {stage0_63[255]},
      {stage1_63[68]}
   );
   gpc2135_5 gpc2905 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc2906 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc2907 (
      {stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[2]},
      {stage1_3[4], stage1_3[5]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc2908 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[3]},
      {stage1_3[6], stage1_3[7]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc606_5 gpc2909 (
      {stage1_0[20], stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24], stage1_0[25]},
      {stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc2910 (
      {stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29], stage1_0[30], stage1_0[31]},
      {stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc2911 (
      {stage1_0[32], stage1_0[33], stage1_0[34], stage1_0[35], stage1_0[36], stage1_0[37]},
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc606_5 gpc2912 (
      {stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41], stage1_0[42], stage1_0[43]},
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc606_5 gpc2913 (
      {stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47], stage1_0[48], stage1_0[49]},
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc606_5 gpc2914 (
      {stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53], stage1_0[54], stage1_0[55]},
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc2915 (
      {stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59], stage1_0[60], stage1_0[61]},
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc606_5 gpc2916 (
      {stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65], stage1_0[66], stage1_0[67]},
      {stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc2917 (
      {stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71], stage1_0[72], stage1_0[73]},
      {stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc2918 (
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13]},
      {stage2_5[0],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc2919 (
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19]},
      {stage2_5[1],stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14]}
   );
   gpc606_5 gpc2920 (
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25]},
      {stage2_5[2],stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15]}
   );
   gpc606_5 gpc2921 (
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage2_5[3],stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16]}
   );
   gpc606_5 gpc2922 (
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37]},
      {stage2_5[4],stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17]}
   );
   gpc606_5 gpc2923 (
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage2_5[5],stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18]}
   );
   gpc606_5 gpc2924 (
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49]},
      {stage2_5[6],stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19]}
   );
   gpc615_5 gpc2925 (
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58]},
      {stage1_2[58]},
      {stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage2_5[7],stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20]}
   );
   gpc615_5 gpc2926 (
      {stage1_1[59], stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63]},
      {stage1_2[59]},
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61]},
      {stage2_5[8],stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21]}
   );
   gpc615_5 gpc2927 (
      {stage1_1[64], stage1_1[65], stage1_1[66], stage1_1[67], stage1_1[68]},
      {stage1_2[60]},
      {stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66], stage1_3[67]},
      {stage2_5[9],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc615_5 gpc2928 (
      {stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage1_3[68]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[10],stage2_4[23],stage2_3[23],stage2_2[23]}
   );
   gpc615_5 gpc2929 (
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70]},
      {stage1_3[69]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[11],stage2_4[24],stage2_3[24],stage2_2[24]}
   );
   gpc615_5 gpc2930 (
      {stage1_2[71], stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75]},
      {stage1_3[70]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[12],stage2_4[25],stage2_3[25],stage2_2[25]}
   );
   gpc615_5 gpc2931 (
      {stage1_2[76], stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80]},
      {stage1_3[71]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[13],stage2_4[26],stage2_3[26],stage2_2[26]}
   );
   gpc615_5 gpc2932 (
      {stage1_2[81], stage1_2[82], stage1_2[83], stage1_2[84], stage1_2[85]},
      {stage1_3[72]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[14],stage2_4[27],stage2_3[27],stage2_2[27]}
   );
   gpc615_5 gpc2933 (
      {stage1_2[86], stage1_2[87], stage1_2[88], stage1_2[89], stage1_2[90]},
      {stage1_3[73]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[15],stage2_4[28],stage2_3[28],stage2_2[28]}
   );
   gpc615_5 gpc2934 (
      {stage1_2[91], stage1_2[92], stage1_2[93], stage1_2[94], stage1_2[95]},
      {stage1_3[74]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[16],stage2_4[29],stage2_3[29],stage2_2[29]}
   );
   gpc615_5 gpc2935 (
      {stage1_2[96], stage1_2[97], stage1_2[98], stage1_2[99], stage1_2[100]},
      {stage1_3[75]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[17],stage2_4[30],stage2_3[30],stage2_2[30]}
   );
   gpc615_5 gpc2936 (
      {stage1_2[101], stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105]},
      {stage1_3[76]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[18],stage2_4[31],stage2_3[31],stage2_2[31]}
   );
   gpc615_5 gpc2937 (
      {stage1_2[106], stage1_2[107], stage1_2[108], stage1_2[109], stage1_2[110]},
      {stage1_3[77]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[19],stage2_4[32],stage2_3[32],stage2_2[32]}
   );
   gpc615_5 gpc2938 (
      {stage1_2[111], stage1_2[112], stage1_2[113], stage1_2[114], stage1_2[115]},
      {stage1_3[78]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[20],stage2_4[33],stage2_3[33],stage2_2[33]}
   );
   gpc615_5 gpc2939 (
      {stage1_2[116], stage1_2[117], stage1_2[118], stage1_2[119], stage1_2[120]},
      {stage1_3[79]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[21],stage2_4[34],stage2_3[34],stage2_2[34]}
   );
   gpc615_5 gpc2940 (
      {stage1_2[121], stage1_2[122], stage1_2[123], stage1_2[124], stage1_2[125]},
      {stage1_3[80]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[22],stage2_4[35],stage2_3[35],stage2_2[35]}
   );
   gpc615_5 gpc2941 (
      {stage1_2[126], stage1_2[127], stage1_2[128], stage1_2[129], stage1_2[130]},
      {stage1_3[81]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[23],stage2_4[36],stage2_3[36],stage2_2[36]}
   );
   gpc615_5 gpc2942 (
      {stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86]},
      {stage1_4[84]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[14],stage2_5[24],stage2_4[37],stage2_3[37]}
   );
   gpc615_5 gpc2943 (
      {stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90], stage1_3[91]},
      {stage1_4[85]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[15],stage2_5[25],stage2_4[38],stage2_3[38]}
   );
   gpc606_5 gpc2944 (
      {stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[2],stage2_6[16],stage2_5[26],stage2_4[39]}
   );
   gpc606_5 gpc2945 (
      {stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96], stage1_4[97]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[3],stage2_6[17],stage2_5[27],stage2_4[40]}
   );
   gpc606_5 gpc2946 (
      {stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101], stage1_4[102], stage1_4[103]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[4],stage2_6[18],stage2_5[28],stage2_4[41]}
   );
   gpc606_5 gpc2947 (
      {stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107], stage1_4[108], stage1_4[109]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[5],stage2_6[19],stage2_5[29],stage2_4[42]}
   );
   gpc606_5 gpc2948 (
      {stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[6],stage2_6[20],stage2_5[30],stage2_4[43]}
   );
   gpc606_5 gpc2949 (
      {stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[7],stage2_6[21],stage2_5[31],stage2_4[44]}
   );
   gpc606_5 gpc2950 (
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[6],stage2_7[8],stage2_6[22],stage2_5[32]}
   );
   gpc606_5 gpc2951 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[7],stage2_7[9],stage2_6[23],stage2_5[33]}
   );
   gpc606_5 gpc2952 (
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[8],stage2_7[10],stage2_6[24],stage2_5[34]}
   );
   gpc606_5 gpc2953 (
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[9],stage2_7[11],stage2_6[25],stage2_5[35]}
   );
   gpc606_5 gpc2954 (
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[10],stage2_7[12],stage2_6[26],stage2_5[36]}
   );
   gpc606_5 gpc2955 (
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[11],stage2_7[13],stage2_6[27],stage2_5[37]}
   );
   gpc606_5 gpc2956 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[12],stage2_7[14],stage2_6[28],stage2_5[38]}
   );
   gpc606_5 gpc2957 (
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[13],stage2_7[15],stage2_6[29],stage2_5[39]}
   );
   gpc606_5 gpc2958 (
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[14],stage2_7[16],stage2_6[30],stage2_5[40]}
   );
   gpc606_5 gpc2959 (
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[15],stage2_7[17],stage2_6[31],stage2_5[41]}
   );
   gpc606_5 gpc2960 (
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[16],stage2_7[18],stage2_6[32],stage2_5[42]}
   );
   gpc606_5 gpc2961 (
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[17],stage2_7[19],stage2_6[33],stage2_5[43]}
   );
   gpc606_5 gpc2962 (
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77]},
      {stage2_9[12],stage2_8[18],stage2_7[20],stage2_6[34],stage2_5[44]}
   );
   gpc606_5 gpc2963 (
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83]},
      {stage2_9[13],stage2_8[19],stage2_7[21],stage2_6[35],stage2_5[45]}
   );
   gpc615_5 gpc2964 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40]},
      {stage1_7[84]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[14],stage2_8[20],stage2_7[22],stage2_6[36]}
   );
   gpc615_5 gpc2965 (
      {stage1_6[41], stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45]},
      {stage1_7[85]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[15],stage2_8[21],stage2_7[23],stage2_6[37]}
   );
   gpc615_5 gpc2966 (
      {stage1_6[46], stage1_6[47], stage1_6[48], stage1_6[49], stage1_6[50]},
      {stage1_7[86]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[16],stage2_8[22],stage2_7[24],stage2_6[38]}
   );
   gpc615_5 gpc2967 (
      {stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54], stage1_6[55]},
      {stage1_7[87]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[17],stage2_8[23],stage2_7[25],stage2_6[39]}
   );
   gpc615_5 gpc2968 (
      {stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage1_7[88]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[18],stage2_8[24],stage2_7[26],stage2_6[40]}
   );
   gpc615_5 gpc2969 (
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage1_7[89]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[19],stage2_8[25],stage2_7[27],stage2_6[41]}
   );
   gpc615_5 gpc2970 (
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70]},
      {stage1_7[90]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[20],stage2_8[26],stage2_7[28],stage2_6[42]}
   );
   gpc615_5 gpc2971 (
      {stage1_6[71], stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75]},
      {stage1_7[91]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[21],stage2_8[27],stage2_7[29],stage2_6[43]}
   );
   gpc615_5 gpc2972 (
      {stage1_6[76], stage1_6[77], stage1_6[78], stage1_6[79], stage1_6[80]},
      {stage1_7[92]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[22],stage2_8[28],stage2_7[30],stage2_6[44]}
   );
   gpc615_5 gpc2973 (
      {stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84], stage1_6[85]},
      {stage1_7[93]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[23],stage2_8[29],stage2_7[31],stage2_6[45]}
   );
   gpc615_5 gpc2974 (
      {stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage1_7[94]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[24],stage2_8[30],stage2_7[32],stage2_6[46]}
   );
   gpc615_5 gpc2975 (
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_7[95]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[25],stage2_8[31],stage2_7[33],stage2_6[47]}
   );
   gpc615_5 gpc2976 (
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100]},
      {stage1_7[96]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[26],stage2_8[32],stage2_7[34],stage2_6[48]}
   );
   gpc615_5 gpc2977 (
      {stage1_6[101], stage1_6[102], stage1_6[103], stage1_6[104], stage1_6[105]},
      {stage1_7[97]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[27],stage2_8[33],stage2_7[35],stage2_6[49]}
   );
   gpc615_5 gpc2978 (
      {stage1_6[106], stage1_6[107], stage1_6[108], stage1_6[109], stage1_6[110]},
      {stage1_7[98]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[28],stage2_8[34],stage2_7[36],stage2_6[50]}
   );
   gpc615_5 gpc2979 (
      {stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114], stage1_6[115]},
      {stage1_7[99]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[29],stage2_8[35],stage2_7[37],stage2_6[51]}
   );
   gpc606_5 gpc2980 (
      {stage1_7[100], stage1_7[101], stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[16],stage2_9[30],stage2_8[36],stage2_7[38]}
   );
   gpc606_5 gpc2981 (
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[17],stage2_9[31],stage2_8[37]}
   );
   gpc606_5 gpc2982 (
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[2],stage2_10[18],stage2_9[32],stage2_8[38]}
   );
   gpc606_5 gpc2983 (
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[3],stage2_10[19],stage2_9[33],stage2_8[39]}
   );
   gpc606_5 gpc2984 (
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[4],stage2_10[20],stage2_9[34],stage2_8[40]}
   );
   gpc606_5 gpc2985 (
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[5],stage2_10[21],stage2_9[35],stage2_8[41]}
   );
   gpc606_5 gpc2986 (
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[6],stage2_10[22],stage2_9[36],stage2_8[42]}
   );
   gpc615_5 gpc2987 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10]},
      {stage1_10[36]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[6],stage2_11[7],stage2_10[23],stage2_9[37]}
   );
   gpc615_5 gpc2988 (
      {stage1_9[11], stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15]},
      {stage1_10[37]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[7],stage2_11[8],stage2_10[24],stage2_9[38]}
   );
   gpc615_5 gpc2989 (
      {stage1_9[16], stage1_9[17], stage1_9[18], stage1_9[19], stage1_9[20]},
      {stage1_10[38]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[8],stage2_11[9],stage2_10[25],stage2_9[39]}
   );
   gpc615_5 gpc2990 (
      {stage1_9[21], stage1_9[22], stage1_9[23], stage1_9[24], stage1_9[25]},
      {stage1_10[39]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[9],stage2_11[10],stage2_10[26],stage2_9[40]}
   );
   gpc615_5 gpc2991 (
      {stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29], stage1_9[30]},
      {stage1_10[40]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[10],stage2_11[11],stage2_10[27],stage2_9[41]}
   );
   gpc615_5 gpc2992 (
      {stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_10[41]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[11],stage2_11[12],stage2_10[28],stage2_9[42]}
   );
   gpc615_5 gpc2993 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40]},
      {stage1_10[42]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[12],stage2_11[13],stage2_10[29],stage2_9[43]}
   );
   gpc615_5 gpc2994 (
      {stage1_9[41], stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45]},
      {stage1_10[43]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[13],stage2_11[14],stage2_10[30],stage2_9[44]}
   );
   gpc615_5 gpc2995 (
      {stage1_9[46], stage1_9[47], stage1_9[48], stage1_9[49], stage1_9[50]},
      {stage1_10[44]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[14],stage2_11[15],stage2_10[31],stage2_9[45]}
   );
   gpc615_5 gpc2996 (
      {stage1_9[51], stage1_9[52], stage1_9[53], stage1_9[54], stage1_9[55]},
      {stage1_10[45]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[15],stage2_11[16],stage2_10[32],stage2_9[46]}
   );
   gpc615_5 gpc2997 (
      {stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59], stage1_9[60]},
      {stage1_10[46]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[16],stage2_11[17],stage2_10[33],stage2_9[47]}
   );
   gpc615_5 gpc2998 (
      {stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage1_10[47]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[17],stage2_11[18],stage2_10[34],stage2_9[48]}
   );
   gpc615_5 gpc2999 (
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70]},
      {stage1_10[48]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[18],stage2_11[19],stage2_10[35],stage2_9[49]}
   );
   gpc615_5 gpc3000 (
      {stage1_9[71], stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75]},
      {stage1_10[49]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[19],stage2_11[20],stage2_10[36],stage2_9[50]}
   );
   gpc615_5 gpc3001 (
      {stage1_9[76], stage1_9[77], stage1_9[78], stage1_9[79], stage1_9[80]},
      {stage1_10[50]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[20],stage2_11[21],stage2_10[37],stage2_9[51]}
   );
   gpc615_5 gpc3002 (
      {stage1_9[81], stage1_9[82], stage1_9[83], stage1_9[84], stage1_9[85]},
      {stage1_10[51]},
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95]},
      {stage2_13[15],stage2_12[21],stage2_11[22],stage2_10[38],stage2_9[52]}
   );
   gpc615_5 gpc3003 (
      {stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89], stage1_9[90]},
      {stage1_10[52]},
      {stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage2_13[16],stage2_12[22],stage2_11[23],stage2_10[39],stage2_9[53]}
   );
   gpc615_5 gpc3004 (
      {stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage1_10[53]},
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107]},
      {stage2_13[17],stage2_12[23],stage2_11[24],stage2_10[40],stage2_9[54]}
   );
   gpc615_5 gpc3005 (
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100]},
      {stage1_10[54]},
      {stage1_11[108], stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113]},
      {stage2_13[18],stage2_12[24],stage2_11[25],stage2_10[41],stage2_9[55]}
   );
   gpc615_5 gpc3006 (
      {stage1_9[101], stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105]},
      {stage1_10[55]},
      {stage1_11[114], stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119]},
      {stage2_13[19],stage2_12[25],stage2_11[26],stage2_10[42],stage2_9[56]}
   );
   gpc615_5 gpc3007 (
      {stage1_9[106], stage1_9[107], stage1_9[108], stage1_9[109], stage1_9[110]},
      {stage1_10[56]},
      {stage1_11[120], stage1_11[121], stage1_11[122], stage1_11[123], stage1_11[124], stage1_11[125]},
      {stage2_13[20],stage2_12[26],stage2_11[27],stage2_10[43],stage2_9[57]}
   );
   gpc615_5 gpc3008 (
      {stage1_9[111], stage1_9[112], stage1_9[113], stage1_9[114], stage1_9[115]},
      {stage1_10[57]},
      {stage1_11[126], stage1_11[127], stage1_11[128], stage1_11[129], stage1_11[130], stage1_11[131]},
      {stage2_13[21],stage2_12[27],stage2_11[28],stage2_10[44],stage2_9[58]}
   );
   gpc615_5 gpc3009 (
      {stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119], 1'b0},
      {stage1_10[58]},
      {stage1_11[132], stage1_11[133], stage1_11[134], stage1_11[135], stage1_11[136], stage1_11[137]},
      {stage2_13[22],stage2_12[28],stage2_11[29],stage2_10[45],stage2_9[59]}
   );
   gpc606_5 gpc3010 (
      {stage1_10[59], stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[23],stage2_12[29],stage2_11[30],stage2_10[46]}
   );
   gpc606_5 gpc3011 (
      {stage1_10[65], stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[24],stage2_12[30],stage2_11[31],stage2_10[47]}
   );
   gpc606_5 gpc3012 (
      {stage1_10[71], stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[25],stage2_12[31],stage2_11[32],stage2_10[48]}
   );
   gpc606_5 gpc3013 (
      {stage1_10[77], stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[26],stage2_12[32],stage2_11[33],stage2_10[49]}
   );
   gpc606_5 gpc3014 (
      {stage1_10[83], stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[27],stage2_12[33],stage2_11[34],stage2_10[50]}
   );
   gpc606_5 gpc3015 (
      {stage1_10[89], stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[28],stage2_12[34],stage2_11[35],stage2_10[51]}
   );
   gpc606_5 gpc3016 (
      {stage1_10[95], stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[29],stage2_12[35],stage2_11[36],stage2_10[52]}
   );
   gpc606_5 gpc3017 (
      {stage1_10[101], stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[30],stage2_12[36],stage2_11[37],stage2_10[53]}
   );
   gpc606_5 gpc3018 (
      {stage1_10[107], stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[31],stage2_12[37],stage2_11[38],stage2_10[54]}
   );
   gpc606_5 gpc3019 (
      {stage1_10[113], stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[32],stage2_12[38],stage2_11[39],stage2_10[55]}
   );
   gpc606_5 gpc3020 (
      {stage1_10[119], stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[33],stage2_12[39],stage2_11[40],stage2_10[56]}
   );
   gpc606_5 gpc3021 (
      {stage1_10[125], stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[34],stage2_12[40],stage2_11[41],stage2_10[57]}
   );
   gpc606_5 gpc3022 (
      {stage1_10[131], stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[35],stage2_12[41],stage2_11[42],stage2_10[58]}
   );
   gpc615_5 gpc3023 (
      {stage1_10[137], stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141]},
      {stage1_11[138]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[36],stage2_12[42],stage2_11[43],stage2_10[59]}
   );
   gpc615_5 gpc3024 (
      {stage1_10[142], stage1_10[143], stage1_10[144], stage1_10[145], stage1_10[146]},
      {stage1_11[139]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[37],stage2_12[43],stage2_11[44],stage2_10[60]}
   );
   gpc1406_5 gpc3025 (
      {stage1_11[140], stage1_11[141], stage1_11[142], stage1_11[143], stage1_11[144], stage1_11[145]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[15],stage2_13[38],stage2_12[44],stage2_11[45]}
   );
   gpc606_5 gpc3026 (
      {stage1_11[146], stage1_11[147], stage1_11[148], stage1_11[149], stage1_11[150], stage1_11[151]},
      {stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9]},
      {stage2_15[1],stage2_14[16],stage2_13[39],stage2_12[45],stage2_11[46]}
   );
   gpc606_5 gpc3027 (
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[0],stage2_15[2],stage2_14[17],stage2_13[40],stage2_12[46]}
   );
   gpc606_5 gpc3028 (
      {stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage2_16[1],stage2_15[3],stage2_14[18],stage2_13[41],stage2_12[47]}
   );
   gpc606_5 gpc3029 (
      {stage1_12[102], stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107]},
      {stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18]},
      {stage2_16[2],stage2_15[4],stage2_14[19],stage2_13[42],stage2_12[48]}
   );
   gpc606_5 gpc3030 (
      {stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113]},
      {stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24]},
      {stage2_16[3],stage2_15[5],stage2_14[20],stage2_13[43],stage2_12[49]}
   );
   gpc606_5 gpc3031 (
      {stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30]},
      {stage2_16[4],stage2_15[6],stage2_14[21],stage2_13[44],stage2_12[50]}
   );
   gpc606_5 gpc3032 (
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125]},
      {stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36]},
      {stage2_16[5],stage2_15[7],stage2_14[22],stage2_13[45],stage2_12[51]}
   );
   gpc606_5 gpc3033 (
      {stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131]},
      {stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42]},
      {stage2_16[6],stage2_15[8],stage2_14[23],stage2_13[46],stage2_12[52]}
   );
   gpc606_5 gpc3034 (
      {stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[7],stage2_15[9],stage2_14[24],stage2_13[47]}
   );
   gpc606_5 gpc3035 (
      {stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[8],stage2_15[10],stage2_14[25],stage2_13[48]}
   );
   gpc606_5 gpc3036 (
      {stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[9],stage2_15[11],stage2_14[26],stage2_13[49]}
   );
   gpc606_5 gpc3037 (
      {stage1_13[28], stage1_13[29], stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[10],stage2_15[12],stage2_14[27],stage2_13[50]}
   );
   gpc606_5 gpc3038 (
      {stage1_13[34], stage1_13[35], stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[11],stage2_15[13],stage2_14[28],stage2_13[51]}
   );
   gpc606_5 gpc3039 (
      {stage1_13[40], stage1_13[41], stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[12],stage2_15[14],stage2_14[29],stage2_13[52]}
   );
   gpc606_5 gpc3040 (
      {stage1_13[46], stage1_13[47], stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[13],stage2_15[15],stage2_14[30],stage2_13[53]}
   );
   gpc606_5 gpc3041 (
      {stage1_13[52], stage1_13[53], stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[14],stage2_15[16],stage2_14[31],stage2_13[54]}
   );
   gpc606_5 gpc3042 (
      {stage1_13[58], stage1_13[59], stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage2_17[8],stage2_16[15],stage2_15[17],stage2_14[32],stage2_13[55]}
   );
   gpc606_5 gpc3043 (
      {stage1_13[64], stage1_13[65], stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage2_17[9],stage2_16[16],stage2_15[18],stage2_14[33],stage2_13[56]}
   );
   gpc606_5 gpc3044 (
      {stage1_13[70], stage1_13[71], stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage2_17[10],stage2_16[17],stage2_15[19],stage2_14[34],stage2_13[57]}
   );
   gpc606_5 gpc3045 (
      {stage1_13[76], stage1_13[77], stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage2_17[11],stage2_16[18],stage2_15[20],stage2_14[35],stage2_13[58]}
   );
   gpc606_5 gpc3046 (
      {stage1_13[82], stage1_13[83], stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage2_17[12],stage2_16[19],stage2_15[21],stage2_14[36],stage2_13[59]}
   );
   gpc606_5 gpc3047 (
      {stage1_13[88], stage1_13[89], stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage2_17[13],stage2_16[20],stage2_15[22],stage2_14[37],stage2_13[60]}
   );
   gpc606_5 gpc3048 (
      {stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[14],stage2_16[21],stage2_15[23],stage2_14[38]}
   );
   gpc606_5 gpc3049 (
      {stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[15],stage2_16[22],stage2_15[24],stage2_14[39]}
   );
   gpc606_5 gpc3050 (
      {stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59], stage1_14[60]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[16],stage2_16[23],stage2_15[25],stage2_14[40]}
   );
   gpc606_5 gpc3051 (
      {stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65], stage1_14[66]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[17],stage2_16[24],stage2_15[26],stage2_14[41]}
   );
   gpc606_5 gpc3052 (
      {stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71], stage1_14[72]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[18],stage2_16[25],stage2_15[27],stage2_14[42]}
   );
   gpc606_5 gpc3053 (
      {stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77], stage1_14[78]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[19],stage2_16[26],stage2_15[28],stage2_14[43]}
   );
   gpc606_5 gpc3054 (
      {stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83], stage1_14[84]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[20],stage2_16[27],stage2_15[29],stage2_14[44]}
   );
   gpc615_5 gpc3055 (
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88]},
      {stage1_16[42]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[7],stage2_17[21],stage2_16[28],stage2_15[30]}
   );
   gpc207_4 gpc3056 (
      {stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49]},
      {stage1_18[0], stage1_18[1]},
      {stage2_19[1],stage2_18[8],stage2_17[22],stage2_16[29]}
   );
   gpc606_5 gpc3057 (
      {stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53], stage1_16[54], stage1_16[55]},
      {stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5], stage1_18[6], stage1_18[7]},
      {stage2_20[0],stage2_19[2],stage2_18[9],stage2_17[23],stage2_16[30]}
   );
   gpc606_5 gpc3058 (
      {stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59], stage1_16[60], stage1_16[61]},
      {stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11], stage1_18[12], stage1_18[13]},
      {stage2_20[1],stage2_19[3],stage2_18[10],stage2_17[24],stage2_16[31]}
   );
   gpc606_5 gpc3059 (
      {stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65], stage1_16[66], stage1_16[67]},
      {stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17], stage1_18[18], stage1_18[19]},
      {stage2_20[2],stage2_19[4],stage2_18[11],stage2_17[25],stage2_16[32]}
   );
   gpc606_5 gpc3060 (
      {stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73]},
      {stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23], stage1_18[24], stage1_18[25]},
      {stage2_20[3],stage2_19[5],stage2_18[12],stage2_17[26],stage2_16[33]}
   );
   gpc606_5 gpc3061 (
      {stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79]},
      {stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29], stage1_18[30], stage1_18[31]},
      {stage2_20[4],stage2_19[6],stage2_18[13],stage2_17[27],stage2_16[34]}
   );
   gpc606_5 gpc3062 (
      {stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83], stage1_16[84], stage1_16[85]},
      {stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35], stage1_18[36], stage1_18[37]},
      {stage2_20[5],stage2_19[7],stage2_18[14],stage2_17[28],stage2_16[35]}
   );
   gpc606_5 gpc3063 (
      {stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89], stage1_16[90], stage1_16[91]},
      {stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41], stage1_18[42], stage1_18[43]},
      {stage2_20[6],stage2_19[8],stage2_18[15],stage2_17[29],stage2_16[36]}
   );
   gpc606_5 gpc3064 (
      {stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95], stage1_16[96], stage1_16[97]},
      {stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47], stage1_18[48], stage1_18[49]},
      {stage2_20[7],stage2_19[9],stage2_18[16],stage2_17[30],stage2_16[37]}
   );
   gpc606_5 gpc3065 (
      {stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101], stage1_16[102], stage1_16[103]},
      {stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53], stage1_18[54], stage1_18[55]},
      {stage2_20[8],stage2_19[10],stage2_18[17],stage2_17[31],stage2_16[38]}
   );
   gpc606_5 gpc3066 (
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[9],stage2_19[11],stage2_18[18],stage2_17[32]}
   );
   gpc606_5 gpc3067 (
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[10],stage2_19[12],stage2_18[19],stage2_17[33]}
   );
   gpc606_5 gpc3068 (
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[11],stage2_19[13],stage2_18[20],stage2_17[34]}
   );
   gpc606_5 gpc3069 (
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[12],stage2_19[14],stage2_18[21],stage2_17[35]}
   );
   gpc606_5 gpc3070 (
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[13],stage2_19[15],stage2_18[22],stage2_17[36]}
   );
   gpc606_5 gpc3071 (
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[14],stage2_19[16],stage2_18[23],stage2_17[37]}
   );
   gpc606_5 gpc3072 (
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[15],stage2_19[17],stage2_18[24],stage2_17[38]}
   );
   gpc606_5 gpc3073 (
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[16],stage2_19[18],stage2_18[25],stage2_17[39]}
   );
   gpc606_5 gpc3074 (
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[17],stage2_19[19],stage2_18[26],stage2_17[40]}
   );
   gpc606_5 gpc3075 (
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[18],stage2_19[20],stage2_18[27],stage2_17[41]}
   );
   gpc606_5 gpc3076 (
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[19],stage2_19[21],stage2_18[28],stage2_17[42]}
   );
   gpc606_5 gpc3077 (
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[20],stage2_19[22],stage2_18[29],stage2_17[43]}
   );
   gpc606_5 gpc3078 (
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage1_19[72], stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage2_21[12],stage2_20[21],stage2_19[23],stage2_18[30],stage2_17[44]}
   );
   gpc606_5 gpc3079 (
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82], stage1_19[83]},
      {stage2_21[13],stage2_20[22],stage2_19[24],stage2_18[31],stage2_17[45]}
   );
   gpc606_5 gpc3080 (
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87], stage1_19[88], stage1_19[89]},
      {stage2_21[14],stage2_20[23],stage2_19[25],stage2_18[32],stage2_17[46]}
   );
   gpc606_5 gpc3081 (
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93], stage1_19[94], stage1_19[95]},
      {stage2_21[15],stage2_20[24],stage2_19[26],stage2_18[33],stage2_17[47]}
   );
   gpc615_5 gpc3082 (
      {stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59], stage1_18[60]},
      {stage1_19[96]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[16],stage2_20[25],stage2_19[27],stage2_18[34]}
   );
   gpc615_5 gpc3083 (
      {stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage1_19[97]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[17],stage2_20[26],stage2_19[28],stage2_18[35]}
   );
   gpc615_5 gpc3084 (
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70]},
      {stage1_19[98]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[18],stage2_20[27],stage2_19[29],stage2_18[36]}
   );
   gpc615_5 gpc3085 (
      {stage1_19[99], stage1_19[100], stage1_19[101], stage1_19[102], stage1_19[103]},
      {stage1_20[18]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[3],stage2_21[19],stage2_20[28],stage2_19[30]}
   );
   gpc615_5 gpc3086 (
      {stage1_19[104], stage1_19[105], stage1_19[106], stage1_19[107], stage1_19[108]},
      {stage1_20[19]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[4],stage2_21[20],stage2_20[29],stage2_19[31]}
   );
   gpc615_5 gpc3087 (
      {stage1_19[109], stage1_19[110], stage1_19[111], stage1_19[112], stage1_19[113]},
      {stage1_20[20]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[5],stage2_21[21],stage2_20[30],stage2_19[32]}
   );
   gpc615_5 gpc3088 (
      {stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117], stage1_19[118]},
      {stage1_20[21]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[6],stage2_21[22],stage2_20[31],stage2_19[33]}
   );
   gpc615_5 gpc3089 (
      {stage1_19[119], stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123]},
      {stage1_20[22]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[7],stage2_21[23],stage2_20[32],stage2_19[34]}
   );
   gpc606_5 gpc3090 (
      {stage1_20[23], stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[5],stage2_22[8],stage2_21[24],stage2_20[33]}
   );
   gpc606_5 gpc3091 (
      {stage1_20[29], stage1_20[30], stage1_20[31], stage1_20[32], stage1_20[33], stage1_20[34]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[6],stage2_22[9],stage2_21[25],stage2_20[34]}
   );
   gpc606_5 gpc3092 (
      {stage1_20[35], stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39], stage1_20[40]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[7],stage2_22[10],stage2_21[26],stage2_20[35]}
   );
   gpc606_5 gpc3093 (
      {stage1_20[41], stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[8],stage2_22[11],stage2_21[27],stage2_20[36]}
   );
   gpc606_5 gpc3094 (
      {stage1_20[47], stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51], stage1_20[52]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[9],stage2_22[12],stage2_21[28],stage2_20[37]}
   );
   gpc606_5 gpc3095 (
      {stage1_20[53], stage1_20[54], stage1_20[55], stage1_20[56], stage1_20[57], stage1_20[58]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[10],stage2_22[13],stage2_21[29],stage2_20[38]}
   );
   gpc606_5 gpc3096 (
      {stage1_20[59], stage1_20[60], stage1_20[61], stage1_20[62], stage1_20[63], stage1_20[64]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[11],stage2_22[14],stage2_21[30],stage2_20[39]}
   );
   gpc606_5 gpc3097 (
      {stage1_20[65], stage1_20[66], stage1_20[67], stage1_20[68], stage1_20[69], stage1_20[70]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[12],stage2_22[15],stage2_21[31],stage2_20[40]}
   );
   gpc606_5 gpc3098 (
      {stage1_20[71], stage1_20[72], stage1_20[73], stage1_20[74], stage1_20[75], stage1_20[76]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[13],stage2_22[16],stage2_21[32],stage2_20[41]}
   );
   gpc606_5 gpc3099 (
      {stage1_20[77], stage1_20[78], stage1_20[79], stage1_20[80], stage1_20[81], stage1_20[82]},
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage2_24[9],stage2_23[14],stage2_22[17],stage2_21[33],stage2_20[42]}
   );
   gpc606_5 gpc3100 (
      {stage1_20[83], stage1_20[84], stage1_20[85], stage1_20[86], stage1_20[87], stage1_20[88]},
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage2_24[10],stage2_23[15],stage2_22[18],stage2_21[34],stage2_20[43]}
   );
   gpc606_5 gpc3101 (
      {stage1_20[89], stage1_20[90], stage1_20[91], stage1_20[92], stage1_20[93], stage1_20[94]},
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage2_24[11],stage2_23[16],stage2_22[19],stage2_21[35],stage2_20[44]}
   );
   gpc606_5 gpc3102 (
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[12],stage2_23[17],stage2_22[20],stage2_21[36]}
   );
   gpc606_5 gpc3103 (
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[13],stage2_23[18],stage2_22[21],stage2_21[37]}
   );
   gpc606_5 gpc3104 (
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[14],stage2_23[19],stage2_22[22],stage2_21[38]}
   );
   gpc606_5 gpc3105 (
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[15],stage2_23[20],stage2_22[23],stage2_21[39]}
   );
   gpc606_5 gpc3106 (
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[16],stage2_23[21],stage2_22[24],stage2_21[40]}
   );
   gpc606_5 gpc3107 (
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage2_25[5],stage2_24[17],stage2_23[22],stage2_22[25],stage2_21[41]}
   );
   gpc606_5 gpc3108 (
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage2_25[6],stage2_24[18],stage2_23[23],stage2_22[26],stage2_21[42]}
   );
   gpc606_5 gpc3109 (
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage2_25[7],stage2_24[19],stage2_23[24],stage2_22[27],stage2_21[43]}
   );
   gpc606_5 gpc3110 (
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage2_25[8],stage2_24[20],stage2_23[25],stage2_22[28],stage2_21[44]}
   );
   gpc606_5 gpc3111 (
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage2_25[9],stage2_24[21],stage2_23[26],stage2_22[29],stage2_21[45]}
   );
   gpc606_5 gpc3112 (
      {stage1_21[90], stage1_21[91], stage1_21[92], stage1_21[93], stage1_21[94], stage1_21[95]},
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage2_25[10],stage2_24[22],stage2_23[27],stage2_22[30],stage2_21[46]}
   );
   gpc606_5 gpc3113 (
      {stage1_21[96], stage1_21[97], stage1_21[98], stage1_21[99], stage1_21[100], stage1_21[101]},
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage2_25[11],stage2_24[23],stage2_23[28],stage2_22[31],stage2_21[47]}
   );
   gpc606_5 gpc3114 (
      {stage1_21[102], stage1_21[103], stage1_21[104], stage1_21[105], stage1_21[106], stage1_21[107]},
      {stage1_23[72], stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage2_25[12],stage2_24[24],stage2_23[29],stage2_22[32],stage2_21[48]}
   );
   gpc615_5 gpc3115 (
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76]},
      {stage1_23[78]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[13],stage2_24[25],stage2_23[30],stage2_22[33]}
   );
   gpc615_5 gpc3116 (
      {stage1_22[77], stage1_22[78], stage1_22[79], stage1_22[80], stage1_22[81]},
      {stage1_23[79]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[14],stage2_24[26],stage2_23[31],stage2_22[34]}
   );
   gpc615_5 gpc3117 (
      {stage1_22[82], stage1_22[83], stage1_22[84], stage1_22[85], stage1_22[86]},
      {stage1_23[80]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[15],stage2_24[27],stage2_23[32],stage2_22[35]}
   );
   gpc615_5 gpc3118 (
      {stage1_23[81], stage1_23[82], stage1_23[83], stage1_23[84], stage1_23[85]},
      {stage1_24[18]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[3],stage2_25[16],stage2_24[28],stage2_23[33]}
   );
   gpc615_5 gpc3119 (
      {stage1_23[86], stage1_23[87], stage1_23[88], stage1_23[89], stage1_23[90]},
      {stage1_24[19]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[4],stage2_25[17],stage2_24[29],stage2_23[34]}
   );
   gpc615_5 gpc3120 (
      {stage1_23[91], stage1_23[92], stage1_23[93], stage1_23[94], stage1_23[95]},
      {stage1_24[20]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[5],stage2_25[18],stage2_24[30],stage2_23[35]}
   );
   gpc615_5 gpc3121 (
      {stage1_23[96], stage1_23[97], stage1_23[98], stage1_23[99], stage1_23[100]},
      {stage1_24[21]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[6],stage2_25[19],stage2_24[31],stage2_23[36]}
   );
   gpc615_5 gpc3122 (
      {stage1_23[101], stage1_23[102], stage1_23[103], stage1_23[104], stage1_23[105]},
      {stage1_24[22]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[7],stage2_25[20],stage2_24[32],stage2_23[37]}
   );
   gpc1163_5 gpc3123 (
      {stage1_24[23], stage1_24[24], stage1_24[25]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage1_26[0]},
      {stage1_27[0]},
      {stage2_28[0],stage2_27[5],stage2_26[8],stage2_25[21],stage2_24[33]}
   );
   gpc1163_5 gpc3124 (
      {stage1_24[26], stage1_24[27], stage1_24[28]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage1_26[1]},
      {stage1_27[1]},
      {stage2_28[1],stage2_27[6],stage2_26[9],stage2_25[22],stage2_24[34]}
   );
   gpc1163_5 gpc3125 (
      {stage1_24[29], stage1_24[30], stage1_24[31]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage1_26[2]},
      {stage1_27[2]},
      {stage2_28[2],stage2_27[7],stage2_26[10],stage2_25[23],stage2_24[35]}
   );
   gpc1163_5 gpc3126 (
      {stage1_24[32], stage1_24[33], stage1_24[34]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage1_26[3]},
      {stage1_27[3]},
      {stage2_28[3],stage2_27[8],stage2_26[11],stage2_25[24],stage2_24[36]}
   );
   gpc615_5 gpc3127 (
      {stage1_24[35], stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39]},
      {stage1_25[54]},
      {stage1_26[4], stage1_26[5], stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9]},
      {stage2_28[4],stage2_27[9],stage2_26[12],stage2_25[25],stage2_24[37]}
   );
   gpc615_5 gpc3128 (
      {stage1_24[40], stage1_24[41], stage1_24[42], stage1_24[43], stage1_24[44]},
      {stage1_25[55]},
      {stage1_26[10], stage1_26[11], stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15]},
      {stage2_28[5],stage2_27[10],stage2_26[13],stage2_25[26],stage2_24[38]}
   );
   gpc615_5 gpc3129 (
      {stage1_24[45], stage1_24[46], stage1_24[47], stage1_24[48], stage1_24[49]},
      {stage1_25[56]},
      {stage1_26[16], stage1_26[17], stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21]},
      {stage2_28[6],stage2_27[11],stage2_26[14],stage2_25[27],stage2_24[39]}
   );
   gpc615_5 gpc3130 (
      {stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53], stage1_24[54]},
      {stage1_25[57]},
      {stage1_26[22], stage1_26[23], stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27]},
      {stage2_28[7],stage2_27[12],stage2_26[15],stage2_25[28],stage2_24[40]}
   );
   gpc615_5 gpc3131 (
      {stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage1_25[58]},
      {stage1_26[28], stage1_26[29], stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33]},
      {stage2_28[8],stage2_27[13],stage2_26[16],stage2_25[29],stage2_24[41]}
   );
   gpc615_5 gpc3132 (
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64]},
      {stage1_25[59]},
      {stage1_26[34], stage1_26[35], stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39]},
      {stage2_28[9],stage2_27[14],stage2_26[17],stage2_25[30],stage2_24[42]}
   );
   gpc615_5 gpc3133 (
      {stage1_24[65], stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69]},
      {stage1_25[60]},
      {stage1_26[40], stage1_26[41], stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45]},
      {stage2_28[10],stage2_27[15],stage2_26[18],stage2_25[31],stage2_24[43]}
   );
   gpc615_5 gpc3134 (
      {stage1_24[70], stage1_24[71], stage1_24[72], stage1_24[73], stage1_24[74]},
      {stage1_25[61]},
      {stage1_26[46], stage1_26[47], stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51]},
      {stage2_28[11],stage2_27[16],stage2_26[19],stage2_25[32],stage2_24[44]}
   );
   gpc615_5 gpc3135 (
      {stage1_24[75], stage1_24[76], stage1_24[77], stage1_24[78], stage1_24[79]},
      {stage1_25[62]},
      {stage1_26[52], stage1_26[53], stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57]},
      {stage2_28[12],stage2_27[17],stage2_26[20],stage2_25[33],stage2_24[45]}
   );
   gpc615_5 gpc3136 (
      {stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83], stage1_24[84]},
      {stage1_25[63]},
      {stage1_26[58], stage1_26[59], stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63]},
      {stage2_28[13],stage2_27[18],stage2_26[21],stage2_25[34],stage2_24[46]}
   );
   gpc615_5 gpc3137 (
      {stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage1_25[64]},
      {stage1_26[64], stage1_26[65], stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69]},
      {stage2_28[14],stage2_27[19],stage2_26[22],stage2_25[35],stage2_24[47]}
   );
   gpc615_5 gpc3138 (
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94]},
      {stage1_25[65]},
      {stage1_26[70], stage1_26[71], stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75]},
      {stage2_28[15],stage2_27[20],stage2_26[23],stage2_25[36],stage2_24[48]}
   );
   gpc615_5 gpc3139 (
      {stage1_24[95], stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99]},
      {stage1_25[66]},
      {stage1_26[76], stage1_26[77], stage1_26[78], stage1_26[79], stage1_26[80], stage1_26[81]},
      {stage2_28[16],stage2_27[21],stage2_26[24],stage2_25[37],stage2_24[49]}
   );
   gpc615_5 gpc3140 (
      {stage1_24[100], stage1_24[101], stage1_24[102], stage1_24[103], stage1_24[104]},
      {stage1_25[67]},
      {stage1_26[82], stage1_26[83], stage1_26[84], stage1_26[85], stage1_26[86], stage1_26[87]},
      {stage2_28[17],stage2_27[22],stage2_26[25],stage2_25[38],stage2_24[50]}
   );
   gpc615_5 gpc3141 (
      {stage1_24[105], stage1_24[106], stage1_24[107], stage1_24[108], stage1_24[109]},
      {stage1_25[68]},
      {stage1_26[88], stage1_26[89], stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93]},
      {stage2_28[18],stage2_27[23],stage2_26[26],stage2_25[39],stage2_24[51]}
   );
   gpc606_5 gpc3142 (
      {stage1_25[69], stage1_25[70], stage1_25[71], stage1_25[72], stage1_25[73], stage1_25[74]},
      {stage1_27[4], stage1_27[5], stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9]},
      {stage2_29[0],stage2_28[19],stage2_27[24],stage2_26[27],stage2_25[40]}
   );
   gpc606_5 gpc3143 (
      {stage1_25[75], stage1_25[76], stage1_25[77], stage1_25[78], stage1_25[79], stage1_25[80]},
      {stage1_27[10], stage1_27[11], stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15]},
      {stage2_29[1],stage2_28[20],stage2_27[25],stage2_26[28],stage2_25[41]}
   );
   gpc606_5 gpc3144 (
      {stage1_25[81], stage1_25[82], stage1_25[83], stage1_25[84], stage1_25[85], stage1_25[86]},
      {stage1_27[16], stage1_27[17], stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21]},
      {stage2_29[2],stage2_28[21],stage2_27[26],stage2_26[29],stage2_25[42]}
   );
   gpc606_5 gpc3145 (
      {stage1_25[87], stage1_25[88], stage1_25[89], stage1_25[90], stage1_25[91], stage1_25[92]},
      {stage1_27[22], stage1_27[23], stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27]},
      {stage2_29[3],stage2_28[22],stage2_27[27],stage2_26[30],stage2_25[43]}
   );
   gpc606_5 gpc3146 (
      {stage1_25[93], stage1_25[94], stage1_25[95], stage1_25[96], stage1_25[97], stage1_25[98]},
      {stage1_27[28], stage1_27[29], stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33]},
      {stage2_29[4],stage2_28[23],stage2_27[28],stage2_26[31],stage2_25[44]}
   );
   gpc606_5 gpc3147 (
      {stage1_25[99], stage1_25[100], stage1_25[101], stage1_25[102], stage1_25[103], stage1_25[104]},
      {stage1_27[34], stage1_27[35], stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39]},
      {stage2_29[5],stage2_28[24],stage2_27[29],stage2_26[32],stage2_25[45]}
   );
   gpc615_5 gpc3148 (
      {stage1_26[94], stage1_26[95], stage1_26[96], stage1_26[97], stage1_26[98]},
      {stage1_27[40]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[6],stage2_28[25],stage2_27[30],stage2_26[33]}
   );
   gpc615_5 gpc3149 (
      {stage1_26[99], stage1_26[100], stage1_26[101], stage1_26[102], stage1_26[103]},
      {stage1_27[41]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[7],stage2_28[26],stage2_27[31],stage2_26[34]}
   );
   gpc615_5 gpc3150 (
      {stage1_26[104], stage1_26[105], stage1_26[106], stage1_26[107], stage1_26[108]},
      {stage1_27[42]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[8],stage2_28[27],stage2_27[32],stage2_26[35]}
   );
   gpc615_5 gpc3151 (
      {stage1_26[109], stage1_26[110], stage1_26[111], stage1_26[112], stage1_26[113]},
      {stage1_27[43]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[9],stage2_28[28],stage2_27[33],stage2_26[36]}
   );
   gpc615_5 gpc3152 (
      {stage1_26[114], stage1_26[115], stage1_26[116], stage1_26[117], stage1_26[118]},
      {stage1_27[44]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[10],stage2_28[29],stage2_27[34],stage2_26[37]}
   );
   gpc615_5 gpc3153 (
      {stage1_26[119], stage1_26[120], stage1_26[121], stage1_26[122], stage1_26[123]},
      {stage1_27[45]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[11],stage2_28[30],stage2_27[35],stage2_26[38]}
   );
   gpc615_5 gpc3154 (
      {stage1_26[124], stage1_26[125], stage1_26[126], stage1_26[127], stage1_26[128]},
      {stage1_27[46]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[12],stage2_28[31],stage2_27[36],stage2_26[39]}
   );
   gpc606_5 gpc3155 (
      {stage1_27[47], stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[7],stage2_29[13],stage2_28[32],stage2_27[37]}
   );
   gpc615_5 gpc3156 (
      {stage1_27[53], stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57]},
      {stage1_28[42]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[8],stage2_29[14],stage2_28[33],stage2_27[38]}
   );
   gpc615_5 gpc3157 (
      {stage1_27[58], stage1_27[59], stage1_27[60], stage1_27[61], stage1_27[62]},
      {stage1_28[43]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[9],stage2_29[15],stage2_28[34],stage2_27[39]}
   );
   gpc615_5 gpc3158 (
      {stage1_27[63], stage1_27[64], stage1_27[65], stage1_27[66], stage1_27[67]},
      {stage1_28[44]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[10],stage2_29[16],stage2_28[35],stage2_27[40]}
   );
   gpc615_5 gpc3159 (
      {stage1_27[68], stage1_27[69], stage1_27[70], stage1_27[71], stage1_27[72]},
      {stage1_28[45]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[11],stage2_29[17],stage2_28[36],stage2_27[41]}
   );
   gpc615_5 gpc3160 (
      {stage1_27[73], stage1_27[74], stage1_27[75], stage1_27[76], stage1_27[77]},
      {stage1_28[46]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[12],stage2_29[18],stage2_28[37],stage2_27[42]}
   );
   gpc615_5 gpc3161 (
      {stage1_27[78], stage1_27[79], stage1_27[80], stage1_27[81], stage1_27[82]},
      {stage1_28[47]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[13],stage2_29[19],stage2_28[38],stage2_27[43]}
   );
   gpc615_5 gpc3162 (
      {stage1_27[83], stage1_27[84], stage1_27[85], stage1_27[86], stage1_27[87]},
      {stage1_28[48]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[14],stage2_29[20],stage2_28[39],stage2_27[44]}
   );
   gpc615_5 gpc3163 (
      {stage1_27[88], stage1_27[89], stage1_27[90], stage1_27[91], stage1_27[92]},
      {stage1_28[49]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[15],stage2_29[21],stage2_28[40],stage2_27[45]}
   );
   gpc606_5 gpc3164 (
      {stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53], stage1_28[54], stage1_28[55]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[9],stage2_30[16],stage2_29[22],stage2_28[41]}
   );
   gpc606_5 gpc3165 (
      {stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59], stage1_28[60], stage1_28[61]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[10],stage2_30[17],stage2_29[23],stage2_28[42]}
   );
   gpc606_5 gpc3166 (
      {stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65], stage1_28[66], stage1_28[67]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[11],stage2_30[18],stage2_29[24],stage2_28[43]}
   );
   gpc606_5 gpc3167 (
      {stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71], stage1_28[72], stage1_28[73]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[12],stage2_30[19],stage2_29[25],stage2_28[44]}
   );
   gpc606_5 gpc3168 (
      {stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77], stage1_28[78], stage1_28[79]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[13],stage2_30[20],stage2_29[26],stage2_28[45]}
   );
   gpc606_5 gpc3169 (
      {stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83], stage1_28[84], stage1_28[85]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[14],stage2_30[21],stage2_29[27],stage2_28[46]}
   );
   gpc606_5 gpc3170 (
      {stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89], stage1_28[90], stage1_28[91]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[15],stage2_30[22],stage2_29[28],stage2_28[47]}
   );
   gpc606_5 gpc3171 (
      {stage1_28[92], stage1_28[93], stage1_28[94], stage1_28[95], stage1_28[96], stage1_28[97]},
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage2_32[7],stage2_31[16],stage2_30[23],stage2_29[29],stage2_28[48]}
   );
   gpc606_5 gpc3172 (
      {stage1_28[98], stage1_28[99], stage1_28[100], stage1_28[101], stage1_28[102], stage1_28[103]},
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage2_32[8],stage2_31[17],stage2_30[24],stage2_29[30],stage2_28[49]}
   );
   gpc1415_5 gpc3173 (
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58]},
      {stage1_30[54]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3]},
      {stage1_32[0]},
      {stage2_33[0],stage2_32[9],stage2_31[18],stage2_30[25],stage2_29[31]}
   );
   gpc606_5 gpc3174 (
      {stage1_29[59], stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64]},
      {stage1_31[4], stage1_31[5], stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9]},
      {stage2_33[1],stage2_32[10],stage2_31[19],stage2_30[26],stage2_29[32]}
   );
   gpc606_5 gpc3175 (
      {stage1_29[65], stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70]},
      {stage1_31[10], stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15]},
      {stage2_33[2],stage2_32[11],stage2_31[20],stage2_30[27],stage2_29[33]}
   );
   gpc606_5 gpc3176 (
      {stage1_29[71], stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76]},
      {stage1_31[16], stage1_31[17], stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21]},
      {stage2_33[3],stage2_32[12],stage2_31[21],stage2_30[28],stage2_29[34]}
   );
   gpc606_5 gpc3177 (
      {stage1_29[77], stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82]},
      {stage1_31[22], stage1_31[23], stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27]},
      {stage2_33[4],stage2_32[13],stage2_31[22],stage2_30[29],stage2_29[35]}
   );
   gpc606_5 gpc3178 (
      {stage1_29[83], stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88]},
      {stage1_31[28], stage1_31[29], stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33]},
      {stage2_33[5],stage2_32[14],stage2_31[23],stage2_30[30],stage2_29[36]}
   );
   gpc615_5 gpc3179 (
      {stage1_29[89], stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93]},
      {stage1_30[55]},
      {stage1_31[34], stage1_31[35], stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39]},
      {stage2_33[6],stage2_32[15],stage2_31[24],stage2_30[31],stage2_29[37]}
   );
   gpc615_5 gpc3180 (
      {stage1_29[94], stage1_29[95], stage1_29[96], stage1_29[97], stage1_29[98]},
      {stage1_30[56]},
      {stage1_31[40], stage1_31[41], stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45]},
      {stage2_33[7],stage2_32[16],stage2_31[25],stage2_30[32],stage2_29[38]}
   );
   gpc615_5 gpc3181 (
      {stage1_29[99], stage1_29[100], stage1_29[101], stage1_29[102], stage1_29[103]},
      {stage1_30[57]},
      {stage1_31[46], stage1_31[47], stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51]},
      {stage2_33[8],stage2_32[17],stage2_31[26],stage2_30[33],stage2_29[39]}
   );
   gpc615_5 gpc3182 (
      {stage1_30[58], stage1_30[59], stage1_30[60], stage1_30[61], stage1_30[62]},
      {stage1_31[52]},
      {stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5], stage1_32[6]},
      {stage2_34[0],stage2_33[9],stage2_32[18],stage2_31[27],stage2_30[34]}
   );
   gpc615_5 gpc3183 (
      {stage1_30[63], stage1_30[64], stage1_30[65], stage1_30[66], stage1_30[67]},
      {stage1_31[53]},
      {stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11], stage1_32[12]},
      {stage2_34[1],stage2_33[10],stage2_32[19],stage2_31[28],stage2_30[35]}
   );
   gpc615_5 gpc3184 (
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58]},
      {stage1_32[13]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[2],stage2_33[11],stage2_32[20],stage2_31[29]}
   );
   gpc615_5 gpc3185 (
      {stage1_31[59], stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63]},
      {stage1_32[14]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[3],stage2_33[12],stage2_32[21],stage2_31[30]}
   );
   gpc615_5 gpc3186 (
      {stage1_31[64], stage1_31[65], stage1_31[66], stage1_31[67], stage1_31[68]},
      {stage1_32[15]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[4],stage2_33[13],stage2_32[22],stage2_31[31]}
   );
   gpc615_5 gpc3187 (
      {stage1_31[69], stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73]},
      {stage1_32[16]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[5],stage2_33[14],stage2_32[23],stage2_31[32]}
   );
   gpc615_5 gpc3188 (
      {stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78]},
      {stage1_32[17]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[6],stage2_33[15],stage2_32[24],stage2_31[33]}
   );
   gpc615_5 gpc3189 (
      {stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage1_32[18]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage2_35[5],stage2_34[7],stage2_33[16],stage2_32[25],stage2_31[34]}
   );
   gpc615_5 gpc3190 (
      {stage1_31[84], stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88]},
      {stage1_32[19]},
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41]},
      {stage2_35[6],stage2_34[8],stage2_33[17],stage2_32[26],stage2_31[35]}
   );
   gpc615_5 gpc3191 (
      {stage1_31[89], stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93]},
      {stage1_32[20]},
      {stage1_33[42], stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47]},
      {stage2_35[7],stage2_34[9],stage2_33[18],stage2_32[27],stage2_31[36]}
   );
   gpc615_5 gpc3192 (
      {stage1_31[94], stage1_31[95], stage1_31[96], stage1_31[97], stage1_31[98]},
      {stage1_32[21]},
      {stage1_33[48], stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53]},
      {stage2_35[8],stage2_34[10],stage2_33[19],stage2_32[28],stage2_31[37]}
   );
   gpc606_5 gpc3193 (
      {stage1_32[22], stage1_32[23], stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[9],stage2_34[11],stage2_33[20],stage2_32[29]}
   );
   gpc606_5 gpc3194 (
      {stage1_32[28], stage1_32[29], stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33]},
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11]},
      {stage2_36[1],stage2_35[10],stage2_34[12],stage2_33[21],stage2_32[30]}
   );
   gpc606_5 gpc3195 (
      {stage1_32[34], stage1_32[35], stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39]},
      {stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17]},
      {stage2_36[2],stage2_35[11],stage2_34[13],stage2_33[22],stage2_32[31]}
   );
   gpc606_5 gpc3196 (
      {stage1_32[40], stage1_32[41], stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45]},
      {stage1_34[18], stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23]},
      {stage2_36[3],stage2_35[12],stage2_34[14],stage2_33[23],stage2_32[32]}
   );
   gpc606_5 gpc3197 (
      {stage1_32[46], stage1_32[47], stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51]},
      {stage1_34[24], stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29]},
      {stage2_36[4],stage2_35[13],stage2_34[15],stage2_33[24],stage2_32[33]}
   );
   gpc606_5 gpc3198 (
      {stage1_32[52], stage1_32[53], stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57]},
      {stage1_34[30], stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35]},
      {stage2_36[5],stage2_35[14],stage2_34[16],stage2_33[25],stage2_32[34]}
   );
   gpc606_5 gpc3199 (
      {stage1_32[58], stage1_32[59], stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63]},
      {stage1_34[36], stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40], stage1_34[41]},
      {stage2_36[6],stage2_35[15],stage2_34[17],stage2_33[26],stage2_32[35]}
   );
   gpc606_5 gpc3200 (
      {stage1_32[64], stage1_32[65], stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69]},
      {stage1_34[42], stage1_34[43], stage1_34[44], stage1_34[45], stage1_34[46], stage1_34[47]},
      {stage2_36[7],stage2_35[16],stage2_34[18],stage2_33[27],stage2_32[36]}
   );
   gpc606_5 gpc3201 (
      {stage1_32[70], stage1_32[71], stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75]},
      {stage1_34[48], stage1_34[49], stage1_34[50], stage1_34[51], stage1_34[52], stage1_34[53]},
      {stage2_36[8],stage2_35[17],stage2_34[19],stage2_33[28],stage2_32[37]}
   );
   gpc606_5 gpc3202 (
      {stage1_32[76], stage1_32[77], stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81]},
      {stage1_34[54], stage1_34[55], stage1_34[56], stage1_34[57], stage1_34[58], stage1_34[59]},
      {stage2_36[9],stage2_35[18],stage2_34[20],stage2_33[29],stage2_32[38]}
   );
   gpc606_5 gpc3203 (
      {stage1_32[82], stage1_32[83], stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87]},
      {stage1_34[60], stage1_34[61], stage1_34[62], stage1_34[63], stage1_34[64], stage1_34[65]},
      {stage2_36[10],stage2_35[19],stage2_34[21],stage2_33[30],stage2_32[39]}
   );
   gpc606_5 gpc3204 (
      {stage1_32[88], stage1_32[89], stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93]},
      {stage1_34[66], stage1_34[67], stage1_34[68], stage1_34[69], stage1_34[70], stage1_34[71]},
      {stage2_36[11],stage2_35[20],stage2_34[22],stage2_33[31],stage2_32[40]}
   );
   gpc606_5 gpc3205 (
      {stage1_32[94], stage1_32[95], stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99]},
      {stage1_34[72], stage1_34[73], stage1_34[74], stage1_34[75], stage1_34[76], stage1_34[77]},
      {stage2_36[12],stage2_35[21],stage2_34[23],stage2_33[32],stage2_32[41]}
   );
   gpc606_5 gpc3206 (
      {stage1_32[100], stage1_32[101], stage1_32[102], stage1_32[103], stage1_32[104], stage1_32[105]},
      {stage1_34[78], stage1_34[79], stage1_34[80], stage1_34[81], stage1_34[82], stage1_34[83]},
      {stage2_36[13],stage2_35[22],stage2_34[24],stage2_33[33],stage2_32[42]}
   );
   gpc606_5 gpc3207 (
      {stage1_32[106], stage1_32[107], stage1_32[108], stage1_32[109], stage1_32[110], stage1_32[111]},
      {stage1_34[84], stage1_34[85], stage1_34[86], stage1_34[87], stage1_34[88], stage1_34[89]},
      {stage2_36[14],stage2_35[23],stage2_34[25],stage2_33[34],stage2_32[43]}
   );
   gpc606_5 gpc3208 (
      {stage1_33[54], stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[15],stage2_35[24],stage2_34[26],stage2_33[35]}
   );
   gpc606_5 gpc3209 (
      {stage1_33[60], stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[16],stage2_35[25],stage2_34[27],stage2_33[36]}
   );
   gpc606_5 gpc3210 (
      {stage1_33[66], stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[17],stage2_35[26],stage2_34[28],stage2_33[37]}
   );
   gpc606_5 gpc3211 (
      {stage1_33[72], stage1_33[73], stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77]},
      {stage1_35[18], stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23]},
      {stage2_37[3],stage2_36[18],stage2_35[27],stage2_34[29],stage2_33[38]}
   );
   gpc606_5 gpc3212 (
      {stage1_33[78], stage1_33[79], stage1_33[80], stage1_33[81], stage1_33[82], stage1_33[83]},
      {stage1_35[24], stage1_35[25], stage1_35[26], stage1_35[27], stage1_35[28], stage1_35[29]},
      {stage2_37[4],stage2_36[19],stage2_35[28],stage2_34[30],stage2_33[39]}
   );
   gpc606_5 gpc3213 (
      {stage1_33[84], stage1_33[85], stage1_33[86], stage1_33[87], stage1_33[88], stage1_33[89]},
      {stage1_35[30], stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35]},
      {stage2_37[5],stage2_36[20],stage2_35[29],stage2_34[31],stage2_33[40]}
   );
   gpc606_5 gpc3214 (
      {stage1_33[90], stage1_33[91], stage1_33[92], stage1_33[93], stage1_33[94], stage1_33[95]},
      {stage1_35[36], stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40], stage1_35[41]},
      {stage2_37[6],stage2_36[21],stage2_35[30],stage2_34[32],stage2_33[41]}
   );
   gpc606_5 gpc3215 (
      {stage1_33[96], stage1_33[97], stage1_33[98], stage1_33[99], stage1_33[100], stage1_33[101]},
      {stage1_35[42], stage1_35[43], stage1_35[44], stage1_35[45], stage1_35[46], stage1_35[47]},
      {stage2_37[7],stage2_36[22],stage2_35[31],stage2_34[33],stage2_33[42]}
   );
   gpc615_5 gpc3216 (
      {stage1_34[90], stage1_34[91], stage1_34[92], stage1_34[93], stage1_34[94]},
      {stage1_35[48]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[8],stage2_36[23],stage2_35[32],stage2_34[34]}
   );
   gpc615_5 gpc3217 (
      {stage1_34[95], stage1_34[96], stage1_34[97], stage1_34[98], stage1_34[99]},
      {stage1_35[49]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[9],stage2_36[24],stage2_35[33],stage2_34[35]}
   );
   gpc615_5 gpc3218 (
      {stage1_34[100], stage1_34[101], stage1_34[102], stage1_34[103], 1'b0},
      {stage1_35[50]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[10],stage2_36[25],stage2_35[34],stage2_34[36]}
   );
   gpc615_5 gpc3219 (
      {stage1_35[51], stage1_35[52], stage1_35[53], stage1_35[54], stage1_35[55]},
      {stage1_36[18]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[3],stage2_37[11],stage2_36[26],stage2_35[35]}
   );
   gpc615_5 gpc3220 (
      {stage1_35[56], stage1_35[57], stage1_35[58], stage1_35[59], stage1_35[60]},
      {stage1_36[19]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[4],stage2_37[12],stage2_36[27],stage2_35[36]}
   );
   gpc615_5 gpc3221 (
      {stage1_35[61], stage1_35[62], stage1_35[63], stage1_35[64], stage1_35[65]},
      {stage1_36[20]},
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage2_39[2],stage2_38[5],stage2_37[13],stage2_36[28],stage2_35[37]}
   );
   gpc615_5 gpc3222 (
      {stage1_35[66], stage1_35[67], stage1_35[68], stage1_35[69], stage1_35[70]},
      {stage1_36[21]},
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage2_39[3],stage2_38[6],stage2_37[14],stage2_36[29],stage2_35[38]}
   );
   gpc615_5 gpc3223 (
      {stage1_35[71], stage1_35[72], stage1_35[73], stage1_35[74], stage1_35[75]},
      {stage1_36[22]},
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28], stage1_37[29]},
      {stage2_39[4],stage2_38[7],stage2_37[15],stage2_36[30],stage2_35[39]}
   );
   gpc615_5 gpc3224 (
      {stage1_35[76], stage1_35[77], stage1_35[78], stage1_35[79], stage1_35[80]},
      {stage1_36[23]},
      {stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33], stage1_37[34], stage1_37[35]},
      {stage2_39[5],stage2_38[8],stage2_37[16],stage2_36[31],stage2_35[40]}
   );
   gpc615_5 gpc3225 (
      {stage1_35[81], stage1_35[82], stage1_35[83], stage1_35[84], stage1_35[85]},
      {stage1_36[24]},
      {stage1_37[36], stage1_37[37], stage1_37[38], stage1_37[39], stage1_37[40], stage1_37[41]},
      {stage2_39[6],stage2_38[9],stage2_37[17],stage2_36[32],stage2_35[41]}
   );
   gpc615_5 gpc3226 (
      {stage1_35[86], stage1_35[87], stage1_35[88], stage1_35[89], stage1_35[90]},
      {stage1_36[25]},
      {stage1_37[42], stage1_37[43], stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47]},
      {stage2_39[7],stage2_38[10],stage2_37[18],stage2_36[33],stage2_35[42]}
   );
   gpc615_5 gpc3227 (
      {stage1_35[91], stage1_35[92], stage1_35[93], stage1_35[94], stage1_35[95]},
      {stage1_36[26]},
      {stage1_37[48], stage1_37[49], stage1_37[50], stage1_37[51], stage1_37[52], stage1_37[53]},
      {stage2_39[8],stage2_38[11],stage2_37[19],stage2_36[34],stage2_35[43]}
   );
   gpc615_5 gpc3228 (
      {stage1_35[96], stage1_35[97], stage1_35[98], stage1_35[99], stage1_35[100]},
      {stage1_36[27]},
      {stage1_37[54], stage1_37[55], stage1_37[56], stage1_37[57], stage1_37[58], stage1_37[59]},
      {stage2_39[9],stage2_38[12],stage2_37[20],stage2_36[35],stage2_35[44]}
   );
   gpc615_5 gpc3229 (
      {stage1_35[101], stage1_35[102], stage1_35[103], stage1_35[104], stage1_35[105]},
      {stage1_36[28]},
      {stage1_37[60], stage1_37[61], stage1_37[62], stage1_37[63], stage1_37[64], stage1_37[65]},
      {stage2_39[10],stage2_38[13],stage2_37[21],stage2_36[36],stage2_35[45]}
   );
   gpc135_4 gpc3230 (
      {stage1_36[29], stage1_36[30], stage1_36[31], stage1_36[32], stage1_36[33]},
      {stage1_37[66], stage1_37[67], stage1_37[68]},
      {stage1_38[0]},
      {stage2_39[11],stage2_38[14],stage2_37[22],stage2_36[37]}
   );
   gpc135_4 gpc3231 (
      {stage1_36[34], stage1_36[35], stage1_36[36], stage1_36[37], stage1_36[38]},
      {stage1_37[69], stage1_37[70], stage1_37[71]},
      {stage1_38[1]},
      {stage2_39[12],stage2_38[15],stage2_37[23],stage2_36[38]}
   );
   gpc135_4 gpc3232 (
      {stage1_36[39], stage1_36[40], stage1_36[41], stage1_36[42], stage1_36[43]},
      {stage1_37[72], stage1_37[73], stage1_37[74]},
      {stage1_38[2]},
      {stage2_39[13],stage2_38[16],stage2_37[24],stage2_36[39]}
   );
   gpc135_4 gpc3233 (
      {stage1_36[44], stage1_36[45], stage1_36[46], stage1_36[47], stage1_36[48]},
      {stage1_37[75], stage1_37[76], stage1_37[77]},
      {stage1_38[3]},
      {stage2_39[14],stage2_38[17],stage2_37[25],stage2_36[40]}
   );
   gpc135_4 gpc3234 (
      {stage1_36[49], stage1_36[50], stage1_36[51], stage1_36[52], stage1_36[53]},
      {stage1_37[78], stage1_37[79], stage1_37[80]},
      {stage1_38[4]},
      {stage2_39[15],stage2_38[18],stage2_37[26],stage2_36[41]}
   );
   gpc606_5 gpc3235 (
      {stage1_36[54], stage1_36[55], stage1_36[56], stage1_36[57], stage1_36[58], stage1_36[59]},
      {stage1_38[5], stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10]},
      {stage2_40[0],stage2_39[16],stage2_38[19],stage2_37[27],stage2_36[42]}
   );
   gpc606_5 gpc3236 (
      {stage1_36[60], stage1_36[61], stage1_36[62], stage1_36[63], stage1_36[64], stage1_36[65]},
      {stage1_38[11], stage1_38[12], stage1_38[13], stage1_38[14], stage1_38[15], stage1_38[16]},
      {stage2_40[1],stage2_39[17],stage2_38[20],stage2_37[28],stage2_36[43]}
   );
   gpc606_5 gpc3237 (
      {stage1_36[66], stage1_36[67], stage1_36[68], stage1_36[69], stage1_36[70], stage1_36[71]},
      {stage1_38[17], stage1_38[18], stage1_38[19], stage1_38[20], stage1_38[21], stage1_38[22]},
      {stage2_40[2],stage2_39[18],stage2_38[21],stage2_37[29],stage2_36[44]}
   );
   gpc606_5 gpc3238 (
      {stage1_36[72], stage1_36[73], stage1_36[74], stage1_36[75], stage1_36[76], stage1_36[77]},
      {stage1_38[23], stage1_38[24], stage1_38[25], stage1_38[26], stage1_38[27], stage1_38[28]},
      {stage2_40[3],stage2_39[19],stage2_38[22],stage2_37[30],stage2_36[45]}
   );
   gpc606_5 gpc3239 (
      {stage1_36[78], stage1_36[79], stage1_36[80], stage1_36[81], stage1_36[82], stage1_36[83]},
      {stage1_38[29], stage1_38[30], stage1_38[31], stage1_38[32], stage1_38[33], stage1_38[34]},
      {stage2_40[4],stage2_39[20],stage2_38[23],stage2_37[31],stage2_36[46]}
   );
   gpc606_5 gpc3240 (
      {stage1_36[84], stage1_36[85], stage1_36[86], stage1_36[87], stage1_36[88], stage1_36[89]},
      {stage1_38[35], stage1_38[36], stage1_38[37], stage1_38[38], stage1_38[39], stage1_38[40]},
      {stage2_40[5],stage2_39[21],stage2_38[24],stage2_37[32],stage2_36[47]}
   );
   gpc606_5 gpc3241 (
      {stage1_36[90], stage1_36[91], stage1_36[92], stage1_36[93], stage1_36[94], stage1_36[95]},
      {stage1_38[41], stage1_38[42], stage1_38[43], stage1_38[44], stage1_38[45], stage1_38[46]},
      {stage2_40[6],stage2_39[22],stage2_38[25],stage2_37[33],stage2_36[48]}
   );
   gpc606_5 gpc3242 (
      {stage1_36[96], stage1_36[97], stage1_36[98], stage1_36[99], stage1_36[100], stage1_36[101]},
      {stage1_38[47], stage1_38[48], stage1_38[49], stage1_38[50], stage1_38[51], stage1_38[52]},
      {stage2_40[7],stage2_39[23],stage2_38[26],stage2_37[34],stage2_36[49]}
   );
   gpc606_5 gpc3243 (
      {stage1_36[102], stage1_36[103], stage1_36[104], stage1_36[105], stage1_36[106], stage1_36[107]},
      {stage1_38[53], stage1_38[54], stage1_38[55], stage1_38[56], stage1_38[57], stage1_38[58]},
      {stage2_40[8],stage2_39[24],stage2_38[27],stage2_37[35],stage2_36[50]}
   );
   gpc606_5 gpc3244 (
      {stage1_36[108], stage1_36[109], stage1_36[110], stage1_36[111], stage1_36[112], stage1_36[113]},
      {stage1_38[59], stage1_38[60], stage1_38[61], stage1_38[62], stage1_38[63], stage1_38[64]},
      {stage2_40[9],stage2_39[25],stage2_38[28],stage2_37[36],stage2_36[51]}
   );
   gpc606_5 gpc3245 (
      {stage1_36[114], stage1_36[115], stage1_36[116], stage1_36[117], stage1_36[118], stage1_36[119]},
      {stage1_38[65], stage1_38[66], stage1_38[67], stage1_38[68], stage1_38[69], stage1_38[70]},
      {stage2_40[10],stage2_39[26],stage2_38[29],stage2_37[37],stage2_36[52]}
   );
   gpc606_5 gpc3246 (
      {stage1_36[120], stage1_36[121], stage1_36[122], stage1_36[123], stage1_36[124], stage1_36[125]},
      {stage1_38[71], stage1_38[72], stage1_38[73], stage1_38[74], stage1_38[75], stage1_38[76]},
      {stage2_40[11],stage2_39[27],stage2_38[30],stage2_37[38],stage2_36[53]}
   );
   gpc606_5 gpc3247 (
      {stage1_36[126], stage1_36[127], stage1_36[128], stage1_36[129], stage1_36[130], stage1_36[131]},
      {stage1_38[77], stage1_38[78], stage1_38[79], stage1_38[80], stage1_38[81], stage1_38[82]},
      {stage2_40[12],stage2_39[28],stage2_38[31],stage2_37[39],stage2_36[54]}
   );
   gpc606_5 gpc3248 (
      {stage1_36[132], stage1_36[133], stage1_36[134], stage1_36[135], stage1_36[136], stage1_36[137]},
      {stage1_38[83], stage1_38[84], stage1_38[85], stage1_38[86], stage1_38[87], stage1_38[88]},
      {stage2_40[13],stage2_39[29],stage2_38[32],stage2_37[40],stage2_36[55]}
   );
   gpc606_5 gpc3249 (
      {stage1_37[81], stage1_37[82], stage1_37[83], stage1_37[84], stage1_37[85], stage1_37[86]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage2_41[0],stage2_40[14],stage2_39[30],stage2_38[33],stage2_37[41]}
   );
   gpc606_5 gpc3250 (
      {stage1_37[87], stage1_37[88], stage1_37[89], stage1_37[90], stage1_37[91], stage1_37[92]},
      {stage1_39[6], stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11]},
      {stage2_41[1],stage2_40[15],stage2_39[31],stage2_38[34],stage2_37[42]}
   );
   gpc615_5 gpc3251 (
      {stage1_38[89], stage1_38[90], stage1_38[91], stage1_38[92], stage1_38[93]},
      {stage1_39[12]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[2],stage2_40[16],stage2_39[32],stage2_38[35]}
   );
   gpc615_5 gpc3252 (
      {stage1_38[94], stage1_38[95], stage1_38[96], stage1_38[97], stage1_38[98]},
      {stage1_39[13]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[3],stage2_40[17],stage2_39[33],stage2_38[36]}
   );
   gpc615_5 gpc3253 (
      {stage1_38[99], stage1_38[100], stage1_38[101], stage1_38[102], stage1_38[103]},
      {stage1_39[14]},
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage2_42[2],stage2_41[4],stage2_40[18],stage2_39[34],stage2_38[37]}
   );
   gpc615_5 gpc3254 (
      {stage1_38[104], stage1_38[105], stage1_38[106], stage1_38[107], stage1_38[108]},
      {stage1_39[15]},
      {stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage2_42[3],stage2_41[5],stage2_40[19],stage2_39[35],stage2_38[38]}
   );
   gpc615_5 gpc3255 (
      {stage1_38[109], stage1_38[110], stage1_38[111], stage1_38[112], stage1_38[113]},
      {stage1_39[16]},
      {stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28], stage1_40[29]},
      {stage2_42[4],stage2_41[6],stage2_40[20],stage2_39[36],stage2_38[39]}
   );
   gpc615_5 gpc3256 (
      {stage1_38[114], stage1_38[115], stage1_38[116], stage1_38[117], stage1_38[118]},
      {stage1_39[17]},
      {stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34], stage1_40[35]},
      {stage2_42[5],stage2_41[7],stage2_40[21],stage2_39[37],stage2_38[40]}
   );
   gpc615_5 gpc3257 (
      {stage1_38[119], stage1_38[120], stage1_38[121], stage1_38[122], stage1_38[123]},
      {stage1_39[18]},
      {stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40], stage1_40[41]},
      {stage2_42[6],stage2_41[8],stage2_40[22],stage2_39[38],stage2_38[41]}
   );
   gpc615_5 gpc3258 (
      {stage1_38[124], stage1_38[125], stage1_38[126], stage1_38[127], stage1_38[128]},
      {stage1_39[19]},
      {stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46], stage1_40[47]},
      {stage2_42[7],stage2_41[9],stage2_40[23],stage2_39[39],stage2_38[42]}
   );
   gpc615_5 gpc3259 (
      {stage1_38[129], stage1_38[130], stage1_38[131], stage1_38[132], stage1_38[133]},
      {stage1_39[20]},
      {stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52], stage1_40[53]},
      {stage2_42[8],stage2_41[10],stage2_40[24],stage2_39[40],stage2_38[43]}
   );
   gpc606_5 gpc3260 (
      {stage1_39[21], stage1_39[22], stage1_39[23], stage1_39[24], stage1_39[25], stage1_39[26]},
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage2_43[0],stage2_42[9],stage2_41[11],stage2_40[25],stage2_39[41]}
   );
   gpc606_5 gpc3261 (
      {stage1_39[27], stage1_39[28], stage1_39[29], stage1_39[30], stage1_39[31], stage1_39[32]},
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11]},
      {stage2_43[1],stage2_42[10],stage2_41[12],stage2_40[26],stage2_39[42]}
   );
   gpc606_5 gpc3262 (
      {stage1_39[33], stage1_39[34], stage1_39[35], stage1_39[36], stage1_39[37], stage1_39[38]},
      {stage1_41[12], stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17]},
      {stage2_43[2],stage2_42[11],stage2_41[13],stage2_40[27],stage2_39[43]}
   );
   gpc606_5 gpc3263 (
      {stage1_39[39], stage1_39[40], stage1_39[41], stage1_39[42], stage1_39[43], stage1_39[44]},
      {stage1_41[18], stage1_41[19], stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23]},
      {stage2_43[3],stage2_42[12],stage2_41[14],stage2_40[28],stage2_39[44]}
   );
   gpc606_5 gpc3264 (
      {stage1_39[45], stage1_39[46], stage1_39[47], stage1_39[48], stage1_39[49], stage1_39[50]},
      {stage1_41[24], stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29]},
      {stage2_43[4],stage2_42[13],stage2_41[15],stage2_40[29],stage2_39[45]}
   );
   gpc606_5 gpc3265 (
      {stage1_39[51], stage1_39[52], stage1_39[53], stage1_39[54], stage1_39[55], stage1_39[56]},
      {stage1_41[30], stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34], stage1_41[35]},
      {stage2_43[5],stage2_42[14],stage2_41[16],stage2_40[30],stage2_39[46]}
   );
   gpc606_5 gpc3266 (
      {stage1_39[57], stage1_39[58], stage1_39[59], stage1_39[60], stage1_39[61], stage1_39[62]},
      {stage1_41[36], stage1_41[37], stage1_41[38], stage1_41[39], stage1_41[40], stage1_41[41]},
      {stage2_43[6],stage2_42[15],stage2_41[17],stage2_40[31],stage2_39[47]}
   );
   gpc606_5 gpc3267 (
      {stage1_39[63], stage1_39[64], stage1_39[65], stage1_39[66], stage1_39[67], stage1_39[68]},
      {stage1_41[42], stage1_41[43], stage1_41[44], stage1_41[45], stage1_41[46], stage1_41[47]},
      {stage2_43[7],stage2_42[16],stage2_41[18],stage2_40[32],stage2_39[48]}
   );
   gpc606_5 gpc3268 (
      {stage1_39[69], stage1_39[70], stage1_39[71], stage1_39[72], stage1_39[73], stage1_39[74]},
      {stage1_41[48], stage1_41[49], stage1_41[50], stage1_41[51], stage1_41[52], stage1_41[53]},
      {stage2_43[8],stage2_42[17],stage2_41[19],stage2_40[33],stage2_39[49]}
   );
   gpc606_5 gpc3269 (
      {stage1_39[75], stage1_39[76], stage1_39[77], stage1_39[78], stage1_39[79], stage1_39[80]},
      {stage1_41[54], stage1_41[55], stage1_41[56], stage1_41[57], stage1_41[58], stage1_41[59]},
      {stage2_43[9],stage2_42[18],stage2_41[20],stage2_40[34],stage2_39[50]}
   );
   gpc606_5 gpc3270 (
      {stage1_39[81], stage1_39[82], stage1_39[83], stage1_39[84], stage1_39[85], stage1_39[86]},
      {stage1_41[60], stage1_41[61], stage1_41[62], stage1_41[63], stage1_41[64], stage1_41[65]},
      {stage2_43[10],stage2_42[19],stage2_41[21],stage2_40[35],stage2_39[51]}
   );
   gpc606_5 gpc3271 (
      {stage1_39[87], stage1_39[88], stage1_39[89], stage1_39[90], stage1_39[91], stage1_39[92]},
      {stage1_41[66], stage1_41[67], stage1_41[68], stage1_41[69], stage1_41[70], stage1_41[71]},
      {stage2_43[11],stage2_42[20],stage2_41[22],stage2_40[36],stage2_39[52]}
   );
   gpc615_5 gpc3272 (
      {stage1_39[93], stage1_39[94], stage1_39[95], stage1_39[96], stage1_39[97]},
      {stage1_40[54]},
      {stage1_41[72], stage1_41[73], stage1_41[74], stage1_41[75], stage1_41[76], stage1_41[77]},
      {stage2_43[12],stage2_42[21],stage2_41[23],stage2_40[37],stage2_39[53]}
   );
   gpc606_5 gpc3273 (
      {stage1_40[55], stage1_40[56], stage1_40[57], stage1_40[58], stage1_40[59], stage1_40[60]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[13],stage2_42[22],stage2_41[24],stage2_40[38]}
   );
   gpc606_5 gpc3274 (
      {stage1_40[61], stage1_40[62], stage1_40[63], stage1_40[64], stage1_40[65], stage1_40[66]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[14],stage2_42[23],stage2_41[25],stage2_40[39]}
   );
   gpc606_5 gpc3275 (
      {stage1_40[67], stage1_40[68], stage1_40[69], stage1_40[70], stage1_40[71], stage1_40[72]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[15],stage2_42[24],stage2_41[26],stage2_40[40]}
   );
   gpc606_5 gpc3276 (
      {stage1_40[73], stage1_40[74], stage1_40[75], stage1_40[76], stage1_40[77], stage1_40[78]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[16],stage2_42[25],stage2_41[27],stage2_40[41]}
   );
   gpc606_5 gpc3277 (
      {stage1_40[79], stage1_40[80], stage1_40[81], stage1_40[82], stage1_40[83], stage1_40[84]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[17],stage2_42[26],stage2_41[28],stage2_40[42]}
   );
   gpc606_5 gpc3278 (
      {stage1_40[85], stage1_40[86], stage1_40[87], stage1_40[88], stage1_40[89], stage1_40[90]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[18],stage2_42[27],stage2_41[29],stage2_40[43]}
   );
   gpc606_5 gpc3279 (
      {stage1_41[78], stage1_41[79], stage1_41[80], stage1_41[81], stage1_41[82], stage1_41[83]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[6],stage2_43[19],stage2_42[28],stage2_41[30]}
   );
   gpc606_5 gpc3280 (
      {stage1_41[84], stage1_41[85], stage1_41[86], stage1_41[87], stage1_41[88], stage1_41[89]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[7],stage2_43[20],stage2_42[29],stage2_41[31]}
   );
   gpc606_5 gpc3281 (
      {stage1_41[90], stage1_41[91], stage1_41[92], stage1_41[93], stage1_41[94], stage1_41[95]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[8],stage2_43[21],stage2_42[30],stage2_41[32]}
   );
   gpc606_5 gpc3282 (
      {stage1_41[96], stage1_41[97], stage1_41[98], stage1_41[99], stage1_41[100], stage1_41[101]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[9],stage2_43[22],stage2_42[31],stage2_41[33]}
   );
   gpc606_5 gpc3283 (
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage2_46[0],stage2_45[4],stage2_44[10],stage2_43[23],stage2_42[32]}
   );
   gpc606_5 gpc3284 (
      {stage1_42[42], stage1_42[43], stage1_42[44], stage1_42[45], stage1_42[46], stage1_42[47]},
      {stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9], stage1_44[10], stage1_44[11]},
      {stage2_46[1],stage2_45[5],stage2_44[11],stage2_43[24],stage2_42[33]}
   );
   gpc606_5 gpc3285 (
      {stage1_42[48], stage1_42[49], stage1_42[50], stage1_42[51], stage1_42[52], stage1_42[53]},
      {stage1_44[12], stage1_44[13], stage1_44[14], stage1_44[15], stage1_44[16], stage1_44[17]},
      {stage2_46[2],stage2_45[6],stage2_44[12],stage2_43[25],stage2_42[34]}
   );
   gpc606_5 gpc3286 (
      {stage1_42[54], stage1_42[55], stage1_42[56], stage1_42[57], stage1_42[58], stage1_42[59]},
      {stage1_44[18], stage1_44[19], stage1_44[20], stage1_44[21], stage1_44[22], stage1_44[23]},
      {stage2_46[3],stage2_45[7],stage2_44[13],stage2_43[26],stage2_42[35]}
   );
   gpc606_5 gpc3287 (
      {stage1_42[60], stage1_42[61], stage1_42[62], stage1_42[63], stage1_42[64], stage1_42[65]},
      {stage1_44[24], stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28], stage1_44[29]},
      {stage2_46[4],stage2_45[8],stage2_44[14],stage2_43[27],stage2_42[36]}
   );
   gpc606_5 gpc3288 (
      {stage1_42[66], stage1_42[67], stage1_42[68], stage1_42[69], stage1_42[70], stage1_42[71]},
      {stage1_44[30], stage1_44[31], stage1_44[32], stage1_44[33], stage1_44[34], stage1_44[35]},
      {stage2_46[5],stage2_45[9],stage2_44[15],stage2_43[28],stage2_42[37]}
   );
   gpc606_5 gpc3289 (
      {stage1_42[72], stage1_42[73], stage1_42[74], stage1_42[75], stage1_42[76], stage1_42[77]},
      {stage1_44[36], stage1_44[37], stage1_44[38], stage1_44[39], stage1_44[40], stage1_44[41]},
      {stage2_46[6],stage2_45[10],stage2_44[16],stage2_43[29],stage2_42[38]}
   );
   gpc606_5 gpc3290 (
      {stage1_42[78], stage1_42[79], stage1_42[80], stage1_42[81], stage1_42[82], stage1_42[83]},
      {stage1_44[42], stage1_44[43], stage1_44[44], stage1_44[45], stage1_44[46], stage1_44[47]},
      {stage2_46[7],stage2_45[11],stage2_44[17],stage2_43[30],stage2_42[39]}
   );
   gpc606_5 gpc3291 (
      {stage1_42[84], stage1_42[85], stage1_42[86], stage1_42[87], stage1_42[88], stage1_42[89]},
      {stage1_44[48], stage1_44[49], stage1_44[50], stage1_44[51], stage1_44[52], stage1_44[53]},
      {stage2_46[8],stage2_45[12],stage2_44[18],stage2_43[31],stage2_42[40]}
   );
   gpc606_5 gpc3292 (
      {stage1_42[90], stage1_42[91], stage1_42[92], stage1_42[93], stage1_42[94], stage1_42[95]},
      {stage1_44[54], stage1_44[55], stage1_44[56], stage1_44[57], stage1_44[58], stage1_44[59]},
      {stage2_46[9],stage2_45[13],stage2_44[19],stage2_43[32],stage2_42[41]}
   );
   gpc606_5 gpc3293 (
      {stage1_42[96], stage1_42[97], stage1_42[98], stage1_42[99], stage1_42[100], stage1_42[101]},
      {stage1_44[60], stage1_44[61], stage1_44[62], stage1_44[63], stage1_44[64], stage1_44[65]},
      {stage2_46[10],stage2_45[14],stage2_44[20],stage2_43[33],stage2_42[42]}
   );
   gpc606_5 gpc3294 (
      {stage1_42[102], stage1_42[103], stage1_42[104], stage1_42[105], stage1_42[106], stage1_42[107]},
      {stage1_44[66], stage1_44[67], stage1_44[68], stage1_44[69], stage1_44[70], stage1_44[71]},
      {stage2_46[11],stage2_45[15],stage2_44[21],stage2_43[34],stage2_42[43]}
   );
   gpc606_5 gpc3295 (
      {stage1_42[108], stage1_42[109], stage1_42[110], stage1_42[111], stage1_42[112], stage1_42[113]},
      {stage1_44[72], stage1_44[73], stage1_44[74], stage1_44[75], stage1_44[76], stage1_44[77]},
      {stage2_46[12],stage2_45[16],stage2_44[22],stage2_43[35],stage2_42[44]}
   );
   gpc606_5 gpc3296 (
      {stage1_42[114], stage1_42[115], stage1_42[116], stage1_42[117], stage1_42[118], stage1_42[119]},
      {stage1_44[78], stage1_44[79], stage1_44[80], stage1_44[81], stage1_44[82], stage1_44[83]},
      {stage2_46[13],stage2_45[17],stage2_44[23],stage2_43[36],stage2_42[45]}
   );
   gpc606_5 gpc3297 (
      {stage1_42[120], stage1_42[121], stage1_42[122], stage1_42[123], stage1_42[124], stage1_42[125]},
      {stage1_44[84], stage1_44[85], stage1_44[86], stage1_44[87], stage1_44[88], stage1_44[89]},
      {stage2_46[14],stage2_45[18],stage2_44[24],stage2_43[37],stage2_42[46]}
   );
   gpc606_5 gpc3298 (
      {stage1_42[126], stage1_42[127], stage1_42[128], stage1_42[129], stage1_42[130], stage1_42[131]},
      {stage1_44[90], stage1_44[91], stage1_44[92], stage1_44[93], stage1_44[94], stage1_44[95]},
      {stage2_46[15],stage2_45[19],stage2_44[25],stage2_43[38],stage2_42[47]}
   );
   gpc606_5 gpc3299 (
      {stage1_42[132], stage1_42[133], stage1_42[134], stage1_42[135], stage1_42[136], stage1_42[137]},
      {stage1_44[96], stage1_44[97], stage1_44[98], stage1_44[99], stage1_44[100], stage1_44[101]},
      {stage2_46[16],stage2_45[20],stage2_44[26],stage2_43[39],stage2_42[48]}
   );
   gpc606_5 gpc3300 (
      {stage1_42[138], stage1_42[139], stage1_42[140], stage1_42[141], stage1_42[142], stage1_42[143]},
      {stage1_44[102], stage1_44[103], stage1_44[104], stage1_44[105], stage1_44[106], stage1_44[107]},
      {stage2_46[17],stage2_45[21],stage2_44[27],stage2_43[40],stage2_42[49]}
   );
   gpc606_5 gpc3301 (
      {stage1_42[144], stage1_42[145], stage1_42[146], stage1_42[147], stage1_42[148], stage1_42[149]},
      {stage1_44[108], stage1_44[109], stage1_44[110], stage1_44[111], stage1_44[112], stage1_44[113]},
      {stage2_46[18],stage2_45[22],stage2_44[28],stage2_43[41],stage2_42[50]}
   );
   gpc606_5 gpc3302 (
      {stage1_42[150], stage1_42[151], stage1_42[152], stage1_42[153], stage1_42[154], stage1_42[155]},
      {stage1_44[114], stage1_44[115], stage1_44[116], stage1_44[117], stage1_44[118], stage1_44[119]},
      {stage2_46[19],stage2_45[23],stage2_44[29],stage2_43[42],stage2_42[51]}
   );
   gpc606_5 gpc3303 (
      {stage1_42[156], stage1_42[157], stage1_42[158], stage1_42[159], stage1_42[160], stage1_42[161]},
      {stage1_44[120], stage1_44[121], stage1_44[122], stage1_44[123], stage1_44[124], stage1_44[125]},
      {stage2_46[20],stage2_45[24],stage2_44[30],stage2_43[43],stage2_42[52]}
   );
   gpc606_5 gpc3304 (
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[21],stage2_45[25],stage2_44[31],stage2_43[44]}
   );
   gpc615_5 gpc3305 (
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34]},
      {stage1_44[126]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[22],stage2_45[26],stage2_44[32],stage2_43[45]}
   );
   gpc615_5 gpc3306 (
      {stage1_43[35], stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39]},
      {stage1_44[127]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[23],stage2_45[27],stage2_44[33],stage2_43[46]}
   );
   gpc615_5 gpc3307 (
      {stage1_43[40], stage1_43[41], stage1_43[42], stage1_43[43], stage1_43[44]},
      {stage1_44[128]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[24],stage2_45[28],stage2_44[34],stage2_43[47]}
   );
   gpc615_5 gpc3308 (
      {stage1_43[45], stage1_43[46], stage1_43[47], stage1_43[48], stage1_43[49]},
      {stage1_44[129]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[25],stage2_45[29],stage2_44[35],stage2_43[48]}
   );
   gpc615_5 gpc3309 (
      {stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53], stage1_43[54]},
      {stage1_44[130]},
      {stage1_45[30], stage1_45[31], stage1_45[32], stage1_45[33], stage1_45[34], stage1_45[35]},
      {stage2_47[5],stage2_46[26],stage2_45[30],stage2_44[36],stage2_43[49]}
   );
   gpc615_5 gpc3310 (
      {stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage1_44[131]},
      {stage1_45[36], stage1_45[37], stage1_45[38], stage1_45[39], stage1_45[40], stage1_45[41]},
      {stage2_47[6],stage2_46[27],stage2_45[31],stage2_44[37],stage2_43[50]}
   );
   gpc615_5 gpc3311 (
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64]},
      {stage1_44[132]},
      {stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46], stage1_45[47]},
      {stage2_47[7],stage2_46[28],stage2_45[32],stage2_44[38],stage2_43[51]}
   );
   gpc615_5 gpc3312 (
      {stage1_43[65], stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69]},
      {stage1_44[133]},
      {stage1_45[48], stage1_45[49], stage1_45[50], stage1_45[51], stage1_45[52], stage1_45[53]},
      {stage2_47[8],stage2_46[29],stage2_45[33],stage2_44[39],stage2_43[52]}
   );
   gpc606_5 gpc3313 (
      {stage1_45[54], stage1_45[55], stage1_45[56], stage1_45[57], stage1_45[58], stage1_45[59]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[0],stage2_47[9],stage2_46[30],stage2_45[34]}
   );
   gpc606_5 gpc3314 (
      {stage1_45[60], stage1_45[61], stage1_45[62], stage1_45[63], stage1_45[64], stage1_45[65]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[1],stage2_47[10],stage2_46[31],stage2_45[35]}
   );
   gpc606_5 gpc3315 (
      {stage1_45[66], stage1_45[67], stage1_45[68], stage1_45[69], stage1_45[70], stage1_45[71]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[2],stage2_47[11],stage2_46[32],stage2_45[36]}
   );
   gpc606_5 gpc3316 (
      {stage1_45[72], stage1_45[73], stage1_45[74], stage1_45[75], stage1_45[76], stage1_45[77]},
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage2_49[3],stage2_48[3],stage2_47[12],stage2_46[33],stage2_45[37]}
   );
   gpc606_5 gpc3317 (
      {stage1_45[78], stage1_45[79], stage1_45[80], stage1_45[81], stage1_45[82], stage1_45[83]},
      {stage1_47[24], stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29]},
      {stage2_49[4],stage2_48[4],stage2_47[13],stage2_46[34],stage2_45[38]}
   );
   gpc606_5 gpc3318 (
      {stage1_45[84], stage1_45[85], stage1_45[86], stage1_45[87], stage1_45[88], stage1_45[89]},
      {stage1_47[30], stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35]},
      {stage2_49[5],stage2_48[5],stage2_47[14],stage2_46[35],stage2_45[39]}
   );
   gpc606_5 gpc3319 (
      {stage1_45[90], stage1_45[91], stage1_45[92], stage1_45[93], stage1_45[94], stage1_45[95]},
      {stage1_47[36], stage1_47[37], stage1_47[38], stage1_47[39], stage1_47[40], stage1_47[41]},
      {stage2_49[6],stage2_48[6],stage2_47[15],stage2_46[36],stage2_45[40]}
   );
   gpc606_5 gpc3320 (
      {stage1_45[96], stage1_45[97], stage1_45[98], stage1_45[99], stage1_45[100], stage1_45[101]},
      {stage1_47[42], stage1_47[43], stage1_47[44], stage1_47[45], stage1_47[46], stage1_47[47]},
      {stage2_49[7],stage2_48[7],stage2_47[16],stage2_46[37],stage2_45[41]}
   );
   gpc606_5 gpc3321 (
      {stage1_45[102], stage1_45[103], stage1_45[104], stage1_45[105], stage1_45[106], stage1_45[107]},
      {stage1_47[48], stage1_47[49], stage1_47[50], stage1_47[51], stage1_47[52], stage1_47[53]},
      {stage2_49[8],stage2_48[8],stage2_47[17],stage2_46[38],stage2_45[42]}
   );
   gpc606_5 gpc3322 (
      {stage1_45[108], stage1_45[109], stage1_45[110], stage1_45[111], stage1_45[112], stage1_45[113]},
      {stage1_47[54], stage1_47[55], stage1_47[56], stage1_47[57], stage1_47[58], stage1_47[59]},
      {stage2_49[9],stage2_48[9],stage2_47[18],stage2_46[39],stage2_45[43]}
   );
   gpc606_5 gpc3323 (
      {stage1_45[114], stage1_45[115], stage1_45[116], stage1_45[117], stage1_45[118], stage1_45[119]},
      {stage1_47[60], stage1_47[61], stage1_47[62], stage1_47[63], stage1_47[64], stage1_47[65]},
      {stage2_49[10],stage2_48[10],stage2_47[19],stage2_46[40],stage2_45[44]}
   );
   gpc606_5 gpc3324 (
      {stage1_45[120], stage1_45[121], stage1_45[122], stage1_45[123], stage1_45[124], stage1_45[125]},
      {stage1_47[66], stage1_47[67], stage1_47[68], stage1_47[69], stage1_47[70], stage1_47[71]},
      {stage2_49[11],stage2_48[11],stage2_47[20],stage2_46[41],stage2_45[45]}
   );
   gpc606_5 gpc3325 (
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[12],stage2_48[12],stage2_47[21],stage2_46[42]}
   );
   gpc606_5 gpc3326 (
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[13],stage2_48[13],stage2_47[22],stage2_46[43]}
   );
   gpc606_5 gpc3327 (
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], stage1_46[17]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[14],stage2_48[14],stage2_47[23],stage2_46[44]}
   );
   gpc606_5 gpc3328 (
      {stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21], stage1_46[22], stage1_46[23]},
      {stage1_48[18], stage1_48[19], stage1_48[20], stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage2_50[3],stage2_49[15],stage2_48[15],stage2_47[24],stage2_46[45]}
   );
   gpc606_5 gpc3329 (
      {stage1_46[24], stage1_46[25], stage1_46[26], stage1_46[27], stage1_46[28], stage1_46[29]},
      {stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27], stage1_48[28], stage1_48[29]},
      {stage2_50[4],stage2_49[16],stage2_48[16],stage2_47[25],stage2_46[46]}
   );
   gpc606_5 gpc3330 (
      {stage1_46[30], stage1_46[31], stage1_46[32], stage1_46[33], stage1_46[34], stage1_46[35]},
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage2_50[5],stage2_49[17],stage2_48[17],stage2_47[26],stage2_46[47]}
   );
   gpc606_5 gpc3331 (
      {stage1_46[36], stage1_46[37], stage1_46[38], stage1_46[39], stage1_46[40], stage1_46[41]},
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage2_50[6],stage2_49[18],stage2_48[18],stage2_47[27],stage2_46[48]}
   );
   gpc606_5 gpc3332 (
      {stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45], stage1_46[46], stage1_46[47]},
      {stage1_48[42], stage1_48[43], stage1_48[44], stage1_48[45], stage1_48[46], stage1_48[47]},
      {stage2_50[7],stage2_49[19],stage2_48[19],stage2_47[28],stage2_46[49]}
   );
   gpc606_5 gpc3333 (
      {stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51], stage1_46[52], stage1_46[53]},
      {stage1_48[48], stage1_48[49], stage1_48[50], stage1_48[51], stage1_48[52], stage1_48[53]},
      {stage2_50[8],stage2_49[20],stage2_48[20],stage2_47[29],stage2_46[50]}
   );
   gpc606_5 gpc3334 (
      {stage1_46[54], stage1_46[55], stage1_46[56], stage1_46[57], stage1_46[58], stage1_46[59]},
      {stage1_48[54], stage1_48[55], stage1_48[56], stage1_48[57], stage1_48[58], stage1_48[59]},
      {stage2_50[9],stage2_49[21],stage2_48[21],stage2_47[30],stage2_46[51]}
   );
   gpc606_5 gpc3335 (
      {stage1_46[60], stage1_46[61], stage1_46[62], stage1_46[63], stage1_46[64], stage1_46[65]},
      {stage1_48[60], stage1_48[61], stage1_48[62], stage1_48[63], stage1_48[64], stage1_48[65]},
      {stage2_50[10],stage2_49[22],stage2_48[22],stage2_47[31],stage2_46[52]}
   );
   gpc606_5 gpc3336 (
      {stage1_46[66], stage1_46[67], stage1_46[68], stage1_46[69], stage1_46[70], stage1_46[71]},
      {stage1_48[66], stage1_48[67], stage1_48[68], stage1_48[69], stage1_48[70], stage1_48[71]},
      {stage2_50[11],stage2_49[23],stage2_48[23],stage2_47[32],stage2_46[53]}
   );
   gpc606_5 gpc3337 (
      {stage1_46[72], stage1_46[73], stage1_46[74], stage1_46[75], stage1_46[76], stage1_46[77]},
      {stage1_48[72], stage1_48[73], stage1_48[74], stage1_48[75], stage1_48[76], stage1_48[77]},
      {stage2_50[12],stage2_49[24],stage2_48[24],stage2_47[33],stage2_46[54]}
   );
   gpc606_5 gpc3338 (
      {stage1_46[78], stage1_46[79], stage1_46[80], stage1_46[81], stage1_46[82], stage1_46[83]},
      {stage1_48[78], stage1_48[79], stage1_48[80], stage1_48[81], stage1_48[82], stage1_48[83]},
      {stage2_50[13],stage2_49[25],stage2_48[25],stage2_47[34],stage2_46[55]}
   );
   gpc606_5 gpc3339 (
      {stage1_46[84], stage1_46[85], stage1_46[86], stage1_46[87], stage1_46[88], stage1_46[89]},
      {stage1_48[84], stage1_48[85], stage1_48[86], stage1_48[87], stage1_48[88], stage1_48[89]},
      {stage2_50[14],stage2_49[26],stage2_48[26],stage2_47[35],stage2_46[56]}
   );
   gpc606_5 gpc3340 (
      {stage1_46[90], stage1_46[91], stage1_46[92], stage1_46[93], stage1_46[94], stage1_46[95]},
      {stage1_48[90], stage1_48[91], stage1_48[92], stage1_48[93], stage1_48[94], stage1_48[95]},
      {stage2_50[15],stage2_49[27],stage2_48[27],stage2_47[36],stage2_46[57]}
   );
   gpc606_5 gpc3341 (
      {stage1_47[72], stage1_47[73], stage1_47[74], stage1_47[75], stage1_47[76], stage1_47[77]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[16],stage2_49[28],stage2_48[28],stage2_47[37]}
   );
   gpc606_5 gpc3342 (
      {stage1_47[78], stage1_47[79], stage1_47[80], stage1_47[81], stage1_47[82], stage1_47[83]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[17],stage2_49[29],stage2_48[29],stage2_47[38]}
   );
   gpc606_5 gpc3343 (
      {stage1_47[84], stage1_47[85], stage1_47[86], stage1_47[87], stage1_47[88], stage1_47[89]},
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage2_51[2],stage2_50[18],stage2_49[30],stage2_48[30],stage2_47[39]}
   );
   gpc606_5 gpc3344 (
      {stage1_47[90], stage1_47[91], stage1_47[92], stage1_47[93], stage1_47[94], stage1_47[95]},
      {stage1_49[18], stage1_49[19], stage1_49[20], stage1_49[21], stage1_49[22], stage1_49[23]},
      {stage2_51[3],stage2_50[19],stage2_49[31],stage2_48[31],stage2_47[40]}
   );
   gpc623_5 gpc3345 (
      {stage1_47[96], stage1_47[97], stage1_47[98]},
      {stage1_48[96], stage1_48[97]},
      {stage1_49[24], stage1_49[25], stage1_49[26], stage1_49[27], stage1_49[28], stage1_49[29]},
      {stage2_51[4],stage2_50[20],stage2_49[32],stage2_48[32],stage2_47[41]}
   );
   gpc623_5 gpc3346 (
      {stage1_47[99], stage1_47[100], stage1_47[101]},
      {stage1_48[98], stage1_48[99]},
      {stage1_49[30], stage1_49[31], stage1_49[32], stage1_49[33], stage1_49[34], stage1_49[35]},
      {stage2_51[5],stage2_50[21],stage2_49[33],stage2_48[33],stage2_47[42]}
   );
   gpc1406_5 gpc3347 (
      {stage1_49[36], stage1_49[37], stage1_49[38], stage1_49[39], stage1_49[40], stage1_49[41]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3]},
      {stage1_52[0]},
      {stage2_53[0],stage2_52[0],stage2_51[6],stage2_50[22],stage2_49[34]}
   );
   gpc606_5 gpc3348 (
      {stage1_49[42], stage1_49[43], stage1_49[44], stage1_49[45], stage1_49[46], stage1_49[47]},
      {stage1_51[4], stage1_51[5], stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9]},
      {stage2_53[1],stage2_52[1],stage2_51[7],stage2_50[23],stage2_49[35]}
   );
   gpc606_5 gpc3349 (
      {stage1_49[48], stage1_49[49], stage1_49[50], stage1_49[51], stage1_49[52], stage1_49[53]},
      {stage1_51[10], stage1_51[11], stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15]},
      {stage2_53[2],stage2_52[2],stage2_51[8],stage2_50[24],stage2_49[36]}
   );
   gpc606_5 gpc3350 (
      {stage1_49[54], stage1_49[55], stage1_49[56], stage1_49[57], stage1_49[58], stage1_49[59]},
      {stage1_51[16], stage1_51[17], stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21]},
      {stage2_53[3],stage2_52[3],stage2_51[9],stage2_50[25],stage2_49[37]}
   );
   gpc606_5 gpc3351 (
      {stage1_49[60], stage1_49[61], stage1_49[62], stage1_49[63], stage1_49[64], stage1_49[65]},
      {stage1_51[22], stage1_51[23], stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27]},
      {stage2_53[4],stage2_52[4],stage2_51[10],stage2_50[26],stage2_49[38]}
   );
   gpc606_5 gpc3352 (
      {stage1_49[66], stage1_49[67], stage1_49[68], stage1_49[69], stage1_49[70], stage1_49[71]},
      {stage1_51[28], stage1_51[29], stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33]},
      {stage2_53[5],stage2_52[5],stage2_51[11],stage2_50[27],stage2_49[39]}
   );
   gpc606_5 gpc3353 (
      {stage1_49[72], stage1_49[73], stage1_49[74], stage1_49[75], stage1_49[76], stage1_49[77]},
      {stage1_51[34], stage1_51[35], stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39]},
      {stage2_53[6],stage2_52[6],stage2_51[12],stage2_50[28],stage2_49[40]}
   );
   gpc615_5 gpc3354 (
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4]},
      {stage1_51[40]},
      {stage1_52[1], stage1_52[2], stage1_52[3], stage1_52[4], stage1_52[5], stage1_52[6]},
      {stage2_54[0],stage2_53[7],stage2_52[7],stage2_51[13],stage2_50[29]}
   );
   gpc615_5 gpc3355 (
      {stage1_50[5], stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9]},
      {stage1_51[41]},
      {stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10], stage1_52[11], stage1_52[12]},
      {stage2_54[1],stage2_53[8],stage2_52[8],stage2_51[14],stage2_50[30]}
   );
   gpc615_5 gpc3356 (
      {stage1_50[10], stage1_50[11], stage1_50[12], stage1_50[13], stage1_50[14]},
      {stage1_51[42]},
      {stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16], stage1_52[17], stage1_52[18]},
      {stage2_54[2],stage2_53[9],stage2_52[9],stage2_51[15],stage2_50[31]}
   );
   gpc615_5 gpc3357 (
      {stage1_50[15], stage1_50[16], stage1_50[17], stage1_50[18], stage1_50[19]},
      {stage1_51[43]},
      {stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22], stage1_52[23], stage1_52[24]},
      {stage2_54[3],stage2_53[10],stage2_52[10],stage2_51[16],stage2_50[32]}
   );
   gpc615_5 gpc3358 (
      {stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23], stage1_50[24]},
      {stage1_51[44]},
      {stage1_52[25], stage1_52[26], stage1_52[27], stage1_52[28], stage1_52[29], stage1_52[30]},
      {stage2_54[4],stage2_53[11],stage2_52[11],stage2_51[17],stage2_50[33]}
   );
   gpc615_5 gpc3359 (
      {stage1_50[25], stage1_50[26], stage1_50[27], stage1_50[28], stage1_50[29]},
      {stage1_51[45]},
      {stage1_52[31], stage1_52[32], stage1_52[33], stage1_52[34], stage1_52[35], stage1_52[36]},
      {stage2_54[5],stage2_53[12],stage2_52[12],stage2_51[18],stage2_50[34]}
   );
   gpc615_5 gpc3360 (
      {stage1_50[30], stage1_50[31], stage1_50[32], stage1_50[33], stage1_50[34]},
      {stage1_51[46]},
      {stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41], stage1_52[42]},
      {stage2_54[6],stage2_53[13],stage2_52[13],stage2_51[19],stage2_50[35]}
   );
   gpc615_5 gpc3361 (
      {stage1_50[35], stage1_50[36], stage1_50[37], stage1_50[38], stage1_50[39]},
      {stage1_51[47]},
      {stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46], stage1_52[47], stage1_52[48]},
      {stage2_54[7],stage2_53[14],stage2_52[14],stage2_51[20],stage2_50[36]}
   );
   gpc615_5 gpc3362 (
      {stage1_50[40], stage1_50[41], stage1_50[42], stage1_50[43], stage1_50[44]},
      {stage1_51[48]},
      {stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52], stage1_52[53], stage1_52[54]},
      {stage2_54[8],stage2_53[15],stage2_52[15],stage2_51[21],stage2_50[37]}
   );
   gpc615_5 gpc3363 (
      {stage1_50[45], stage1_50[46], stage1_50[47], stage1_50[48], stage1_50[49]},
      {stage1_51[49]},
      {stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58], stage1_52[59], stage1_52[60]},
      {stage2_54[9],stage2_53[16],stage2_52[16],stage2_51[22],stage2_50[38]}
   );
   gpc615_5 gpc3364 (
      {stage1_50[50], stage1_50[51], stage1_50[52], stage1_50[53], stage1_50[54]},
      {stage1_51[50]},
      {stage1_52[61], stage1_52[62], stage1_52[63], stage1_52[64], stage1_52[65], stage1_52[66]},
      {stage2_54[10],stage2_53[17],stage2_52[17],stage2_51[23],stage2_50[39]}
   );
   gpc615_5 gpc3365 (
      {stage1_50[55], stage1_50[56], stage1_50[57], stage1_50[58], stage1_50[59]},
      {stage1_51[51]},
      {stage1_52[67], stage1_52[68], stage1_52[69], stage1_52[70], stage1_52[71], stage1_52[72]},
      {stage2_54[11],stage2_53[18],stage2_52[18],stage2_51[24],stage2_50[40]}
   );
   gpc615_5 gpc3366 (
      {stage1_50[60], stage1_50[61], stage1_50[62], stage1_50[63], stage1_50[64]},
      {stage1_51[52]},
      {stage1_52[73], stage1_52[74], stage1_52[75], stage1_52[76], stage1_52[77], stage1_52[78]},
      {stage2_54[12],stage2_53[19],stage2_52[19],stage2_51[25],stage2_50[41]}
   );
   gpc615_5 gpc3367 (
      {stage1_50[65], stage1_50[66], stage1_50[67], stage1_50[68], stage1_50[69]},
      {stage1_51[53]},
      {stage1_52[79], stage1_52[80], stage1_52[81], stage1_52[82], stage1_52[83], stage1_52[84]},
      {stage2_54[13],stage2_53[20],stage2_52[20],stage2_51[26],stage2_50[42]}
   );
   gpc615_5 gpc3368 (
      {stage1_50[70], stage1_50[71], stage1_50[72], stage1_50[73], stage1_50[74]},
      {stage1_51[54]},
      {stage1_52[85], stage1_52[86], stage1_52[87], stage1_52[88], stage1_52[89], stage1_52[90]},
      {stage2_54[14],stage2_53[21],stage2_52[21],stage2_51[27],stage2_50[43]}
   );
   gpc615_5 gpc3369 (
      {stage1_52[91], stage1_52[92], stage1_52[93], stage1_52[94], stage1_52[95]},
      {stage1_53[0]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[0],stage2_54[15],stage2_53[22],stage2_52[22]}
   );
   gpc615_5 gpc3370 (
      {stage1_52[96], stage1_52[97], stage1_52[98], stage1_52[99], stage1_52[100]},
      {stage1_53[1]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[1],stage2_54[16],stage2_53[23],stage2_52[23]}
   );
   gpc615_5 gpc3371 (
      {stage1_52[101], stage1_52[102], stage1_52[103], stage1_52[104], stage1_52[105]},
      {stage1_53[2]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[2],stage2_54[17],stage2_53[24],stage2_52[24]}
   );
   gpc615_5 gpc3372 (
      {stage1_52[106], stage1_52[107], stage1_52[108], stage1_52[109], stage1_52[110]},
      {stage1_53[3]},
      {stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21], stage1_54[22], stage1_54[23]},
      {stage2_56[3],stage2_55[3],stage2_54[18],stage2_53[25],stage2_52[25]}
   );
   gpc615_5 gpc3373 (
      {stage1_52[111], stage1_52[112], stage1_52[113], stage1_52[114], stage1_52[115]},
      {stage1_53[4]},
      {stage1_54[24], stage1_54[25], stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29]},
      {stage2_56[4],stage2_55[4],stage2_54[19],stage2_53[26],stage2_52[26]}
   );
   gpc615_5 gpc3374 (
      {stage1_53[5], stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9]},
      {stage1_54[30]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[5],stage2_55[5],stage2_54[20],stage2_53[27]}
   );
   gpc615_5 gpc3375 (
      {stage1_53[10], stage1_53[11], stage1_53[12], stage1_53[13], stage1_53[14]},
      {stage1_54[31]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage2_57[1],stage2_56[6],stage2_55[6],stage2_54[21],stage2_53[28]}
   );
   gpc615_5 gpc3376 (
      {stage1_53[15], stage1_53[16], stage1_53[17], stage1_53[18], stage1_53[19]},
      {stage1_54[32]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage2_57[2],stage2_56[7],stage2_55[7],stage2_54[22],stage2_53[29]}
   );
   gpc615_5 gpc3377 (
      {stage1_53[20], stage1_53[21], stage1_53[22], stage1_53[23], stage1_53[24]},
      {stage1_54[33]},
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22], stage1_55[23]},
      {stage2_57[3],stage2_56[8],stage2_55[8],stage2_54[23],stage2_53[30]}
   );
   gpc615_5 gpc3378 (
      {stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28], stage1_53[29]},
      {stage1_54[34]},
      {stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27], stage1_55[28], stage1_55[29]},
      {stage2_57[4],stage2_56[9],stage2_55[9],stage2_54[24],stage2_53[31]}
   );
   gpc615_5 gpc3379 (
      {stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34]},
      {stage1_54[35]},
      {stage1_55[30], stage1_55[31], stage1_55[32], stage1_55[33], stage1_55[34], stage1_55[35]},
      {stage2_57[5],stage2_56[10],stage2_55[10],stage2_54[25],stage2_53[32]}
   );
   gpc615_5 gpc3380 (
      {stage1_53[35], stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39]},
      {stage1_54[36]},
      {stage1_55[36], stage1_55[37], stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41]},
      {stage2_57[6],stage2_56[11],stage2_55[11],stage2_54[26],stage2_53[33]}
   );
   gpc615_5 gpc3381 (
      {stage1_53[40], stage1_53[41], stage1_53[42], stage1_53[43], stage1_53[44]},
      {stage1_54[37]},
      {stage1_55[42], stage1_55[43], stage1_55[44], stage1_55[45], stage1_55[46], stage1_55[47]},
      {stage2_57[7],stage2_56[12],stage2_55[12],stage2_54[27],stage2_53[34]}
   );
   gpc615_5 gpc3382 (
      {stage1_53[45], stage1_53[46], stage1_53[47], stage1_53[48], stage1_53[49]},
      {stage1_54[38]},
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52], stage1_55[53]},
      {stage2_57[8],stage2_56[13],stage2_55[13],stage2_54[28],stage2_53[35]}
   );
   gpc615_5 gpc3383 (
      {stage1_53[50], stage1_53[51], stage1_53[52], stage1_53[53], stage1_53[54]},
      {stage1_54[39]},
      {stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57], stage1_55[58], stage1_55[59]},
      {stage2_57[9],stage2_56[14],stage2_55[14],stage2_54[29],stage2_53[36]}
   );
   gpc615_5 gpc3384 (
      {stage1_53[55], stage1_53[56], stage1_53[57], stage1_53[58], stage1_53[59]},
      {stage1_54[40]},
      {stage1_55[60], stage1_55[61], stage1_55[62], stage1_55[63], stage1_55[64], stage1_55[65]},
      {stage2_57[10],stage2_56[15],stage2_55[15],stage2_54[30],stage2_53[37]}
   );
   gpc615_5 gpc3385 (
      {stage1_53[60], stage1_53[61], stage1_53[62], stage1_53[63], stage1_53[64]},
      {stage1_54[41]},
      {stage1_55[66], stage1_55[67], stage1_55[68], stage1_55[69], stage1_55[70], stage1_55[71]},
      {stage2_57[11],stage2_56[16],stage2_55[16],stage2_54[31],stage2_53[38]}
   );
   gpc615_5 gpc3386 (
      {stage1_53[65], stage1_53[66], stage1_53[67], stage1_53[68], stage1_53[69]},
      {stage1_54[42]},
      {stage1_55[72], stage1_55[73], stage1_55[74], stage1_55[75], stage1_55[76], stage1_55[77]},
      {stage2_57[12],stage2_56[17],stage2_55[17],stage2_54[32],stage2_53[39]}
   );
   gpc606_5 gpc3387 (
      {stage1_54[43], stage1_54[44], stage1_54[45], stage1_54[46], stage1_54[47], stage1_54[48]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[13],stage2_56[18],stage2_55[18],stage2_54[33]}
   );
   gpc606_5 gpc3388 (
      {stage1_54[49], stage1_54[50], stage1_54[51], stage1_54[52], stage1_54[53], stage1_54[54]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[14],stage2_56[19],stage2_55[19],stage2_54[34]}
   );
   gpc606_5 gpc3389 (
      {stage1_54[55], stage1_54[56], stage1_54[57], stage1_54[58], stage1_54[59], stage1_54[60]},
      {stage1_56[12], stage1_56[13], stage1_56[14], stage1_56[15], stage1_56[16], stage1_56[17]},
      {stage2_58[2],stage2_57[15],stage2_56[20],stage2_55[20],stage2_54[35]}
   );
   gpc606_5 gpc3390 (
      {stage1_54[61], stage1_54[62], stage1_54[63], stage1_54[64], stage1_54[65], stage1_54[66]},
      {stage1_56[18], stage1_56[19], stage1_56[20], stage1_56[21], stage1_56[22], stage1_56[23]},
      {stage2_58[3],stage2_57[16],stage2_56[21],stage2_55[21],stage2_54[36]}
   );
   gpc606_5 gpc3391 (
      {stage1_54[67], stage1_54[68], stage1_54[69], stage1_54[70], stage1_54[71], stage1_54[72]},
      {stage1_56[24], stage1_56[25], stage1_56[26], stage1_56[27], stage1_56[28], stage1_56[29]},
      {stage2_58[4],stage2_57[17],stage2_56[22],stage2_55[22],stage2_54[37]}
   );
   gpc606_5 gpc3392 (
      {stage1_54[73], stage1_54[74], stage1_54[75], stage1_54[76], stage1_54[77], stage1_54[78]},
      {stage1_56[30], stage1_56[31], stage1_56[32], stage1_56[33], stage1_56[34], stage1_56[35]},
      {stage2_58[5],stage2_57[18],stage2_56[23],stage2_55[23],stage2_54[38]}
   );
   gpc606_5 gpc3393 (
      {stage1_54[79], stage1_54[80], stage1_54[81], stage1_54[82], stage1_54[83], stage1_54[84]},
      {stage1_56[36], stage1_56[37], stage1_56[38], stage1_56[39], stage1_56[40], stage1_56[41]},
      {stage2_58[6],stage2_57[19],stage2_56[24],stage2_55[24],stage2_54[39]}
   );
   gpc606_5 gpc3394 (
      {stage1_54[85], stage1_54[86], stage1_54[87], stage1_54[88], stage1_54[89], stage1_54[90]},
      {stage1_56[42], stage1_56[43], stage1_56[44], stage1_56[45], stage1_56[46], stage1_56[47]},
      {stage2_58[7],stage2_57[20],stage2_56[25],stage2_55[25],stage2_54[40]}
   );
   gpc606_5 gpc3395 (
      {stage1_54[91], stage1_54[92], stage1_54[93], stage1_54[94], stage1_54[95], stage1_54[96]},
      {stage1_56[48], stage1_56[49], stage1_56[50], stage1_56[51], stage1_56[52], stage1_56[53]},
      {stage2_58[8],stage2_57[21],stage2_56[26],stage2_55[26],stage2_54[41]}
   );
   gpc606_5 gpc3396 (
      {stage1_54[97], stage1_54[98], stage1_54[99], stage1_54[100], stage1_54[101], stage1_54[102]},
      {stage1_56[54], stage1_56[55], stage1_56[56], stage1_56[57], stage1_56[58], stage1_56[59]},
      {stage2_58[9],stage2_57[22],stage2_56[27],stage2_55[27],stage2_54[42]}
   );
   gpc606_5 gpc3397 (
      {stage1_54[103], stage1_54[104], stage1_54[105], stage1_54[106], stage1_54[107], stage1_54[108]},
      {stage1_56[60], stage1_56[61], stage1_56[62], stage1_56[63], stage1_56[64], stage1_56[65]},
      {stage2_58[10],stage2_57[23],stage2_56[28],stage2_55[28],stage2_54[43]}
   );
   gpc606_5 gpc3398 (
      {stage1_54[109], stage1_54[110], stage1_54[111], stage1_54[112], stage1_54[113], stage1_54[114]},
      {stage1_56[66], stage1_56[67], stage1_56[68], stage1_56[69], stage1_56[70], stage1_56[71]},
      {stage2_58[11],stage2_57[24],stage2_56[29],stage2_55[29],stage2_54[44]}
   );
   gpc606_5 gpc3399 (
      {stage1_54[115], stage1_54[116], stage1_54[117], stage1_54[118], stage1_54[119], stage1_54[120]},
      {stage1_56[72], stage1_56[73], stage1_56[74], stage1_56[75], stage1_56[76], stage1_56[77]},
      {stage2_58[12],stage2_57[25],stage2_56[30],stage2_55[30],stage2_54[45]}
   );
   gpc606_5 gpc3400 (
      {stage1_54[121], stage1_54[122], stage1_54[123], stage1_54[124], stage1_54[125], stage1_54[126]},
      {stage1_56[78], stage1_56[79], stage1_56[80], stage1_56[81], stage1_56[82], stage1_56[83]},
      {stage2_58[13],stage2_57[26],stage2_56[31],stage2_55[31],stage2_54[46]}
   );
   gpc606_5 gpc3401 (
      {stage1_54[127], stage1_54[128], stage1_54[129], stage1_54[130], stage1_54[131], stage1_54[132]},
      {stage1_56[84], stage1_56[85], stage1_56[86], stage1_56[87], stage1_56[88], stage1_56[89]},
      {stage2_58[14],stage2_57[27],stage2_56[32],stage2_55[32],stage2_54[47]}
   );
   gpc606_5 gpc3402 (
      {stage1_55[78], stage1_55[79], stage1_55[80], stage1_55[81], stage1_55[82], stage1_55[83]},
      {stage1_57[0], stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage2_59[0],stage2_58[15],stage2_57[28],stage2_56[33],stage2_55[33]}
   );
   gpc606_5 gpc3403 (
      {stage1_55[84], stage1_55[85], stage1_55[86], stage1_55[87], stage1_55[88], stage1_55[89]},
      {stage1_57[6], stage1_57[7], stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11]},
      {stage2_59[1],stage2_58[16],stage2_57[29],stage2_56[34],stage2_55[34]}
   );
   gpc606_5 gpc3404 (
      {stage1_56[90], stage1_56[91], stage1_56[92], stage1_56[93], stage1_56[94], stage1_56[95]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[2],stage2_58[17],stage2_57[30],stage2_56[35]}
   );
   gpc606_5 gpc3405 (
      {stage1_56[96], stage1_56[97], stage1_56[98], stage1_56[99], stage1_56[100], stage1_56[101]},
      {stage1_58[6], stage1_58[7], stage1_58[8], stage1_58[9], stage1_58[10], stage1_58[11]},
      {stage2_60[1],stage2_59[3],stage2_58[18],stage2_57[31],stage2_56[36]}
   );
   gpc606_5 gpc3406 (
      {stage1_56[102], stage1_56[103], stage1_56[104], stage1_56[105], stage1_56[106], stage1_56[107]},
      {stage1_58[12], stage1_58[13], stage1_58[14], stage1_58[15], stage1_58[16], stage1_58[17]},
      {stage2_60[2],stage2_59[4],stage2_58[19],stage2_57[32],stage2_56[37]}
   );
   gpc606_5 gpc3407 (
      {stage1_56[108], stage1_56[109], stage1_56[110], stage1_56[111], stage1_56[112], stage1_56[113]},
      {stage1_58[18], stage1_58[19], stage1_58[20], stage1_58[21], stage1_58[22], stage1_58[23]},
      {stage2_60[3],stage2_59[5],stage2_58[20],stage2_57[33],stage2_56[38]}
   );
   gpc606_5 gpc3408 (
      {stage1_56[114], stage1_56[115], stage1_56[116], stage1_56[117], stage1_56[118], stage1_56[119]},
      {stage1_58[24], stage1_58[25], stage1_58[26], stage1_58[27], stage1_58[28], stage1_58[29]},
      {stage2_60[4],stage2_59[6],stage2_58[21],stage2_57[34],stage2_56[39]}
   );
   gpc606_5 gpc3409 (
      {stage1_56[120], stage1_56[121], stage1_56[122], stage1_56[123], stage1_56[124], stage1_56[125]},
      {stage1_58[30], stage1_58[31], stage1_58[32], stage1_58[33], stage1_58[34], stage1_58[35]},
      {stage2_60[5],stage2_59[7],stage2_58[22],stage2_57[35],stage2_56[40]}
   );
   gpc606_5 gpc3410 (
      {stage1_56[126], stage1_56[127], stage1_56[128], stage1_56[129], stage1_56[130], stage1_56[131]},
      {stage1_58[36], stage1_58[37], stage1_58[38], stage1_58[39], stage1_58[40], stage1_58[41]},
      {stage2_60[6],stage2_59[8],stage2_58[23],stage2_57[36],stage2_56[41]}
   );
   gpc606_5 gpc3411 (
      {stage1_56[132], stage1_56[133], stage1_56[134], stage1_56[135], stage1_56[136], stage1_56[137]},
      {stage1_58[42], stage1_58[43], stage1_58[44], stage1_58[45], stage1_58[46], stage1_58[47]},
      {stage2_60[7],stage2_59[9],stage2_58[24],stage2_57[37],stage2_56[42]}
   );
   gpc606_5 gpc3412 (
      {stage1_56[138], stage1_56[139], stage1_56[140], stage1_56[141], stage1_56[142], stage1_56[143]},
      {stage1_58[48], stage1_58[49], stage1_58[50], stage1_58[51], stage1_58[52], stage1_58[53]},
      {stage2_60[8],stage2_59[10],stage2_58[25],stage2_57[38],stage2_56[43]}
   );
   gpc606_5 gpc3413 (
      {stage1_56[144], stage1_56[145], stage1_56[146], stage1_56[147], stage1_56[148], stage1_56[149]},
      {stage1_58[54], stage1_58[55], stage1_58[56], stage1_58[57], stage1_58[58], stage1_58[59]},
      {stage2_60[9],stage2_59[11],stage2_58[26],stage2_57[39],stage2_56[44]}
   );
   gpc606_5 gpc3414 (
      {stage1_57[12], stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[10],stage2_59[12],stage2_58[27],stage2_57[40]}
   );
   gpc606_5 gpc3415 (
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[11],stage2_59[13],stage2_58[28],stage2_57[41]}
   );
   gpc606_5 gpc3416 (
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17]},
      {stage2_61[2],stage2_60[12],stage2_59[14],stage2_58[29],stage2_57[42]}
   );
   gpc606_5 gpc3417 (
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage1_59[18], stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23]},
      {stage2_61[3],stage2_60[13],stage2_59[15],stage2_58[30],stage2_57[43]}
   );
   gpc606_5 gpc3418 (
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage1_59[24], stage1_59[25], stage1_59[26], stage1_59[27], stage1_59[28], stage1_59[29]},
      {stage2_61[4],stage2_60[14],stage2_59[16],stage2_58[31],stage2_57[44]}
   );
   gpc606_5 gpc3419 (
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage1_59[30], stage1_59[31], stage1_59[32], stage1_59[33], stage1_59[34], stage1_59[35]},
      {stage2_61[5],stage2_60[15],stage2_59[17],stage2_58[32],stage2_57[45]}
   );
   gpc606_5 gpc3420 (
      {stage1_57[48], stage1_57[49], stage1_57[50], stage1_57[51], stage1_57[52], stage1_57[53]},
      {stage1_59[36], stage1_59[37], stage1_59[38], stage1_59[39], stage1_59[40], stage1_59[41]},
      {stage2_61[6],stage2_60[16],stage2_59[18],stage2_58[33],stage2_57[46]}
   );
   gpc606_5 gpc3421 (
      {stage1_57[54], stage1_57[55], stage1_57[56], stage1_57[57], stage1_57[58], stage1_57[59]},
      {stage1_59[42], stage1_59[43], stage1_59[44], stage1_59[45], stage1_59[46], stage1_59[47]},
      {stage2_61[7],stage2_60[17],stage2_59[19],stage2_58[34],stage2_57[47]}
   );
   gpc606_5 gpc3422 (
      {stage1_57[60], stage1_57[61], stage1_57[62], stage1_57[63], stage1_57[64], stage1_57[65]},
      {stage1_59[48], stage1_59[49], stage1_59[50], stage1_59[51], stage1_59[52], stage1_59[53]},
      {stage2_61[8],stage2_60[18],stage2_59[20],stage2_58[35],stage2_57[48]}
   );
   gpc606_5 gpc3423 (
      {stage1_57[66], stage1_57[67], stage1_57[68], stage1_57[69], stage1_57[70], stage1_57[71]},
      {stage1_59[54], stage1_59[55], stage1_59[56], stage1_59[57], stage1_59[58], stage1_59[59]},
      {stage2_61[9],stage2_60[19],stage2_59[21],stage2_58[36],stage2_57[49]}
   );
   gpc606_5 gpc3424 (
      {stage1_58[60], stage1_58[61], stage1_58[62], stage1_58[63], stage1_58[64], stage1_58[65]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[10],stage2_60[20],stage2_59[22],stage2_58[37]}
   );
   gpc606_5 gpc3425 (
      {stage1_58[66], stage1_58[67], stage1_58[68], stage1_58[69], stage1_58[70], stage1_58[71]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[11],stage2_60[21],stage2_59[23],stage2_58[38]}
   );
   gpc606_5 gpc3426 (
      {stage1_58[72], stage1_58[73], stage1_58[74], stage1_58[75], stage1_58[76], stage1_58[77]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[12],stage2_60[22],stage2_59[24],stage2_58[39]}
   );
   gpc606_5 gpc3427 (
      {stage1_59[60], stage1_59[61], stage1_59[62], stage1_59[63], stage1_59[64], stage1_59[65]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[3],stage2_61[13],stage2_60[23],stage2_59[25]}
   );
   gpc606_5 gpc3428 (
      {stage1_59[66], stage1_59[67], stage1_59[68], stage1_59[69], stage1_59[70], stage1_59[71]},
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage2_63[1],stage2_62[4],stage2_61[14],stage2_60[24],stage2_59[26]}
   );
   gpc606_5 gpc3429 (
      {stage1_59[72], stage1_59[73], stage1_59[74], stage1_59[75], stage1_59[76], stage1_59[77]},
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage2_63[2],stage2_62[5],stage2_61[15],stage2_60[25],stage2_59[27]}
   );
   gpc606_5 gpc3430 (
      {stage1_59[78], stage1_59[79], stage1_59[80], stage1_59[81], stage1_59[82], stage1_59[83]},
      {stage1_61[18], stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23]},
      {stage2_63[3],stage2_62[6],stage2_61[16],stage2_60[26],stage2_59[28]}
   );
   gpc606_5 gpc3431 (
      {stage1_59[84], stage1_59[85], stage1_59[86], stage1_59[87], stage1_59[88], stage1_59[89]},
      {stage1_61[24], stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29]},
      {stage2_63[4],stage2_62[7],stage2_61[17],stage2_60[27],stage2_59[29]}
   );
   gpc606_5 gpc3432 (
      {stage1_59[90], stage1_59[91], stage1_59[92], stage1_59[93], stage1_59[94], stage1_59[95]},
      {stage1_61[30], stage1_61[31], stage1_61[32], stage1_61[33], stage1_61[34], stage1_61[35]},
      {stage2_63[5],stage2_62[8],stage2_61[18],stage2_60[28],stage2_59[30]}
   );
   gpc606_5 gpc3433 (
      {stage1_59[96], stage1_59[97], stage1_59[98], stage1_59[99], stage1_59[100], stage1_59[101]},
      {stage1_61[36], stage1_61[37], stage1_61[38], stage1_61[39], stage1_61[40], stage1_61[41]},
      {stage2_63[6],stage2_62[9],stage2_61[19],stage2_60[29],stage2_59[31]}
   );
   gpc606_5 gpc3434 (
      {stage1_59[102], stage1_59[103], stage1_59[104], stage1_59[105], stage1_59[106], stage1_59[107]},
      {stage1_61[42], stage1_61[43], stage1_61[44], stage1_61[45], stage1_61[46], stage1_61[47]},
      {stage2_63[7],stage2_62[10],stage2_61[20],stage2_60[30],stage2_59[32]}
   );
   gpc606_5 gpc3435 (
      {stage1_59[108], stage1_59[109], stage1_59[110], stage1_59[111], stage1_59[112], stage1_59[113]},
      {stage1_61[48], stage1_61[49], stage1_61[50], stage1_61[51], stage1_61[52], stage1_61[53]},
      {stage2_63[8],stage2_62[11],stage2_61[21],stage2_60[31],stage2_59[33]}
   );
   gpc606_5 gpc3436 (
      {stage1_59[114], stage1_59[115], stage1_59[116], stage1_59[117], stage1_59[118], stage1_59[119]},
      {stage1_61[54], stage1_61[55], stage1_61[56], stage1_61[57], stage1_61[58], stage1_61[59]},
      {stage2_63[9],stage2_62[12],stage2_61[22],stage2_60[32],stage2_59[34]}
   );
   gpc606_5 gpc3437 (
      {stage1_59[120], stage1_59[121], stage1_59[122], stage1_59[123], stage1_59[124], stage1_59[125]},
      {stage1_61[60], stage1_61[61], stage1_61[62], stage1_61[63], stage1_61[64], stage1_61[65]},
      {stage2_63[10],stage2_62[13],stage2_61[23],stage2_60[33],stage2_59[35]}
   );
   gpc606_5 gpc3438 (
      {stage1_59[126], stage1_59[127], stage1_59[128], stage1_59[129], stage1_59[130], stage1_59[131]},
      {stage1_61[66], stage1_61[67], stage1_61[68], stage1_61[69], stage1_61[70], stage1_61[71]},
      {stage2_63[11],stage2_62[14],stage2_61[24],stage2_60[34],stage2_59[36]}
   );
   gpc606_5 gpc3439 (
      {stage1_59[132], stage1_59[133], stage1_59[134], stage1_59[135], stage1_59[136], stage1_59[137]},
      {stage1_61[72], stage1_61[73], stage1_61[74], stage1_61[75], stage1_61[76], stage1_61[77]},
      {stage2_63[12],stage2_62[15],stage2_61[25],stage2_60[35],stage2_59[37]}
   );
   gpc606_5 gpc3440 (
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22], stage1_60[23]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage2_64[0],stage2_63[13],stage2_62[16],stage2_61[26],stage2_60[36]}
   );
   gpc606_5 gpc3441 (
      {stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27], stage1_60[28], stage1_60[29]},
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage2_64[1],stage2_63[14],stage2_62[17],stage2_61[27],stage2_60[37]}
   );
   gpc606_5 gpc3442 (
      {stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33], stage1_60[34], stage1_60[35]},
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage2_64[2],stage2_63[15],stage2_62[18],stage2_61[28],stage2_60[38]}
   );
   gpc606_5 gpc3443 (
      {stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39], stage1_60[40], stage1_60[41]},
      {stage1_62[18], stage1_62[19], stage1_62[20], stage1_62[21], stage1_62[22], stage1_62[23]},
      {stage2_64[3],stage2_63[16],stage2_62[19],stage2_61[29],stage2_60[39]}
   );
   gpc606_5 gpc3444 (
      {stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45], stage1_60[46], stage1_60[47]},
      {stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29]},
      {stage2_64[4],stage2_63[17],stage2_62[20],stage2_61[30],stage2_60[40]}
   );
   gpc615_5 gpc3445 (
      {stage1_60[48], stage1_60[49], stage1_60[50], stage1_60[51], stage1_60[52]},
      {stage1_61[78]},
      {stage1_62[30], stage1_62[31], stage1_62[32], stage1_62[33], stage1_62[34], stage1_62[35]},
      {stage2_64[5],stage2_63[18],stage2_62[21],stage2_61[31],stage2_60[41]}
   );
   gpc615_5 gpc3446 (
      {stage1_60[53], stage1_60[54], stage1_60[55], stage1_60[56], stage1_60[57]},
      {stage1_61[79]},
      {stage1_62[36], stage1_62[37], stage1_62[38], stage1_62[39], stage1_62[40], stage1_62[41]},
      {stage2_64[6],stage2_63[19],stage2_62[22],stage2_61[32],stage2_60[42]}
   );
   gpc615_5 gpc3447 (
      {stage1_60[58], stage1_60[59], stage1_60[60], stage1_60[61], stage1_60[62]},
      {stage1_61[80]},
      {stage1_62[42], stage1_62[43], stage1_62[44], stage1_62[45], stage1_62[46], stage1_62[47]},
      {stage2_64[7],stage2_63[20],stage2_62[23],stage2_61[33],stage2_60[43]}
   );
   gpc615_5 gpc3448 (
      {stage1_60[63], stage1_60[64], stage1_60[65], stage1_60[66], stage1_60[67]},
      {stage1_61[81]},
      {stage1_62[48], stage1_62[49], stage1_62[50], stage1_62[51], stage1_62[52], stage1_62[53]},
      {stage2_64[8],stage2_63[21],stage2_62[24],stage2_61[34],stage2_60[44]}
   );
   gpc615_5 gpc3449 (
      {stage1_60[68], stage1_60[69], stage1_60[70], stage1_60[71], stage1_60[72]},
      {stage1_61[82]},
      {stage1_62[54], stage1_62[55], stage1_62[56], stage1_62[57], stage1_62[58], stage1_62[59]},
      {stage2_64[9],stage2_63[22],stage2_62[25],stage2_61[35],stage2_60[45]}
   );
   gpc615_5 gpc3450 (
      {stage1_60[73], stage1_60[74], stage1_60[75], stage1_60[76], stage1_60[77]},
      {stage1_61[83]},
      {stage1_62[60], stage1_62[61], stage1_62[62], stage1_62[63], stage1_62[64], stage1_62[65]},
      {stage2_64[10],stage2_63[23],stage2_62[26],stage2_61[36],stage2_60[46]}
   );
   gpc615_5 gpc3451 (
      {stage1_60[78], stage1_60[79], stage1_60[80], stage1_60[81], stage1_60[82]},
      {stage1_61[84]},
      {stage1_62[66], stage1_62[67], stage1_62[68], stage1_62[69], stage1_62[70], stage1_62[71]},
      {stage2_64[11],stage2_63[24],stage2_62[27],stage2_61[37],stage2_60[47]}
   );
   gpc615_5 gpc3452 (
      {stage1_60[83], stage1_60[84], stage1_60[85], stage1_60[86], stage1_60[87]},
      {stage1_61[85]},
      {stage1_62[72], stage1_62[73], stage1_62[74], stage1_62[75], stage1_62[76], stage1_62[77]},
      {stage2_64[12],stage2_63[25],stage2_62[28],stage2_61[38],stage2_60[48]}
   );
   gpc615_5 gpc3453 (
      {stage1_60[88], stage1_60[89], stage1_60[90], stage1_60[91], stage1_60[92]},
      {stage1_61[86]},
      {stage1_62[78], stage1_62[79], stage1_62[80], stage1_62[81], stage1_62[82], stage1_62[83]},
      {stage2_64[13],stage2_63[26],stage2_62[29],stage2_61[39],stage2_60[49]}
   );
   gpc615_5 gpc3454 (
      {stage1_60[93], stage1_60[94], stage1_60[95], stage1_60[96], stage1_60[97]},
      {stage1_61[87]},
      {stage1_62[84], stage1_62[85], stage1_62[86], stage1_62[87], stage1_62[88], stage1_62[89]},
      {stage2_64[14],stage2_63[27],stage2_62[30],stage2_61[40],stage2_60[50]}
   );
   gpc615_5 gpc3455 (
      {stage1_60[98], stage1_60[99], stage1_60[100], stage1_60[101], stage1_60[102]},
      {stage1_61[88]},
      {stage1_62[90], stage1_62[91], stage1_62[92], stage1_62[93], stage1_62[94], stage1_62[95]},
      {stage2_64[15],stage2_63[28],stage2_62[31],stage2_61[41],stage2_60[51]}
   );
   gpc615_5 gpc3456 (
      {stage1_60[103], stage1_60[104], stage1_60[105], stage1_60[106], stage1_60[107]},
      {stage1_61[89]},
      {stage1_62[96], stage1_62[97], stage1_62[98], stage1_62[99], stage1_62[100], stage1_62[101]},
      {stage2_64[16],stage2_63[29],stage2_62[32],stage2_61[42],stage2_60[52]}
   );
   gpc615_5 gpc3457 (
      {stage1_60[108], stage1_60[109], stage1_60[110], stage1_60[111], stage1_60[112]},
      {stage1_61[90]},
      {stage1_62[102], stage1_62[103], stage1_62[104], stage1_62[105], stage1_62[106], stage1_62[107]},
      {stage2_64[17],stage2_63[30],stage2_62[33],stage2_61[43],stage2_60[53]}
   );
   gpc615_5 gpc3458 (
      {stage1_60[113], stage1_60[114], stage1_60[115], stage1_60[116], stage1_60[117]},
      {stage1_61[91]},
      {stage1_62[108], stage1_62[109], stage1_62[110], stage1_62[111], stage1_62[112], stage1_62[113]},
      {stage2_64[18],stage2_63[31],stage2_62[34],stage2_61[44],stage2_60[54]}
   );
   gpc615_5 gpc3459 (
      {stage1_60[118], stage1_60[119], stage1_60[120], stage1_60[121], stage1_60[122]},
      {stage1_61[92]},
      {stage1_62[114], stage1_62[115], stage1_62[116], stage1_62[117], stage1_62[118], stage1_62[119]},
      {stage2_64[19],stage2_63[32],stage2_62[35],stage2_61[45],stage2_60[55]}
   );
   gpc615_5 gpc3460 (
      {stage1_60[123], stage1_60[124], stage1_60[125], stage1_60[126], stage1_60[127]},
      {stage1_61[93]},
      {stage1_62[120], stage1_62[121], stage1_62[122], stage1_62[123], stage1_62[124], stage1_62[125]},
      {stage2_64[20],stage2_63[33],stage2_62[36],stage2_61[46],stage2_60[56]}
   );
   gpc615_5 gpc3461 (
      {stage1_60[128], stage1_60[129], stage1_60[130], stage1_60[131], stage1_60[132]},
      {stage1_61[94]},
      {stage1_62[126], stage1_62[127], stage1_62[128], stage1_62[129], stage1_62[130], stage1_62[131]},
      {stage2_64[21],stage2_63[34],stage2_62[37],stage2_61[47],stage2_60[57]}
   );
   gpc615_5 gpc3462 (
      {stage1_60[133], stage1_60[134], stage1_60[135], stage1_60[136], stage1_60[137]},
      {stage1_61[95]},
      {stage1_62[132], stage1_62[133], stage1_62[134], stage1_62[135], stage1_62[136], stage1_62[137]},
      {stage2_64[22],stage2_63[35],stage2_62[38],stage2_61[48],stage2_60[58]}
   );
   gpc606_5 gpc3463 (
      {stage1_61[96], stage1_61[97], stage1_61[98], stage1_61[99], stage1_61[100], stage1_61[101]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[23],stage2_63[36],stage2_62[39],stage2_61[49]}
   );
   gpc606_5 gpc3464 (
      {stage1_62[138], stage1_62[139], stage1_62[140], stage1_62[141], stage1_62[142], stage1_62[143]},
      {stage1_64[0], stage1_64[1], stage1_64[2], stage1_64[3], stage1_64[4], stage1_64[5]},
      {stage2_66[0],stage2_65[1],stage2_64[24],stage2_63[37],stage2_62[40]}
   );
   gpc606_5 gpc3465 (
      {stage1_62[144], stage1_62[145], stage1_62[146], stage1_62[147], stage1_62[148], stage1_62[149]},
      {stage1_64[6], stage1_64[7], stage1_64[8], stage1_64[9], stage1_64[10], stage1_64[11]},
      {stage2_66[1],stage2_65[2],stage2_64[25],stage2_63[38],stage2_62[41]}
   );
   gpc606_5 gpc3466 (
      {stage1_62[150], stage1_62[151], stage1_62[152], stage1_62[153], stage1_62[154], stage1_62[155]},
      {stage1_64[12], stage1_64[13], stage1_64[14], stage1_64[15], stage1_64[16], stage1_64[17]},
      {stage2_66[2],stage2_65[3],stage2_64[26],stage2_63[39],stage2_62[42]}
   );
   gpc606_5 gpc3467 (
      {stage1_62[156], stage1_62[157], stage1_62[158], stage1_62[159], stage1_62[160], stage1_62[161]},
      {stage1_64[18], stage1_64[19], stage1_64[20], stage1_64[21], stage1_64[22], stage1_64[23]},
      {stage2_66[3],stage2_65[4],stage2_64[27],stage2_63[40],stage2_62[43]}
   );
   gpc606_5 gpc3468 (
      {stage1_62[162], stage1_62[163], stage1_62[164], stage1_62[165], stage1_62[166], stage1_62[167]},
      {stage1_64[24], stage1_64[25], stage1_64[26], stage1_64[27], stage1_64[28], stage1_64[29]},
      {stage2_66[4],stage2_65[5],stage2_64[28],stage2_63[41],stage2_62[44]}
   );
   gpc606_5 gpc3469 (
      {stage1_62[168], stage1_62[169], stage1_62[170], stage1_62[171], stage1_62[172], stage1_62[173]},
      {stage1_64[30], stage1_64[31], stage1_64[32], stage1_64[33], stage1_64[34], stage1_64[35]},
      {stage2_66[5],stage2_65[6],stage2_64[29],stage2_63[42],stage2_62[45]}
   );
   gpc606_5 gpc3470 (
      {stage1_62[174], stage1_62[175], stage1_62[176], stage1_62[177], stage1_62[178], stage1_62[179]},
      {stage1_64[36], stage1_64[37], stage1_64[38], stage1_64[39], stage1_64[40], stage1_64[41]},
      {stage2_66[6],stage2_65[7],stage2_64[30],stage2_63[43],stage2_62[46]}
   );
   gpc606_5 gpc3471 (
      {stage1_62[180], stage1_62[181], stage1_62[182], stage1_62[183], stage1_62[184], stage1_62[185]},
      {stage1_64[42], stage1_64[43], stage1_64[44], stage1_64[45], stage1_64[46], stage1_64[47]},
      {stage2_66[7],stage2_65[8],stage2_64[31],stage2_63[44],stage2_62[47]}
   );
   gpc606_5 gpc3472 (
      {stage1_62[186], stage1_62[187], stage1_62[188], stage1_62[189], stage1_62[190], stage1_62[191]},
      {stage1_64[48], stage1_64[49], stage1_64[50], stage1_64[51], stage1_64[52], stage1_64[53]},
      {stage2_66[8],stage2_65[9],stage2_64[32],stage2_63[45],stage2_62[48]}
   );
   gpc606_5 gpc3473 (
      {stage1_62[192], stage1_62[193], stage1_62[194], stage1_62[195], stage1_62[196], stage1_62[197]},
      {stage1_64[54], stage1_64[55], stage1_64[56], stage1_64[57], stage1_64[58], stage1_64[59]},
      {stage2_66[9],stage2_65[10],stage2_64[33],stage2_63[46],stage2_62[49]}
   );
   gpc606_5 gpc3474 (
      {stage1_63[6], stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11]},
      {stage1_65[0], stage1_65[1], stage1_65[2], stage1_65[3], stage1_65[4], stage1_65[5]},
      {stage2_67[0],stage2_66[10],stage2_65[11],stage2_64[34],stage2_63[47]}
   );
   gpc606_5 gpc3475 (
      {stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17]},
      {stage1_65[6], stage1_65[7], stage1_65[8], stage1_65[9], stage1_65[10], stage1_65[11]},
      {stage2_67[1],stage2_66[11],stage2_65[12],stage2_64[35],stage2_63[48]}
   );
   gpc606_5 gpc3476 (
      {stage1_63[18], stage1_63[19], stage1_63[20], stage1_63[21], stage1_63[22], stage1_63[23]},
      {stage1_65[12], stage1_65[13], stage1_65[14], stage1_65[15], stage1_65[16], stage1_65[17]},
      {stage2_67[2],stage2_66[12],stage2_65[13],stage2_64[36],stage2_63[49]}
   );
   gpc606_5 gpc3477 (
      {stage1_63[24], stage1_63[25], stage1_63[26], stage1_63[27], stage1_63[28], stage1_63[29]},
      {stage1_65[18], stage1_65[19], stage1_65[20], stage1_65[21], stage1_65[22], stage1_65[23]},
      {stage2_67[3],stage2_66[13],stage2_65[14],stage2_64[37],stage2_63[50]}
   );
   gpc606_5 gpc3478 (
      {stage1_63[30], stage1_63[31], stage1_63[32], stage1_63[33], stage1_63[34], stage1_63[35]},
      {stage1_65[24], stage1_65[25], stage1_65[26], stage1_65[27], stage1_65[28], stage1_65[29]},
      {stage2_67[4],stage2_66[14],stage2_65[15],stage2_64[38],stage2_63[51]}
   );
   gpc606_5 gpc3479 (
      {stage1_63[36], stage1_63[37], stage1_63[38], stage1_63[39], stage1_63[40], stage1_63[41]},
      {stage1_65[30], stage1_65[31], stage1_65[32], stage1_65[33], stage1_65[34], stage1_65[35]},
      {stage2_67[5],stage2_66[15],stage2_65[16],stage2_64[39],stage2_63[52]}
   );
   gpc606_5 gpc3480 (
      {stage1_63[42], stage1_63[43], stage1_63[44], stage1_63[45], stage1_63[46], stage1_63[47]},
      {stage1_65[36], stage1_65[37], stage1_65[38], stage1_65[39], stage1_65[40], stage1_65[41]},
      {stage2_67[6],stage2_66[16],stage2_65[17],stage2_64[40],stage2_63[53]}
   );
   gpc1_1 gpc3481 (
      {stage1_0[74]},
      {stage2_0[13]}
   );
   gpc1_1 gpc3482 (
      {stage1_0[75]},
      {stage2_0[14]}
   );
   gpc1_1 gpc3483 (
      {stage1_0[76]},
      {stage2_0[15]}
   );
   gpc1_1 gpc3484 (
      {stage1_0[77]},
      {stage2_0[16]}
   );
   gpc1_1 gpc3485 (
      {stage1_0[78]},
      {stage2_0[17]}
   );
   gpc1_1 gpc3486 (
      {stage1_0[79]},
      {stage2_0[18]}
   );
   gpc1_1 gpc3487 (
      {stage1_0[80]},
      {stage2_0[19]}
   );
   gpc1_1 gpc3488 (
      {stage1_0[81]},
      {stage2_0[20]}
   );
   gpc1_1 gpc3489 (
      {stage1_0[82]},
      {stage2_0[21]}
   );
   gpc1_1 gpc3490 (
      {stage1_0[83]},
      {stage2_0[22]}
   );
   gpc1_1 gpc3491 (
      {stage1_0[84]},
      {stage2_0[23]}
   );
   gpc1_1 gpc3492 (
      {stage1_0[85]},
      {stage2_0[24]}
   );
   gpc1_1 gpc3493 (
      {stage1_0[86]},
      {stage2_0[25]}
   );
   gpc1_1 gpc3494 (
      {stage1_0[87]},
      {stage2_0[26]}
   );
   gpc1_1 gpc3495 (
      {stage1_0[88]},
      {stage2_0[27]}
   );
   gpc1_1 gpc3496 (
      {stage1_0[89]},
      {stage2_0[28]}
   );
   gpc1_1 gpc3497 (
      {stage1_0[90]},
      {stage2_0[29]}
   );
   gpc1_1 gpc3498 (
      {stage1_1[69]},
      {stage2_1[23]}
   );
   gpc1_1 gpc3499 (
      {stage1_1[70]},
      {stage2_1[24]}
   );
   gpc1_1 gpc3500 (
      {stage1_1[71]},
      {stage2_1[25]}
   );
   gpc1_1 gpc3501 (
      {stage1_1[72]},
      {stage2_1[26]}
   );
   gpc1_1 gpc3502 (
      {stage1_1[73]},
      {stage2_1[27]}
   );
   gpc1_1 gpc3503 (
      {stage1_1[74]},
      {stage2_1[28]}
   );
   gpc1_1 gpc3504 (
      {stage1_1[75]},
      {stage2_1[29]}
   );
   gpc1_1 gpc3505 (
      {stage1_1[76]},
      {stage2_1[30]}
   );
   gpc1_1 gpc3506 (
      {stage1_1[77]},
      {stage2_1[31]}
   );
   gpc1_1 gpc3507 (
      {stage1_1[78]},
      {stage2_1[32]}
   );
   gpc1_1 gpc3508 (
      {stage1_1[79]},
      {stage2_1[33]}
   );
   gpc1_1 gpc3509 (
      {stage1_1[80]},
      {stage2_1[34]}
   );
   gpc1_1 gpc3510 (
      {stage1_1[81]},
      {stage2_1[35]}
   );
   gpc1_1 gpc3511 (
      {stage1_1[82]},
      {stage2_1[36]}
   );
   gpc1_1 gpc3512 (
      {stage1_3[92]},
      {stage2_3[39]}
   );
   gpc1_1 gpc3513 (
      {stage1_3[93]},
      {stage2_3[40]}
   );
   gpc1_1 gpc3514 (
      {stage1_3[94]},
      {stage2_3[41]}
   );
   gpc1_1 gpc3515 (
      {stage1_3[95]},
      {stage2_3[42]}
   );
   gpc1_1 gpc3516 (
      {stage1_3[96]},
      {stage2_3[43]}
   );
   gpc1_1 gpc3517 (
      {stage1_3[97]},
      {stage2_3[44]}
   );
   gpc1_1 gpc3518 (
      {stage1_3[98]},
      {stage2_3[45]}
   );
   gpc1_1 gpc3519 (
      {stage1_3[99]},
      {stage2_3[46]}
   );
   gpc1_1 gpc3520 (
      {stage1_3[100]},
      {stage2_3[47]}
   );
   gpc1_1 gpc3521 (
      {stage1_3[101]},
      {stage2_3[48]}
   );
   gpc1_1 gpc3522 (
      {stage1_3[102]},
      {stage2_3[49]}
   );
   gpc1_1 gpc3523 (
      {stage1_3[103]},
      {stage2_3[50]}
   );
   gpc1_1 gpc3524 (
      {stage1_3[104]},
      {stage2_3[51]}
   );
   gpc1_1 gpc3525 (
      {stage1_3[105]},
      {stage2_3[52]}
   );
   gpc1_1 gpc3526 (
      {stage1_3[106]},
      {stage2_3[53]}
   );
   gpc1_1 gpc3527 (
      {stage1_7[106]},
      {stage2_7[39]}
   );
   gpc1_1 gpc3528 (
      {stage1_7[107]},
      {stage2_7[40]}
   );
   gpc1_1 gpc3529 (
      {stage1_7[108]},
      {stage2_7[41]}
   );
   gpc1_1 gpc3530 (
      {stage1_7[109]},
      {stage2_7[42]}
   );
   gpc1_1 gpc3531 (
      {stage1_10[147]},
      {stage2_10[61]}
   );
   gpc1_1 gpc3532 (
      {stage1_10[148]},
      {stage2_10[62]}
   );
   gpc1_1 gpc3533 (
      {stage1_10[149]},
      {stage2_10[63]}
   );
   gpc1_1 gpc3534 (
      {stage1_10[150]},
      {stage2_10[64]}
   );
   gpc1_1 gpc3535 (
      {stage1_10[151]},
      {stage2_10[65]}
   );
   gpc1_1 gpc3536 (
      {stage1_10[152]},
      {stage2_10[66]}
   );
   gpc1_1 gpc3537 (
      {stage1_10[153]},
      {stage2_10[67]}
   );
   gpc1_1 gpc3538 (
      {stage1_10[154]},
      {stage2_10[68]}
   );
   gpc1_1 gpc3539 (
      {stage1_10[155]},
      {stage2_10[69]}
   );
   gpc1_1 gpc3540 (
      {stage1_11[152]},
      {stage2_11[47]}
   );
   gpc1_1 gpc3541 (
      {stage1_11[153]},
      {stage2_11[48]}
   );
   gpc1_1 gpc3542 (
      {stage1_12[132]},
      {stage2_12[53]}
   );
   gpc1_1 gpc3543 (
      {stage1_13[94]},
      {stage2_13[61]}
   );
   gpc1_1 gpc3544 (
      {stage1_13[95]},
      {stage2_13[62]}
   );
   gpc1_1 gpc3545 (
      {stage1_13[96]},
      {stage2_13[63]}
   );
   gpc1_1 gpc3546 (
      {stage1_15[89]},
      {stage2_15[31]}
   );
   gpc1_1 gpc3547 (
      {stage1_15[90]},
      {stage2_15[32]}
   );
   gpc1_1 gpc3548 (
      {stage1_15[91]},
      {stage2_15[33]}
   );
   gpc1_1 gpc3549 (
      {stage1_15[92]},
      {stage2_15[34]}
   );
   gpc1_1 gpc3550 (
      {stage1_15[93]},
      {stage2_15[35]}
   );
   gpc1_1 gpc3551 (
      {stage1_15[94]},
      {stage2_15[36]}
   );
   gpc1_1 gpc3552 (
      {stage1_15[95]},
      {stage2_15[37]}
   );
   gpc1_1 gpc3553 (
      {stage1_15[96]},
      {stage2_15[38]}
   );
   gpc1_1 gpc3554 (
      {stage1_15[97]},
      {stage2_15[39]}
   );
   gpc1_1 gpc3555 (
      {stage1_15[98]},
      {stage2_15[40]}
   );
   gpc1_1 gpc3556 (
      {stage1_15[99]},
      {stage2_15[41]}
   );
   gpc1_1 gpc3557 (
      {stage1_15[100]},
      {stage2_15[42]}
   );
   gpc1_1 gpc3558 (
      {stage1_15[101]},
      {stage2_15[43]}
   );
   gpc1_1 gpc3559 (
      {stage1_15[102]},
      {stage2_15[44]}
   );
   gpc1_1 gpc3560 (
      {stage1_15[103]},
      {stage2_15[45]}
   );
   gpc1_1 gpc3561 (
      {stage1_15[104]},
      {stage2_15[46]}
   );
   gpc1_1 gpc3562 (
      {stage1_15[105]},
      {stage2_15[47]}
   );
   gpc1_1 gpc3563 (
      {stage1_15[106]},
      {stage2_15[48]}
   );
   gpc1_1 gpc3564 (
      {stage1_15[107]},
      {stage2_15[49]}
   );
   gpc1_1 gpc3565 (
      {stage1_15[108]},
      {stage2_15[50]}
   );
   gpc1_1 gpc3566 (
      {stage1_15[109]},
      {stage2_15[51]}
   );
   gpc1_1 gpc3567 (
      {stage1_15[110]},
      {stage2_15[52]}
   );
   gpc1_1 gpc3568 (
      {stage1_15[111]},
      {stage2_15[53]}
   );
   gpc1_1 gpc3569 (
      {stage1_15[112]},
      {stage2_15[54]}
   );
   gpc1_1 gpc3570 (
      {stage1_15[113]},
      {stage2_15[55]}
   );
   gpc1_1 gpc3571 (
      {stage1_15[114]},
      {stage2_15[56]}
   );
   gpc1_1 gpc3572 (
      {stage1_15[115]},
      {stage2_15[57]}
   );
   gpc1_1 gpc3573 (
      {stage1_15[116]},
      {stage2_15[58]}
   );
   gpc1_1 gpc3574 (
      {stage1_15[117]},
      {stage2_15[59]}
   );
   gpc1_1 gpc3575 (
      {stage1_15[118]},
      {stage2_15[60]}
   );
   gpc1_1 gpc3576 (
      {stage1_15[119]},
      {stage2_15[61]}
   );
   gpc1_1 gpc3577 (
      {stage1_15[120]},
      {stage2_15[62]}
   );
   gpc1_1 gpc3578 (
      {stage1_15[121]},
      {stage2_15[63]}
   );
   gpc1_1 gpc3579 (
      {stage1_15[122]},
      {stage2_15[64]}
   );
   gpc1_1 gpc3580 (
      {stage1_15[123]},
      {stage2_15[65]}
   );
   gpc1_1 gpc3581 (
      {stage1_15[124]},
      {stage2_15[66]}
   );
   gpc1_1 gpc3582 (
      {stage1_15[125]},
      {stage2_15[67]}
   );
   gpc1_1 gpc3583 (
      {stage1_15[126]},
      {stage2_15[68]}
   );
   gpc1_1 gpc3584 (
      {stage1_15[127]},
      {stage2_15[69]}
   );
   gpc1_1 gpc3585 (
      {stage1_15[128]},
      {stage2_15[70]}
   );
   gpc1_1 gpc3586 (
      {stage1_15[129]},
      {stage2_15[71]}
   );
   gpc1_1 gpc3587 (
      {stage1_15[130]},
      {stage2_15[72]}
   );
   gpc1_1 gpc3588 (
      {stage1_15[131]},
      {stage2_15[73]}
   );
   gpc1_1 gpc3589 (
      {stage1_16[104]},
      {stage2_16[39]}
   );
   gpc1_1 gpc3590 (
      {stage1_16[105]},
      {stage2_16[40]}
   );
   gpc1_1 gpc3591 (
      {stage1_16[106]},
      {stage2_16[41]}
   );
   gpc1_1 gpc3592 (
      {stage1_16[107]},
      {stage2_16[42]}
   );
   gpc1_1 gpc3593 (
      {stage1_16[108]},
      {stage2_16[43]}
   );
   gpc1_1 gpc3594 (
      {stage1_16[109]},
      {stage2_16[44]}
   );
   gpc1_1 gpc3595 (
      {stage1_16[110]},
      {stage2_16[45]}
   );
   gpc1_1 gpc3596 (
      {stage1_16[111]},
      {stage2_16[46]}
   );
   gpc1_1 gpc3597 (
      {stage1_16[112]},
      {stage2_16[47]}
   );
   gpc1_1 gpc3598 (
      {stage1_16[113]},
      {stage2_16[48]}
   );
   gpc1_1 gpc3599 (
      {stage1_16[114]},
      {stage2_16[49]}
   );
   gpc1_1 gpc3600 (
      {stage1_16[115]},
      {stage2_16[50]}
   );
   gpc1_1 gpc3601 (
      {stage1_16[116]},
      {stage2_16[51]}
   );
   gpc1_1 gpc3602 (
      {stage1_16[117]},
      {stage2_16[52]}
   );
   gpc1_1 gpc3603 (
      {stage1_16[118]},
      {stage2_16[53]}
   );
   gpc1_1 gpc3604 (
      {stage1_16[119]},
      {stage2_16[54]}
   );
   gpc1_1 gpc3605 (
      {stage1_17[102]},
      {stage2_17[48]}
   );
   gpc1_1 gpc3606 (
      {stage1_17[103]},
      {stage2_17[49]}
   );
   gpc1_1 gpc3607 (
      {stage1_17[104]},
      {stage2_17[50]}
   );
   gpc1_1 gpc3608 (
      {stage1_17[105]},
      {stage2_17[51]}
   );
   gpc1_1 gpc3609 (
      {stage1_17[106]},
      {stage2_17[52]}
   );
   gpc1_1 gpc3610 (
      {stage1_17[107]},
      {stage2_17[53]}
   );
   gpc1_1 gpc3611 (
      {stage1_17[108]},
      {stage2_17[54]}
   );
   gpc1_1 gpc3612 (
      {stage1_17[109]},
      {stage2_17[55]}
   );
   gpc1_1 gpc3613 (
      {stage1_17[110]},
      {stage2_17[56]}
   );
   gpc1_1 gpc3614 (
      {stage1_18[71]},
      {stage2_18[37]}
   );
   gpc1_1 gpc3615 (
      {stage1_18[72]},
      {stage2_18[38]}
   );
   gpc1_1 gpc3616 (
      {stage1_18[73]},
      {stage2_18[39]}
   );
   gpc1_1 gpc3617 (
      {stage1_18[74]},
      {stage2_18[40]}
   );
   gpc1_1 gpc3618 (
      {stage1_18[75]},
      {stage2_18[41]}
   );
   gpc1_1 gpc3619 (
      {stage1_18[76]},
      {stage2_18[42]}
   );
   gpc1_1 gpc3620 (
      {stage1_18[77]},
      {stage2_18[43]}
   );
   gpc1_1 gpc3621 (
      {stage1_18[78]},
      {stage2_18[44]}
   );
   gpc1_1 gpc3622 (
      {stage1_18[79]},
      {stage2_18[45]}
   );
   gpc1_1 gpc3623 (
      {stage1_18[80]},
      {stage2_18[46]}
   );
   gpc1_1 gpc3624 (
      {stage1_18[81]},
      {stage2_18[47]}
   );
   gpc1_1 gpc3625 (
      {stage1_18[82]},
      {stage2_18[48]}
   );
   gpc1_1 gpc3626 (
      {stage1_18[83]},
      {stage2_18[49]}
   );
   gpc1_1 gpc3627 (
      {stage1_18[84]},
      {stage2_18[50]}
   );
   gpc1_1 gpc3628 (
      {stage1_18[85]},
      {stage2_18[51]}
   );
   gpc1_1 gpc3629 (
      {stage1_18[86]},
      {stage2_18[52]}
   );
   gpc1_1 gpc3630 (
      {stage1_18[87]},
      {stage2_18[53]}
   );
   gpc1_1 gpc3631 (
      {stage1_18[88]},
      {stage2_18[54]}
   );
   gpc1_1 gpc3632 (
      {stage1_18[89]},
      {stage2_18[55]}
   );
   gpc1_1 gpc3633 (
      {stage1_18[90]},
      {stage2_18[56]}
   );
   gpc1_1 gpc3634 (
      {stage1_18[91]},
      {stage2_18[57]}
   );
   gpc1_1 gpc3635 (
      {stage1_18[92]},
      {stage2_18[58]}
   );
   gpc1_1 gpc3636 (
      {stage1_18[93]},
      {stage2_18[59]}
   );
   gpc1_1 gpc3637 (
      {stage1_18[94]},
      {stage2_18[60]}
   );
   gpc1_1 gpc3638 (
      {stage1_18[95]},
      {stage2_18[61]}
   );
   gpc1_1 gpc3639 (
      {stage1_18[96]},
      {stage2_18[62]}
   );
   gpc1_1 gpc3640 (
      {stage1_18[97]},
      {stage2_18[63]}
   );
   gpc1_1 gpc3641 (
      {stage1_18[98]},
      {stage2_18[64]}
   );
   gpc1_1 gpc3642 (
      {stage1_18[99]},
      {stage2_18[65]}
   );
   gpc1_1 gpc3643 (
      {stage1_19[124]},
      {stage2_19[35]}
   );
   gpc1_1 gpc3644 (
      {stage1_19[125]},
      {stage2_19[36]}
   );
   gpc1_1 gpc3645 (
      {stage1_20[95]},
      {stage2_20[45]}
   );
   gpc1_1 gpc3646 (
      {stage1_20[96]},
      {stage2_20[46]}
   );
   gpc1_1 gpc3647 (
      {stage1_20[97]},
      {stage2_20[47]}
   );
   gpc1_1 gpc3648 (
      {stage1_20[98]},
      {stage2_20[48]}
   );
   gpc1_1 gpc3649 (
      {stage1_20[99]},
      {stage2_20[49]}
   );
   gpc1_1 gpc3650 (
      {stage1_20[100]},
      {stage2_20[50]}
   );
   gpc1_1 gpc3651 (
      {stage1_20[101]},
      {stage2_20[51]}
   );
   gpc1_1 gpc3652 (
      {stage1_20[102]},
      {stage2_20[52]}
   );
   gpc1_1 gpc3653 (
      {stage1_20[103]},
      {stage2_20[53]}
   );
   gpc1_1 gpc3654 (
      {stage1_20[104]},
      {stage2_20[54]}
   );
   gpc1_1 gpc3655 (
      {stage1_20[105]},
      {stage2_20[55]}
   );
   gpc1_1 gpc3656 (
      {stage1_20[106]},
      {stage2_20[56]}
   );
   gpc1_1 gpc3657 (
      {stage1_20[107]},
      {stage2_20[57]}
   );
   gpc1_1 gpc3658 (
      {stage1_20[108]},
      {stage2_20[58]}
   );
   gpc1_1 gpc3659 (
      {stage1_20[109]},
      {stage2_20[59]}
   );
   gpc1_1 gpc3660 (
      {stage1_20[110]},
      {stage2_20[60]}
   );
   gpc1_1 gpc3661 (
      {stage1_20[111]},
      {stage2_20[61]}
   );
   gpc1_1 gpc3662 (
      {stage1_20[112]},
      {stage2_20[62]}
   );
   gpc1_1 gpc3663 (
      {stage1_20[113]},
      {stage2_20[63]}
   );
   gpc1_1 gpc3664 (
      {stage1_20[114]},
      {stage2_20[64]}
   );
   gpc1_1 gpc3665 (
      {stage1_20[115]},
      {stage2_20[65]}
   );
   gpc1_1 gpc3666 (
      {stage1_20[116]},
      {stage2_20[66]}
   );
   gpc1_1 gpc3667 (
      {stage1_20[117]},
      {stage2_20[67]}
   );
   gpc1_1 gpc3668 (
      {stage1_20[118]},
      {stage2_20[68]}
   );
   gpc1_1 gpc3669 (
      {stage1_20[119]},
      {stage2_20[69]}
   );
   gpc1_1 gpc3670 (
      {stage1_20[120]},
      {stage2_20[70]}
   );
   gpc1_1 gpc3671 (
      {stage1_20[121]},
      {stage2_20[71]}
   );
   gpc1_1 gpc3672 (
      {stage1_20[122]},
      {stage2_20[72]}
   );
   gpc1_1 gpc3673 (
      {stage1_20[123]},
      {stage2_20[73]}
   );
   gpc1_1 gpc3674 (
      {stage1_20[124]},
      {stage2_20[74]}
   );
   gpc1_1 gpc3675 (
      {stage1_20[125]},
      {stage2_20[75]}
   );
   gpc1_1 gpc3676 (
      {stage1_20[126]},
      {stage2_20[76]}
   );
   gpc1_1 gpc3677 (
      {stage1_20[127]},
      {stage2_20[77]}
   );
   gpc1_1 gpc3678 (
      {stage1_20[128]},
      {stage2_20[78]}
   );
   gpc1_1 gpc3679 (
      {stage1_20[129]},
      {stage2_20[79]}
   );
   gpc1_1 gpc3680 (
      {stage1_22[87]},
      {stage2_22[36]}
   );
   gpc1_1 gpc3681 (
      {stage1_22[88]},
      {stage2_22[37]}
   );
   gpc1_1 gpc3682 (
      {stage1_22[89]},
      {stage2_22[38]}
   );
   gpc1_1 gpc3683 (
      {stage1_22[90]},
      {stage2_22[39]}
   );
   gpc1_1 gpc3684 (
      {stage1_22[91]},
      {stage2_22[40]}
   );
   gpc1_1 gpc3685 (
      {stage1_23[106]},
      {stage2_23[38]}
   );
   gpc1_1 gpc3686 (
      {stage1_23[107]},
      {stage2_23[39]}
   );
   gpc1_1 gpc3687 (
      {stage1_23[108]},
      {stage2_23[40]}
   );
   gpc1_1 gpc3688 (
      {stage1_23[109]},
      {stage2_23[41]}
   );
   gpc1_1 gpc3689 (
      {stage1_23[110]},
      {stage2_23[42]}
   );
   gpc1_1 gpc3690 (
      {stage1_23[111]},
      {stage2_23[43]}
   );
   gpc1_1 gpc3691 (
      {stage1_23[112]},
      {stage2_23[44]}
   );
   gpc1_1 gpc3692 (
      {stage1_23[113]},
      {stage2_23[45]}
   );
   gpc1_1 gpc3693 (
      {stage1_23[114]},
      {stage2_23[46]}
   );
   gpc1_1 gpc3694 (
      {stage1_23[115]},
      {stage2_23[47]}
   );
   gpc1_1 gpc3695 (
      {stage1_23[116]},
      {stage2_23[48]}
   );
   gpc1_1 gpc3696 (
      {stage1_23[117]},
      {stage2_23[49]}
   );
   gpc1_1 gpc3697 (
      {stage1_23[118]},
      {stage2_23[50]}
   );
   gpc1_1 gpc3698 (
      {stage1_23[119]},
      {stage2_23[51]}
   );
   gpc1_1 gpc3699 (
      {stage1_23[120]},
      {stage2_23[52]}
   );
   gpc1_1 gpc3700 (
      {stage1_23[121]},
      {stage2_23[53]}
   );
   gpc1_1 gpc3701 (
      {stage1_23[122]},
      {stage2_23[54]}
   );
   gpc1_1 gpc3702 (
      {stage1_23[123]},
      {stage2_23[55]}
   );
   gpc1_1 gpc3703 (
      {stage1_23[124]},
      {stage2_23[56]}
   );
   gpc1_1 gpc3704 (
      {stage1_23[125]},
      {stage2_23[57]}
   );
   gpc1_1 gpc3705 (
      {stage1_23[126]},
      {stage2_23[58]}
   );
   gpc1_1 gpc3706 (
      {stage1_23[127]},
      {stage2_23[59]}
   );
   gpc1_1 gpc3707 (
      {stage1_23[128]},
      {stage2_23[60]}
   );
   gpc1_1 gpc3708 (
      {stage1_24[110]},
      {stage2_24[52]}
   );
   gpc1_1 gpc3709 (
      {stage1_24[111]},
      {stage2_24[53]}
   );
   gpc1_1 gpc3710 (
      {stage1_24[112]},
      {stage2_24[54]}
   );
   gpc1_1 gpc3711 (
      {stage1_24[113]},
      {stage2_24[55]}
   );
   gpc1_1 gpc3712 (
      {stage1_24[114]},
      {stage2_24[56]}
   );
   gpc1_1 gpc3713 (
      {stage1_24[115]},
      {stage2_24[57]}
   );
   gpc1_1 gpc3714 (
      {stage1_24[116]},
      {stage2_24[58]}
   );
   gpc1_1 gpc3715 (
      {stage1_24[117]},
      {stage2_24[59]}
   );
   gpc1_1 gpc3716 (
      {stage1_24[118]},
      {stage2_24[60]}
   );
   gpc1_1 gpc3717 (
      {stage1_24[119]},
      {stage2_24[61]}
   );
   gpc1_1 gpc3718 (
      {stage1_24[120]},
      {stage2_24[62]}
   );
   gpc1_1 gpc3719 (
      {stage1_24[121]},
      {stage2_24[63]}
   );
   gpc1_1 gpc3720 (
      {stage1_24[122]},
      {stage2_24[64]}
   );
   gpc1_1 gpc3721 (
      {stage1_24[123]},
      {stage2_24[65]}
   );
   gpc1_1 gpc3722 (
      {stage1_24[124]},
      {stage2_24[66]}
   );
   gpc1_1 gpc3723 (
      {stage1_24[125]},
      {stage2_24[67]}
   );
   gpc1_1 gpc3724 (
      {stage1_24[126]},
      {stage2_24[68]}
   );
   gpc1_1 gpc3725 (
      {stage1_24[127]},
      {stage2_24[69]}
   );
   gpc1_1 gpc3726 (
      {stage1_24[128]},
      {stage2_24[70]}
   );
   gpc1_1 gpc3727 (
      {stage1_24[129]},
      {stage2_24[71]}
   );
   gpc1_1 gpc3728 (
      {stage1_24[130]},
      {stage2_24[72]}
   );
   gpc1_1 gpc3729 (
      {stage1_24[131]},
      {stage2_24[73]}
   );
   gpc1_1 gpc3730 (
      {stage1_24[132]},
      {stage2_24[74]}
   );
   gpc1_1 gpc3731 (
      {stage1_24[133]},
      {stage2_24[75]}
   );
   gpc1_1 gpc3732 (
      {stage1_24[134]},
      {stage2_24[76]}
   );
   gpc1_1 gpc3733 (
      {stage1_24[135]},
      {stage2_24[77]}
   );
   gpc1_1 gpc3734 (
      {stage1_24[136]},
      {stage2_24[78]}
   );
   gpc1_1 gpc3735 (
      {stage1_24[137]},
      {stage2_24[79]}
   );
   gpc1_1 gpc3736 (
      {stage1_24[138]},
      {stage2_24[80]}
   );
   gpc1_1 gpc3737 (
      {stage1_24[139]},
      {stage2_24[81]}
   );
   gpc1_1 gpc3738 (
      {stage1_25[105]},
      {stage2_25[46]}
   );
   gpc1_1 gpc3739 (
      {stage1_25[106]},
      {stage2_25[47]}
   );
   gpc1_1 gpc3740 (
      {stage1_25[107]},
      {stage2_25[48]}
   );
   gpc1_1 gpc3741 (
      {stage1_25[108]},
      {stage2_25[49]}
   );
   gpc1_1 gpc3742 (
      {stage1_25[109]},
      {stage2_25[50]}
   );
   gpc1_1 gpc3743 (
      {stage1_26[129]},
      {stage2_26[40]}
   );
   gpc1_1 gpc3744 (
      {stage1_26[130]},
      {stage2_26[41]}
   );
   gpc1_1 gpc3745 (
      {stage1_26[131]},
      {stage2_26[42]}
   );
   gpc1_1 gpc3746 (
      {stage1_26[132]},
      {stage2_26[43]}
   );
   gpc1_1 gpc3747 (
      {stage1_26[133]},
      {stage2_26[44]}
   );
   gpc1_1 gpc3748 (
      {stage1_26[134]},
      {stage2_26[45]}
   );
   gpc1_1 gpc3749 (
      {stage1_26[135]},
      {stage2_26[46]}
   );
   gpc1_1 gpc3750 (
      {stage1_26[136]},
      {stage2_26[47]}
   );
   gpc1_1 gpc3751 (
      {stage1_26[137]},
      {stage2_26[48]}
   );
   gpc1_1 gpc3752 (
      {stage1_26[138]},
      {stage2_26[49]}
   );
   gpc1_1 gpc3753 (
      {stage1_26[139]},
      {stage2_26[50]}
   );
   gpc1_1 gpc3754 (
      {stage1_26[140]},
      {stage2_26[51]}
   );
   gpc1_1 gpc3755 (
      {stage1_27[93]},
      {stage2_27[46]}
   );
   gpc1_1 gpc3756 (
      {stage1_27[94]},
      {stage2_27[47]}
   );
   gpc1_1 gpc3757 (
      {stage1_27[95]},
      {stage2_27[48]}
   );
   gpc1_1 gpc3758 (
      {stage1_27[96]},
      {stage2_27[49]}
   );
   gpc1_1 gpc3759 (
      {stage1_27[97]},
      {stage2_27[50]}
   );
   gpc1_1 gpc3760 (
      {stage1_27[98]},
      {stage2_27[51]}
   );
   gpc1_1 gpc3761 (
      {stage1_27[99]},
      {stage2_27[52]}
   );
   gpc1_1 gpc3762 (
      {stage1_27[100]},
      {stage2_27[53]}
   );
   gpc1_1 gpc3763 (
      {stage1_27[101]},
      {stage2_27[54]}
   );
   gpc1_1 gpc3764 (
      {stage1_27[102]},
      {stage2_27[55]}
   );
   gpc1_1 gpc3765 (
      {stage1_27[103]},
      {stage2_27[56]}
   );
   gpc1_1 gpc3766 (
      {stage1_27[104]},
      {stage2_27[57]}
   );
   gpc1_1 gpc3767 (
      {stage1_27[105]},
      {stage2_27[58]}
   );
   gpc1_1 gpc3768 (
      {stage1_27[106]},
      {stage2_27[59]}
   );
   gpc1_1 gpc3769 (
      {stage1_27[107]},
      {stage2_27[60]}
   );
   gpc1_1 gpc3770 (
      {stage1_27[108]},
      {stage2_27[61]}
   );
   gpc1_1 gpc3771 (
      {stage1_27[109]},
      {stage2_27[62]}
   );
   gpc1_1 gpc3772 (
      {stage1_27[110]},
      {stage2_27[63]}
   );
   gpc1_1 gpc3773 (
      {stage1_27[111]},
      {stage2_27[64]}
   );
   gpc1_1 gpc3774 (
      {stage1_27[112]},
      {stage2_27[65]}
   );
   gpc1_1 gpc3775 (
      {stage1_27[113]},
      {stage2_27[66]}
   );
   gpc1_1 gpc3776 (
      {stage1_27[114]},
      {stage2_27[67]}
   );
   gpc1_1 gpc3777 (
      {stage1_27[115]},
      {stage2_27[68]}
   );
   gpc1_1 gpc3778 (
      {stage1_27[116]},
      {stage2_27[69]}
   );
   gpc1_1 gpc3779 (
      {stage1_27[117]},
      {stage2_27[70]}
   );
   gpc1_1 gpc3780 (
      {stage1_27[118]},
      {stage2_27[71]}
   );
   gpc1_1 gpc3781 (
      {stage1_28[104]},
      {stage2_28[50]}
   );
   gpc1_1 gpc3782 (
      {stage1_28[105]},
      {stage2_28[51]}
   );
   gpc1_1 gpc3783 (
      {stage1_28[106]},
      {stage2_28[52]}
   );
   gpc1_1 gpc3784 (
      {stage1_28[107]},
      {stage2_28[53]}
   );
   gpc1_1 gpc3785 (
      {stage1_28[108]},
      {stage2_28[54]}
   );
   gpc1_1 gpc3786 (
      {stage1_28[109]},
      {stage2_28[55]}
   );
   gpc1_1 gpc3787 (
      {stage1_28[110]},
      {stage2_28[56]}
   );
   gpc1_1 gpc3788 (
      {stage1_28[111]},
      {stage2_28[57]}
   );
   gpc1_1 gpc3789 (
      {stage1_28[112]},
      {stage2_28[58]}
   );
   gpc1_1 gpc3790 (
      {stage1_28[113]},
      {stage2_28[59]}
   );
   gpc1_1 gpc3791 (
      {stage1_28[114]},
      {stage2_28[60]}
   );
   gpc1_1 gpc3792 (
      {stage1_28[115]},
      {stage2_28[61]}
   );
   gpc1_1 gpc3793 (
      {stage1_28[116]},
      {stage2_28[62]}
   );
   gpc1_1 gpc3794 (
      {stage1_28[117]},
      {stage2_28[63]}
   );
   gpc1_1 gpc3795 (
      {stage1_28[118]},
      {stage2_28[64]}
   );
   gpc1_1 gpc3796 (
      {stage1_28[119]},
      {stage2_28[65]}
   );
   gpc1_1 gpc3797 (
      {stage1_28[120]},
      {stage2_28[66]}
   );
   gpc1_1 gpc3798 (
      {stage1_28[121]},
      {stage2_28[67]}
   );
   gpc1_1 gpc3799 (
      {stage1_28[122]},
      {stage2_28[68]}
   );
   gpc1_1 gpc3800 (
      {stage1_28[123]},
      {stage2_28[69]}
   );
   gpc1_1 gpc3801 (
      {stage1_28[124]},
      {stage2_28[70]}
   );
   gpc1_1 gpc3802 (
      {stage1_28[125]},
      {stage2_28[71]}
   );
   gpc1_1 gpc3803 (
      {stage1_28[126]},
      {stage2_28[72]}
   );
   gpc1_1 gpc3804 (
      {stage1_29[104]},
      {stage2_29[40]}
   );
   gpc1_1 gpc3805 (
      {stage1_29[105]},
      {stage2_29[41]}
   );
   gpc1_1 gpc3806 (
      {stage1_29[106]},
      {stage2_29[42]}
   );
   gpc1_1 gpc3807 (
      {stage1_29[107]},
      {stage2_29[43]}
   );
   gpc1_1 gpc3808 (
      {stage1_29[108]},
      {stage2_29[44]}
   );
   gpc1_1 gpc3809 (
      {stage1_29[109]},
      {stage2_29[45]}
   );
   gpc1_1 gpc3810 (
      {stage1_30[68]},
      {stage2_30[36]}
   );
   gpc1_1 gpc3811 (
      {stage1_30[69]},
      {stage2_30[37]}
   );
   gpc1_1 gpc3812 (
      {stage1_30[70]},
      {stage2_30[38]}
   );
   gpc1_1 gpc3813 (
      {stage1_30[71]},
      {stage2_30[39]}
   );
   gpc1_1 gpc3814 (
      {stage1_30[72]},
      {stage2_30[40]}
   );
   gpc1_1 gpc3815 (
      {stage1_30[73]},
      {stage2_30[41]}
   );
   gpc1_1 gpc3816 (
      {stage1_30[74]},
      {stage2_30[42]}
   );
   gpc1_1 gpc3817 (
      {stage1_30[75]},
      {stage2_30[43]}
   );
   gpc1_1 gpc3818 (
      {stage1_30[76]},
      {stage2_30[44]}
   );
   gpc1_1 gpc3819 (
      {stage1_30[77]},
      {stage2_30[45]}
   );
   gpc1_1 gpc3820 (
      {stage1_30[78]},
      {stage2_30[46]}
   );
   gpc1_1 gpc3821 (
      {stage1_30[79]},
      {stage2_30[47]}
   );
   gpc1_1 gpc3822 (
      {stage1_30[80]},
      {stage2_30[48]}
   );
   gpc1_1 gpc3823 (
      {stage1_30[81]},
      {stage2_30[49]}
   );
   gpc1_1 gpc3824 (
      {stage1_30[82]},
      {stage2_30[50]}
   );
   gpc1_1 gpc3825 (
      {stage1_30[83]},
      {stage2_30[51]}
   );
   gpc1_1 gpc3826 (
      {stage1_30[84]},
      {stage2_30[52]}
   );
   gpc1_1 gpc3827 (
      {stage1_30[85]},
      {stage2_30[53]}
   );
   gpc1_1 gpc3828 (
      {stage1_30[86]},
      {stage2_30[54]}
   );
   gpc1_1 gpc3829 (
      {stage1_30[87]},
      {stage2_30[55]}
   );
   gpc1_1 gpc3830 (
      {stage1_30[88]},
      {stage2_30[56]}
   );
   gpc1_1 gpc3831 (
      {stage1_30[89]},
      {stage2_30[57]}
   );
   gpc1_1 gpc3832 (
      {stage1_30[90]},
      {stage2_30[58]}
   );
   gpc1_1 gpc3833 (
      {stage1_31[99]},
      {stage2_31[38]}
   );
   gpc1_1 gpc3834 (
      {stage1_31[100]},
      {stage2_31[39]}
   );
   gpc1_1 gpc3835 (
      {stage1_31[101]},
      {stage2_31[40]}
   );
   gpc1_1 gpc3836 (
      {stage1_31[102]},
      {stage2_31[41]}
   );
   gpc1_1 gpc3837 (
      {stage1_31[103]},
      {stage2_31[42]}
   );
   gpc1_1 gpc3838 (
      {stage1_31[104]},
      {stage2_31[43]}
   );
   gpc1_1 gpc3839 (
      {stage1_31[105]},
      {stage2_31[44]}
   );
   gpc1_1 gpc3840 (
      {stage1_31[106]},
      {stage2_31[45]}
   );
   gpc1_1 gpc3841 (
      {stage1_31[107]},
      {stage2_31[46]}
   );
   gpc1_1 gpc3842 (
      {stage1_31[108]},
      {stage2_31[47]}
   );
   gpc1_1 gpc3843 (
      {stage1_31[109]},
      {stage2_31[48]}
   );
   gpc1_1 gpc3844 (
      {stage1_31[110]},
      {stage2_31[49]}
   );
   gpc1_1 gpc3845 (
      {stage1_31[111]},
      {stage2_31[50]}
   );
   gpc1_1 gpc3846 (
      {stage1_31[112]},
      {stage2_31[51]}
   );
   gpc1_1 gpc3847 (
      {stage1_31[113]},
      {stage2_31[52]}
   );
   gpc1_1 gpc3848 (
      {stage1_31[114]},
      {stage2_31[53]}
   );
   gpc1_1 gpc3849 (
      {stage1_32[112]},
      {stage2_32[44]}
   );
   gpc1_1 gpc3850 (
      {stage1_32[113]},
      {stage2_32[45]}
   );
   gpc1_1 gpc3851 (
      {stage1_32[114]},
      {stage2_32[46]}
   );
   gpc1_1 gpc3852 (
      {stage1_33[102]},
      {stage2_33[43]}
   );
   gpc1_1 gpc3853 (
      {stage1_33[103]},
      {stage2_33[44]}
   );
   gpc1_1 gpc3854 (
      {stage1_33[104]},
      {stage2_33[45]}
   );
   gpc1_1 gpc3855 (
      {stage1_33[105]},
      {stage2_33[46]}
   );
   gpc1_1 gpc3856 (
      {stage1_33[106]},
      {stage2_33[47]}
   );
   gpc1_1 gpc3857 (
      {stage1_33[107]},
      {stage2_33[48]}
   );
   gpc1_1 gpc3858 (
      {stage1_33[108]},
      {stage2_33[49]}
   );
   gpc1_1 gpc3859 (
      {stage1_33[109]},
      {stage2_33[50]}
   );
   gpc1_1 gpc3860 (
      {stage1_33[110]},
      {stage2_33[51]}
   );
   gpc1_1 gpc3861 (
      {stage1_35[106]},
      {stage2_35[46]}
   );
   gpc1_1 gpc3862 (
      {stage1_35[107]},
      {stage2_35[47]}
   );
   gpc1_1 gpc3863 (
      {stage1_35[108]},
      {stage2_35[48]}
   );
   gpc1_1 gpc3864 (
      {stage1_35[109]},
      {stage2_35[49]}
   );
   gpc1_1 gpc3865 (
      {stage1_35[110]},
      {stage2_35[50]}
   );
   gpc1_1 gpc3866 (
      {stage1_35[111]},
      {stage2_35[51]}
   );
   gpc1_1 gpc3867 (
      {stage1_35[112]},
      {stage2_35[52]}
   );
   gpc1_1 gpc3868 (
      {stage1_35[113]},
      {stage2_35[53]}
   );
   gpc1_1 gpc3869 (
      {stage1_35[114]},
      {stage2_35[54]}
   );
   gpc1_1 gpc3870 (
      {stage1_35[115]},
      {stage2_35[55]}
   );
   gpc1_1 gpc3871 (
      {stage1_35[116]},
      {stage2_35[56]}
   );
   gpc1_1 gpc3872 (
      {stage1_35[117]},
      {stage2_35[57]}
   );
   gpc1_1 gpc3873 (
      {stage1_35[118]},
      {stage2_35[58]}
   );
   gpc1_1 gpc3874 (
      {stage1_36[138]},
      {stage2_36[56]}
   );
   gpc1_1 gpc3875 (
      {stage1_36[139]},
      {stage2_36[57]}
   );
   gpc1_1 gpc3876 (
      {stage1_36[140]},
      {stage2_36[58]}
   );
   gpc1_1 gpc3877 (
      {stage1_36[141]},
      {stage2_36[59]}
   );
   gpc1_1 gpc3878 (
      {stage1_36[142]},
      {stage2_36[60]}
   );
   gpc1_1 gpc3879 (
      {stage1_36[143]},
      {stage2_36[61]}
   );
   gpc1_1 gpc3880 (
      {stage1_36[144]},
      {stage2_36[62]}
   );
   gpc1_1 gpc3881 (
      {stage1_37[93]},
      {stage2_37[43]}
   );
   gpc1_1 gpc3882 (
      {stage1_37[94]},
      {stage2_37[44]}
   );
   gpc1_1 gpc3883 (
      {stage1_37[95]},
      {stage2_37[45]}
   );
   gpc1_1 gpc3884 (
      {stage1_37[96]},
      {stage2_37[46]}
   );
   gpc1_1 gpc3885 (
      {stage1_37[97]},
      {stage2_37[47]}
   );
   gpc1_1 gpc3886 (
      {stage1_37[98]},
      {stage2_37[48]}
   );
   gpc1_1 gpc3887 (
      {stage1_37[99]},
      {stage2_37[49]}
   );
   gpc1_1 gpc3888 (
      {stage1_37[100]},
      {stage2_37[50]}
   );
   gpc1_1 gpc3889 (
      {stage1_37[101]},
      {stage2_37[51]}
   );
   gpc1_1 gpc3890 (
      {stage1_37[102]},
      {stage2_37[52]}
   );
   gpc1_1 gpc3891 (
      {stage1_37[103]},
      {stage2_37[53]}
   );
   gpc1_1 gpc3892 (
      {stage1_37[104]},
      {stage2_37[54]}
   );
   gpc1_1 gpc3893 (
      {stage1_38[134]},
      {stage2_38[44]}
   );
   gpc1_1 gpc3894 (
      {stage1_38[135]},
      {stage2_38[45]}
   );
   gpc1_1 gpc3895 (
      {stage1_38[136]},
      {stage2_38[46]}
   );
   gpc1_1 gpc3896 (
      {stage1_39[98]},
      {stage2_39[54]}
   );
   gpc1_1 gpc3897 (
      {stage1_39[99]},
      {stage2_39[55]}
   );
   gpc1_1 gpc3898 (
      {stage1_39[100]},
      {stage2_39[56]}
   );
   gpc1_1 gpc3899 (
      {stage1_39[101]},
      {stage2_39[57]}
   );
   gpc1_1 gpc3900 (
      {stage1_39[102]},
      {stage2_39[58]}
   );
   gpc1_1 gpc3901 (
      {stage1_39[103]},
      {stage2_39[59]}
   );
   gpc1_1 gpc3902 (
      {stage1_39[104]},
      {stage2_39[60]}
   );
   gpc1_1 gpc3903 (
      {stage1_39[105]},
      {stage2_39[61]}
   );
   gpc1_1 gpc3904 (
      {stage1_39[106]},
      {stage2_39[62]}
   );
   gpc1_1 gpc3905 (
      {stage1_39[107]},
      {stage2_39[63]}
   );
   gpc1_1 gpc3906 (
      {stage1_39[108]},
      {stage2_39[64]}
   );
   gpc1_1 gpc3907 (
      {stage1_39[109]},
      {stage2_39[65]}
   );
   gpc1_1 gpc3908 (
      {stage1_39[110]},
      {stage2_39[66]}
   );
   gpc1_1 gpc3909 (
      {stage1_39[111]},
      {stage2_39[67]}
   );
   gpc1_1 gpc3910 (
      {stage1_39[112]},
      {stage2_39[68]}
   );
   gpc1_1 gpc3911 (
      {stage1_39[113]},
      {stage2_39[69]}
   );
   gpc1_1 gpc3912 (
      {stage1_39[114]},
      {stage2_39[70]}
   );
   gpc1_1 gpc3913 (
      {stage1_39[115]},
      {stage2_39[71]}
   );
   gpc1_1 gpc3914 (
      {stage1_39[116]},
      {stage2_39[72]}
   );
   gpc1_1 gpc3915 (
      {stage1_39[117]},
      {stage2_39[73]}
   );
   gpc1_1 gpc3916 (
      {stage1_39[118]},
      {stage2_39[74]}
   );
   gpc1_1 gpc3917 (
      {stage1_39[119]},
      {stage2_39[75]}
   );
   gpc1_1 gpc3918 (
      {stage1_39[120]},
      {stage2_39[76]}
   );
   gpc1_1 gpc3919 (
      {stage1_39[121]},
      {stage2_39[77]}
   );
   gpc1_1 gpc3920 (
      {stage1_39[122]},
      {stage2_39[78]}
   );
   gpc1_1 gpc3921 (
      {stage1_39[123]},
      {stage2_39[79]}
   );
   gpc1_1 gpc3922 (
      {stage1_39[124]},
      {stage2_39[80]}
   );
   gpc1_1 gpc3923 (
      {stage1_40[91]},
      {stage2_40[44]}
   );
   gpc1_1 gpc3924 (
      {stage1_41[102]},
      {stage2_41[34]}
   );
   gpc1_1 gpc3925 (
      {stage1_41[103]},
      {stage2_41[35]}
   );
   gpc1_1 gpc3926 (
      {stage1_41[104]},
      {stage2_41[36]}
   );
   gpc1_1 gpc3927 (
      {stage1_41[105]},
      {stage2_41[37]}
   );
   gpc1_1 gpc3928 (
      {stage1_41[106]},
      {stage2_41[38]}
   );
   gpc1_1 gpc3929 (
      {stage1_41[107]},
      {stage2_41[39]}
   );
   gpc1_1 gpc3930 (
      {stage1_41[108]},
      {stage2_41[40]}
   );
   gpc1_1 gpc3931 (
      {stage1_41[109]},
      {stage2_41[41]}
   );
   gpc1_1 gpc3932 (
      {stage1_41[110]},
      {stage2_41[42]}
   );
   gpc1_1 gpc3933 (
      {stage1_41[111]},
      {stage2_41[43]}
   );
   gpc1_1 gpc3934 (
      {stage1_41[112]},
      {stage2_41[44]}
   );
   gpc1_1 gpc3935 (
      {stage1_41[113]},
      {stage2_41[45]}
   );
   gpc1_1 gpc3936 (
      {stage1_41[114]},
      {stage2_41[46]}
   );
   gpc1_1 gpc3937 (
      {stage1_41[115]},
      {stage2_41[47]}
   );
   gpc1_1 gpc3938 (
      {stage1_41[116]},
      {stage2_41[48]}
   );
   gpc1_1 gpc3939 (
      {stage1_41[117]},
      {stage2_41[49]}
   );
   gpc1_1 gpc3940 (
      {stage1_41[118]},
      {stage2_41[50]}
   );
   gpc1_1 gpc3941 (
      {stage1_41[119]},
      {stage2_41[51]}
   );
   gpc1_1 gpc3942 (
      {stage1_41[120]},
      {stage2_41[52]}
   );
   gpc1_1 gpc3943 (
      {stage1_41[121]},
      {stage2_41[53]}
   );
   gpc1_1 gpc3944 (
      {stage1_41[122]},
      {stage2_41[54]}
   );
   gpc1_1 gpc3945 (
      {stage1_41[123]},
      {stage2_41[55]}
   );
   gpc1_1 gpc3946 (
      {stage1_41[124]},
      {stage2_41[56]}
   );
   gpc1_1 gpc3947 (
      {stage1_41[125]},
      {stage2_41[57]}
   );
   gpc1_1 gpc3948 (
      {stage1_41[126]},
      {stage2_41[58]}
   );
   gpc1_1 gpc3949 (
      {stage1_41[127]},
      {stage2_41[59]}
   );
   gpc1_1 gpc3950 (
      {stage1_41[128]},
      {stage2_41[60]}
   );
   gpc1_1 gpc3951 (
      {stage1_41[129]},
      {stage2_41[61]}
   );
   gpc1_1 gpc3952 (
      {stage1_41[130]},
      {stage2_41[62]}
   );
   gpc1_1 gpc3953 (
      {stage1_41[131]},
      {stage2_41[63]}
   );
   gpc1_1 gpc3954 (
      {stage1_41[132]},
      {stage2_41[64]}
   );
   gpc1_1 gpc3955 (
      {stage1_41[133]},
      {stage2_41[65]}
   );
   gpc1_1 gpc3956 (
      {stage1_41[134]},
      {stage2_41[66]}
   );
   gpc1_1 gpc3957 (
      {stage1_41[135]},
      {stage2_41[67]}
   );
   gpc1_1 gpc3958 (
      {stage1_41[136]},
      {stage2_41[68]}
   );
   gpc1_1 gpc3959 (
      {stage1_41[137]},
      {stage2_41[69]}
   );
   gpc1_1 gpc3960 (
      {stage1_41[138]},
      {stage2_41[70]}
   );
   gpc1_1 gpc3961 (
      {stage1_41[139]},
      {stage2_41[71]}
   );
   gpc1_1 gpc3962 (
      {stage1_41[140]},
      {stage2_41[72]}
   );
   gpc1_1 gpc3963 (
      {stage1_41[141]},
      {stage2_41[73]}
   );
   gpc1_1 gpc3964 (
      {stage1_41[142]},
      {stage2_41[74]}
   );
   gpc1_1 gpc3965 (
      {stage1_42[162]},
      {stage2_42[53]}
   );
   gpc1_1 gpc3966 (
      {stage1_42[163]},
      {stage2_42[54]}
   );
   gpc1_1 gpc3967 (
      {stage1_42[164]},
      {stage2_42[55]}
   );
   gpc1_1 gpc3968 (
      {stage1_42[165]},
      {stage2_42[56]}
   );
   gpc1_1 gpc3969 (
      {stage1_42[166]},
      {stage2_42[57]}
   );
   gpc1_1 gpc3970 (
      {stage1_42[167]},
      {stage2_42[58]}
   );
   gpc1_1 gpc3971 (
      {stage1_42[168]},
      {stage2_42[59]}
   );
   gpc1_1 gpc3972 (
      {stage1_42[169]},
      {stage2_42[60]}
   );
   gpc1_1 gpc3973 (
      {stage1_42[170]},
      {stage2_42[61]}
   );
   gpc1_1 gpc3974 (
      {stage1_42[171]},
      {stage2_42[62]}
   );
   gpc1_1 gpc3975 (
      {stage1_43[70]},
      {stage2_43[53]}
   );
   gpc1_1 gpc3976 (
      {stage1_43[71]},
      {stage2_43[54]}
   );
   gpc1_1 gpc3977 (
      {stage1_43[72]},
      {stage2_43[55]}
   );
   gpc1_1 gpc3978 (
      {stage1_43[73]},
      {stage2_43[56]}
   );
   gpc1_1 gpc3979 (
      {stage1_43[74]},
      {stage2_43[57]}
   );
   gpc1_1 gpc3980 (
      {stage1_43[75]},
      {stage2_43[58]}
   );
   gpc1_1 gpc3981 (
      {stage1_43[76]},
      {stage2_43[59]}
   );
   gpc1_1 gpc3982 (
      {stage1_43[77]},
      {stage2_43[60]}
   );
   gpc1_1 gpc3983 (
      {stage1_43[78]},
      {stage2_43[61]}
   );
   gpc1_1 gpc3984 (
      {stage1_44[134]},
      {stage2_44[40]}
   );
   gpc1_1 gpc3985 (
      {stage1_44[135]},
      {stage2_44[41]}
   );
   gpc1_1 gpc3986 (
      {stage1_44[136]},
      {stage2_44[42]}
   );
   gpc1_1 gpc3987 (
      {stage1_44[137]},
      {stage2_44[43]}
   );
   gpc1_1 gpc3988 (
      {stage1_44[138]},
      {stage2_44[44]}
   );
   gpc1_1 gpc3989 (
      {stage1_44[139]},
      {stage2_44[45]}
   );
   gpc1_1 gpc3990 (
      {stage1_44[140]},
      {stage2_44[46]}
   );
   gpc1_1 gpc3991 (
      {stage1_44[141]},
      {stage2_44[47]}
   );
   gpc1_1 gpc3992 (
      {stage1_44[142]},
      {stage2_44[48]}
   );
   gpc1_1 gpc3993 (
      {stage1_44[143]},
      {stage2_44[49]}
   );
   gpc1_1 gpc3994 (
      {stage1_44[144]},
      {stage2_44[50]}
   );
   gpc1_1 gpc3995 (
      {stage1_44[145]},
      {stage2_44[51]}
   );
   gpc1_1 gpc3996 (
      {stage1_45[126]},
      {stage2_45[46]}
   );
   gpc1_1 gpc3997 (
      {stage1_45[127]},
      {stage2_45[47]}
   );
   gpc1_1 gpc3998 (
      {stage1_45[128]},
      {stage2_45[48]}
   );
   gpc1_1 gpc3999 (
      {stage1_45[129]},
      {stage2_45[49]}
   );
   gpc1_1 gpc4000 (
      {stage1_45[130]},
      {stage2_45[50]}
   );
   gpc1_1 gpc4001 (
      {stage1_45[131]},
      {stage2_45[51]}
   );
   gpc1_1 gpc4002 (
      {stage1_45[132]},
      {stage2_45[52]}
   );
   gpc1_1 gpc4003 (
      {stage1_45[133]},
      {stage2_45[53]}
   );
   gpc1_1 gpc4004 (
      {stage1_45[134]},
      {stage2_45[54]}
   );
   gpc1_1 gpc4005 (
      {stage1_45[135]},
      {stage2_45[55]}
   );
   gpc1_1 gpc4006 (
      {stage1_45[136]},
      {stage2_45[56]}
   );
   gpc1_1 gpc4007 (
      {stage1_45[137]},
      {stage2_45[57]}
   );
   gpc1_1 gpc4008 (
      {stage1_45[138]},
      {stage2_45[58]}
   );
   gpc1_1 gpc4009 (
      {stage1_45[139]},
      {stage2_45[59]}
   );
   gpc1_1 gpc4010 (
      {stage1_45[140]},
      {stage2_45[60]}
   );
   gpc1_1 gpc4011 (
      {stage1_45[141]},
      {stage2_45[61]}
   );
   gpc1_1 gpc4012 (
      {stage1_45[142]},
      {stage2_45[62]}
   );
   gpc1_1 gpc4013 (
      {stage1_45[143]},
      {stage2_45[63]}
   );
   gpc1_1 gpc4014 (
      {stage1_45[144]},
      {stage2_45[64]}
   );
   gpc1_1 gpc4015 (
      {stage1_45[145]},
      {stage2_45[65]}
   );
   gpc1_1 gpc4016 (
      {stage1_45[146]},
      {stage2_45[66]}
   );
   gpc1_1 gpc4017 (
      {stage1_45[147]},
      {stage2_45[67]}
   );
   gpc1_1 gpc4018 (
      {stage1_45[148]},
      {stage2_45[68]}
   );
   gpc1_1 gpc4019 (
      {stage1_45[149]},
      {stage2_45[69]}
   );
   gpc1_1 gpc4020 (
      {stage1_45[150]},
      {stage2_45[70]}
   );
   gpc1_1 gpc4021 (
      {stage1_45[151]},
      {stage2_45[71]}
   );
   gpc1_1 gpc4022 (
      {stage1_45[152]},
      {stage2_45[72]}
   );
   gpc1_1 gpc4023 (
      {stage1_45[153]},
      {stage2_45[73]}
   );
   gpc1_1 gpc4024 (
      {stage1_45[154]},
      {stage2_45[74]}
   );
   gpc1_1 gpc4025 (
      {stage1_45[155]},
      {stage2_45[75]}
   );
   gpc1_1 gpc4026 (
      {stage1_45[156]},
      {stage2_45[76]}
   );
   gpc1_1 gpc4027 (
      {stage1_45[157]},
      {stage2_45[77]}
   );
   gpc1_1 gpc4028 (
      {stage1_45[158]},
      {stage2_45[78]}
   );
   gpc1_1 gpc4029 (
      {stage1_46[96]},
      {stage2_46[58]}
   );
   gpc1_1 gpc4030 (
      {stage1_46[97]},
      {stage2_46[59]}
   );
   gpc1_1 gpc4031 (
      {stage1_46[98]},
      {stage2_46[60]}
   );
   gpc1_1 gpc4032 (
      {stage1_46[99]},
      {stage2_46[61]}
   );
   gpc1_1 gpc4033 (
      {stage1_46[100]},
      {stage2_46[62]}
   );
   gpc1_1 gpc4034 (
      {stage1_47[102]},
      {stage2_47[43]}
   );
   gpc1_1 gpc4035 (
      {stage1_47[103]},
      {stage2_47[44]}
   );
   gpc1_1 gpc4036 (
      {stage1_47[104]},
      {stage2_47[45]}
   );
   gpc1_1 gpc4037 (
      {stage1_47[105]},
      {stage2_47[46]}
   );
   gpc1_1 gpc4038 (
      {stage1_47[106]},
      {stage2_47[47]}
   );
   gpc1_1 gpc4039 (
      {stage1_47[107]},
      {stage2_47[48]}
   );
   gpc1_1 gpc4040 (
      {stage1_47[108]},
      {stage2_47[49]}
   );
   gpc1_1 gpc4041 (
      {stage1_47[109]},
      {stage2_47[50]}
   );
   gpc1_1 gpc4042 (
      {stage1_47[110]},
      {stage2_47[51]}
   );
   gpc1_1 gpc4043 (
      {stage1_47[111]},
      {stage2_47[52]}
   );
   gpc1_1 gpc4044 (
      {stage1_47[112]},
      {stage2_47[53]}
   );
   gpc1_1 gpc4045 (
      {stage1_47[113]},
      {stage2_47[54]}
   );
   gpc1_1 gpc4046 (
      {stage1_47[114]},
      {stage2_47[55]}
   );
   gpc1_1 gpc4047 (
      {stage1_47[115]},
      {stage2_47[56]}
   );
   gpc1_1 gpc4048 (
      {stage1_47[116]},
      {stage2_47[57]}
   );
   gpc1_1 gpc4049 (
      {stage1_47[117]},
      {stage2_47[58]}
   );
   gpc1_1 gpc4050 (
      {stage1_47[118]},
      {stage2_47[59]}
   );
   gpc1_1 gpc4051 (
      {stage1_47[119]},
      {stage2_47[60]}
   );
   gpc1_1 gpc4052 (
      {stage1_47[120]},
      {stage2_47[61]}
   );
   gpc1_1 gpc4053 (
      {stage1_47[121]},
      {stage2_47[62]}
   );
   gpc1_1 gpc4054 (
      {stage1_47[122]},
      {stage2_47[63]}
   );
   gpc1_1 gpc4055 (
      {stage1_47[123]},
      {stage2_47[64]}
   );
   gpc1_1 gpc4056 (
      {stage1_47[124]},
      {stage2_47[65]}
   );
   gpc1_1 gpc4057 (
      {stage1_47[125]},
      {stage2_47[66]}
   );
   gpc1_1 gpc4058 (
      {stage1_47[126]},
      {stage2_47[67]}
   );
   gpc1_1 gpc4059 (
      {stage1_47[127]},
      {stage2_47[68]}
   );
   gpc1_1 gpc4060 (
      {stage1_47[128]},
      {stage2_47[69]}
   );
   gpc1_1 gpc4061 (
      {stage1_47[129]},
      {stage2_47[70]}
   );
   gpc1_1 gpc4062 (
      {stage1_48[100]},
      {stage2_48[34]}
   );
   gpc1_1 gpc4063 (
      {stage1_48[101]},
      {stage2_48[35]}
   );
   gpc1_1 gpc4064 (
      {stage1_48[102]},
      {stage2_48[36]}
   );
   gpc1_1 gpc4065 (
      {stage1_48[103]},
      {stage2_48[37]}
   );
   gpc1_1 gpc4066 (
      {stage1_48[104]},
      {stage2_48[38]}
   );
   gpc1_1 gpc4067 (
      {stage1_48[105]},
      {stage2_48[39]}
   );
   gpc1_1 gpc4068 (
      {stage1_48[106]},
      {stage2_48[40]}
   );
   gpc1_1 gpc4069 (
      {stage1_48[107]},
      {stage2_48[41]}
   );
   gpc1_1 gpc4070 (
      {stage1_49[78]},
      {stage2_49[41]}
   );
   gpc1_1 gpc4071 (
      {stage1_49[79]},
      {stage2_49[42]}
   );
   gpc1_1 gpc4072 (
      {stage1_49[80]},
      {stage2_49[43]}
   );
   gpc1_1 gpc4073 (
      {stage1_49[81]},
      {stage2_49[44]}
   );
   gpc1_1 gpc4074 (
      {stage1_49[82]},
      {stage2_49[45]}
   );
   gpc1_1 gpc4075 (
      {stage1_49[83]},
      {stage2_49[46]}
   );
   gpc1_1 gpc4076 (
      {stage1_49[84]},
      {stage2_49[47]}
   );
   gpc1_1 gpc4077 (
      {stage1_49[85]},
      {stage2_49[48]}
   );
   gpc1_1 gpc4078 (
      {stage1_49[86]},
      {stage2_49[49]}
   );
   gpc1_1 gpc4079 (
      {stage1_49[87]},
      {stage2_49[50]}
   );
   gpc1_1 gpc4080 (
      {stage1_49[88]},
      {stage2_49[51]}
   );
   gpc1_1 gpc4081 (
      {stage1_49[89]},
      {stage2_49[52]}
   );
   gpc1_1 gpc4082 (
      {stage1_49[90]},
      {stage2_49[53]}
   );
   gpc1_1 gpc4083 (
      {stage1_49[91]},
      {stage2_49[54]}
   );
   gpc1_1 gpc4084 (
      {stage1_49[92]},
      {stage2_49[55]}
   );
   gpc1_1 gpc4085 (
      {stage1_49[93]},
      {stage2_49[56]}
   );
   gpc1_1 gpc4086 (
      {stage1_49[94]},
      {stage2_49[57]}
   );
   gpc1_1 gpc4087 (
      {stage1_49[95]},
      {stage2_49[58]}
   );
   gpc1_1 gpc4088 (
      {stage1_49[96]},
      {stage2_49[59]}
   );
   gpc1_1 gpc4089 (
      {stage1_49[97]},
      {stage2_49[60]}
   );
   gpc1_1 gpc4090 (
      {stage1_49[98]},
      {stage2_49[61]}
   );
   gpc1_1 gpc4091 (
      {stage1_49[99]},
      {stage2_49[62]}
   );
   gpc1_1 gpc4092 (
      {stage1_49[100]},
      {stage2_49[63]}
   );
   gpc1_1 gpc4093 (
      {stage1_49[101]},
      {stage2_49[64]}
   );
   gpc1_1 gpc4094 (
      {stage1_49[102]},
      {stage2_49[65]}
   );
   gpc1_1 gpc4095 (
      {stage1_49[103]},
      {stage2_49[66]}
   );
   gpc1_1 gpc4096 (
      {stage1_49[104]},
      {stage2_49[67]}
   );
   gpc1_1 gpc4097 (
      {stage1_49[105]},
      {stage2_49[68]}
   );
   gpc1_1 gpc4098 (
      {stage1_49[106]},
      {stage2_49[69]}
   );
   gpc1_1 gpc4099 (
      {stage1_49[107]},
      {stage2_49[70]}
   );
   gpc1_1 gpc4100 (
      {stage1_49[108]},
      {stage2_49[71]}
   );
   gpc1_1 gpc4101 (
      {stage1_49[109]},
      {stage2_49[72]}
   );
   gpc1_1 gpc4102 (
      {stage1_49[110]},
      {stage2_49[73]}
   );
   gpc1_1 gpc4103 (
      {stage1_49[111]},
      {stage2_49[74]}
   );
   gpc1_1 gpc4104 (
      {stage1_49[112]},
      {stage2_49[75]}
   );
   gpc1_1 gpc4105 (
      {stage1_49[113]},
      {stage2_49[76]}
   );
   gpc1_1 gpc4106 (
      {stage1_49[114]},
      {stage2_49[77]}
   );
   gpc1_1 gpc4107 (
      {stage1_49[115]},
      {stage2_49[78]}
   );
   gpc1_1 gpc4108 (
      {stage1_49[116]},
      {stage2_49[79]}
   );
   gpc1_1 gpc4109 (
      {stage1_49[117]},
      {stage2_49[80]}
   );
   gpc1_1 gpc4110 (
      {stage1_49[118]},
      {stage2_49[81]}
   );
   gpc1_1 gpc4111 (
      {stage1_49[119]},
      {stage2_49[82]}
   );
   gpc1_1 gpc4112 (
      {stage1_49[120]},
      {stage2_49[83]}
   );
   gpc1_1 gpc4113 (
      {stage1_49[121]},
      {stage2_49[84]}
   );
   gpc1_1 gpc4114 (
      {stage1_49[122]},
      {stage2_49[85]}
   );
   gpc1_1 gpc4115 (
      {stage1_49[123]},
      {stage2_49[86]}
   );
   gpc1_1 gpc4116 (
      {stage1_49[124]},
      {stage2_49[87]}
   );
   gpc1_1 gpc4117 (
      {stage1_49[125]},
      {stage2_49[88]}
   );
   gpc1_1 gpc4118 (
      {stage1_49[126]},
      {stage2_49[89]}
   );
   gpc1_1 gpc4119 (
      {stage1_49[127]},
      {stage2_49[90]}
   );
   gpc1_1 gpc4120 (
      {stage1_49[128]},
      {stage2_49[91]}
   );
   gpc1_1 gpc4121 (
      {stage1_49[129]},
      {stage2_49[92]}
   );
   gpc1_1 gpc4122 (
      {stage1_49[130]},
      {stage2_49[93]}
   );
   gpc1_1 gpc4123 (
      {stage1_49[131]},
      {stage2_49[94]}
   );
   gpc1_1 gpc4124 (
      {stage1_49[132]},
      {stage2_49[95]}
   );
   gpc1_1 gpc4125 (
      {stage1_49[133]},
      {stage2_49[96]}
   );
   gpc1_1 gpc4126 (
      {stage1_49[134]},
      {stage2_49[97]}
   );
   gpc1_1 gpc4127 (
      {stage1_49[135]},
      {stage2_49[98]}
   );
   gpc1_1 gpc4128 (
      {stage1_49[136]},
      {stage2_49[99]}
   );
   gpc1_1 gpc4129 (
      {stage1_49[137]},
      {stage2_49[100]}
   );
   gpc1_1 gpc4130 (
      {stage1_49[138]},
      {stage2_49[101]}
   );
   gpc1_1 gpc4131 (
      {stage1_49[139]},
      {stage2_49[102]}
   );
   gpc1_1 gpc4132 (
      {stage1_49[140]},
      {stage2_49[103]}
   );
   gpc1_1 gpc4133 (
      {stage1_49[141]},
      {stage2_49[104]}
   );
   gpc1_1 gpc4134 (
      {stage1_49[142]},
      {stage2_49[105]}
   );
   gpc1_1 gpc4135 (
      {stage1_49[143]},
      {stage2_49[106]}
   );
   gpc1_1 gpc4136 (
      {stage1_49[144]},
      {stage2_49[107]}
   );
   gpc1_1 gpc4137 (
      {stage1_49[145]},
      {stage2_49[108]}
   );
   gpc1_1 gpc4138 (
      {stage1_49[146]},
      {stage2_49[109]}
   );
   gpc1_1 gpc4139 (
      {stage1_49[147]},
      {stage2_49[110]}
   );
   gpc1_1 gpc4140 (
      {stage1_49[148]},
      {stage2_49[111]}
   );
   gpc1_1 gpc4141 (
      {stage1_49[149]},
      {stage2_49[112]}
   );
   gpc1_1 gpc4142 (
      {stage1_49[150]},
      {stage2_49[113]}
   );
   gpc1_1 gpc4143 (
      {stage1_49[151]},
      {stage2_49[114]}
   );
   gpc1_1 gpc4144 (
      {stage1_50[75]},
      {stage2_50[44]}
   );
   gpc1_1 gpc4145 (
      {stage1_50[76]},
      {stage2_50[45]}
   );
   gpc1_1 gpc4146 (
      {stage1_50[77]},
      {stage2_50[46]}
   );
   gpc1_1 gpc4147 (
      {stage1_50[78]},
      {stage2_50[47]}
   );
   gpc1_1 gpc4148 (
      {stage1_50[79]},
      {stage2_50[48]}
   );
   gpc1_1 gpc4149 (
      {stage1_50[80]},
      {stage2_50[49]}
   );
   gpc1_1 gpc4150 (
      {stage1_50[81]},
      {stage2_50[50]}
   );
   gpc1_1 gpc4151 (
      {stage1_50[82]},
      {stage2_50[51]}
   );
   gpc1_1 gpc4152 (
      {stage1_50[83]},
      {stage2_50[52]}
   );
   gpc1_1 gpc4153 (
      {stage1_50[84]},
      {stage2_50[53]}
   );
   gpc1_1 gpc4154 (
      {stage1_50[85]},
      {stage2_50[54]}
   );
   gpc1_1 gpc4155 (
      {stage1_50[86]},
      {stage2_50[55]}
   );
   gpc1_1 gpc4156 (
      {stage1_50[87]},
      {stage2_50[56]}
   );
   gpc1_1 gpc4157 (
      {stage1_50[88]},
      {stage2_50[57]}
   );
   gpc1_1 gpc4158 (
      {stage1_50[89]},
      {stage2_50[58]}
   );
   gpc1_1 gpc4159 (
      {stage1_50[90]},
      {stage2_50[59]}
   );
   gpc1_1 gpc4160 (
      {stage1_50[91]},
      {stage2_50[60]}
   );
   gpc1_1 gpc4161 (
      {stage1_50[92]},
      {stage2_50[61]}
   );
   gpc1_1 gpc4162 (
      {stage1_50[93]},
      {stage2_50[62]}
   );
   gpc1_1 gpc4163 (
      {stage1_50[94]},
      {stage2_50[63]}
   );
   gpc1_1 gpc4164 (
      {stage1_50[95]},
      {stage2_50[64]}
   );
   gpc1_1 gpc4165 (
      {stage1_50[96]},
      {stage2_50[65]}
   );
   gpc1_1 gpc4166 (
      {stage1_50[97]},
      {stage2_50[66]}
   );
   gpc1_1 gpc4167 (
      {stage1_50[98]},
      {stage2_50[67]}
   );
   gpc1_1 gpc4168 (
      {stage1_51[55]},
      {stage2_51[28]}
   );
   gpc1_1 gpc4169 (
      {stage1_51[56]},
      {stage2_51[29]}
   );
   gpc1_1 gpc4170 (
      {stage1_51[57]},
      {stage2_51[30]}
   );
   gpc1_1 gpc4171 (
      {stage1_51[58]},
      {stage2_51[31]}
   );
   gpc1_1 gpc4172 (
      {stage1_51[59]},
      {stage2_51[32]}
   );
   gpc1_1 gpc4173 (
      {stage1_51[60]},
      {stage2_51[33]}
   );
   gpc1_1 gpc4174 (
      {stage1_51[61]},
      {stage2_51[34]}
   );
   gpc1_1 gpc4175 (
      {stage1_51[62]},
      {stage2_51[35]}
   );
   gpc1_1 gpc4176 (
      {stage1_51[63]},
      {stage2_51[36]}
   );
   gpc1_1 gpc4177 (
      {stage1_51[64]},
      {stage2_51[37]}
   );
   gpc1_1 gpc4178 (
      {stage1_51[65]},
      {stage2_51[38]}
   );
   gpc1_1 gpc4179 (
      {stage1_51[66]},
      {stage2_51[39]}
   );
   gpc1_1 gpc4180 (
      {stage1_51[67]},
      {stage2_51[40]}
   );
   gpc1_1 gpc4181 (
      {stage1_51[68]},
      {stage2_51[41]}
   );
   gpc1_1 gpc4182 (
      {stage1_51[69]},
      {stage2_51[42]}
   );
   gpc1_1 gpc4183 (
      {stage1_51[70]},
      {stage2_51[43]}
   );
   gpc1_1 gpc4184 (
      {stage1_51[71]},
      {stage2_51[44]}
   );
   gpc1_1 gpc4185 (
      {stage1_51[72]},
      {stage2_51[45]}
   );
   gpc1_1 gpc4186 (
      {stage1_51[73]},
      {stage2_51[46]}
   );
   gpc1_1 gpc4187 (
      {stage1_51[74]},
      {stage2_51[47]}
   );
   gpc1_1 gpc4188 (
      {stage1_51[75]},
      {stage2_51[48]}
   );
   gpc1_1 gpc4189 (
      {stage1_51[76]},
      {stage2_51[49]}
   );
   gpc1_1 gpc4190 (
      {stage1_51[77]},
      {stage2_51[50]}
   );
   gpc1_1 gpc4191 (
      {stage1_51[78]},
      {stage2_51[51]}
   );
   gpc1_1 gpc4192 (
      {stage1_51[79]},
      {stage2_51[52]}
   );
   gpc1_1 gpc4193 (
      {stage1_51[80]},
      {stage2_51[53]}
   );
   gpc1_1 gpc4194 (
      {stage1_51[81]},
      {stage2_51[54]}
   );
   gpc1_1 gpc4195 (
      {stage1_51[82]},
      {stage2_51[55]}
   );
   gpc1_1 gpc4196 (
      {stage1_51[83]},
      {stage2_51[56]}
   );
   gpc1_1 gpc4197 (
      {stage1_51[84]},
      {stage2_51[57]}
   );
   gpc1_1 gpc4198 (
      {stage1_51[85]},
      {stage2_51[58]}
   );
   gpc1_1 gpc4199 (
      {stage1_51[86]},
      {stage2_51[59]}
   );
   gpc1_1 gpc4200 (
      {stage1_51[87]},
      {stage2_51[60]}
   );
   gpc1_1 gpc4201 (
      {stage1_51[88]},
      {stage2_51[61]}
   );
   gpc1_1 gpc4202 (
      {stage1_51[89]},
      {stage2_51[62]}
   );
   gpc1_1 gpc4203 (
      {stage1_51[90]},
      {stage2_51[63]}
   );
   gpc1_1 gpc4204 (
      {stage1_51[91]},
      {stage2_51[64]}
   );
   gpc1_1 gpc4205 (
      {stage1_51[92]},
      {stage2_51[65]}
   );
   gpc1_1 gpc4206 (
      {stage1_51[93]},
      {stage2_51[66]}
   );
   gpc1_1 gpc4207 (
      {stage1_51[94]},
      {stage2_51[67]}
   );
   gpc1_1 gpc4208 (
      {stage1_51[95]},
      {stage2_51[68]}
   );
   gpc1_1 gpc4209 (
      {stage1_51[96]},
      {stage2_51[69]}
   );
   gpc1_1 gpc4210 (
      {stage1_51[97]},
      {stage2_51[70]}
   );
   gpc1_1 gpc4211 (
      {stage1_51[98]},
      {stage2_51[71]}
   );
   gpc1_1 gpc4212 (
      {stage1_51[99]},
      {stage2_51[72]}
   );
   gpc1_1 gpc4213 (
      {stage1_51[100]},
      {stage2_51[73]}
   );
   gpc1_1 gpc4214 (
      {stage1_51[101]},
      {stage2_51[74]}
   );
   gpc1_1 gpc4215 (
      {stage1_51[102]},
      {stage2_51[75]}
   );
   gpc1_1 gpc4216 (
      {stage1_51[103]},
      {stage2_51[76]}
   );
   gpc1_1 gpc4217 (
      {stage1_51[104]},
      {stage2_51[77]}
   );
   gpc1_1 gpc4218 (
      {stage1_51[105]},
      {stage2_51[78]}
   );
   gpc1_1 gpc4219 (
      {stage1_52[116]},
      {stage2_52[27]}
   );
   gpc1_1 gpc4220 (
      {stage1_52[117]},
      {stage2_52[28]}
   );
   gpc1_1 gpc4221 (
      {stage1_52[118]},
      {stage2_52[29]}
   );
   gpc1_1 gpc4222 (
      {stage1_52[119]},
      {stage2_52[30]}
   );
   gpc1_1 gpc4223 (
      {stage1_52[120]},
      {stage2_52[31]}
   );
   gpc1_1 gpc4224 (
      {stage1_52[121]},
      {stage2_52[32]}
   );
   gpc1_1 gpc4225 (
      {stage1_52[122]},
      {stage2_52[33]}
   );
   gpc1_1 gpc4226 (
      {stage1_52[123]},
      {stage2_52[34]}
   );
   gpc1_1 gpc4227 (
      {stage1_52[124]},
      {stage2_52[35]}
   );
   gpc1_1 gpc4228 (
      {stage1_52[125]},
      {stage2_52[36]}
   );
   gpc1_1 gpc4229 (
      {stage1_52[126]},
      {stage2_52[37]}
   );
   gpc1_1 gpc4230 (
      {stage1_52[127]},
      {stage2_52[38]}
   );
   gpc1_1 gpc4231 (
      {stage1_52[128]},
      {stage2_52[39]}
   );
   gpc1_1 gpc4232 (
      {stage1_52[129]},
      {stage2_52[40]}
   );
   gpc1_1 gpc4233 (
      {stage1_52[130]},
      {stage2_52[41]}
   );
   gpc1_1 gpc4234 (
      {stage1_52[131]},
      {stage2_52[42]}
   );
   gpc1_1 gpc4235 (
      {stage1_52[132]},
      {stage2_52[43]}
   );
   gpc1_1 gpc4236 (
      {stage1_52[133]},
      {stage2_52[44]}
   );
   gpc1_1 gpc4237 (
      {stage1_52[134]},
      {stage2_52[45]}
   );
   gpc1_1 gpc4238 (
      {stage1_52[135]},
      {stage2_52[46]}
   );
   gpc1_1 gpc4239 (
      {stage1_52[136]},
      {stage2_52[47]}
   );
   gpc1_1 gpc4240 (
      {stage1_52[137]},
      {stage2_52[48]}
   );
   gpc1_1 gpc4241 (
      {stage1_52[138]},
      {stage2_52[49]}
   );
   gpc1_1 gpc4242 (
      {stage1_52[139]},
      {stage2_52[50]}
   );
   gpc1_1 gpc4243 (
      {stage1_53[70]},
      {stage2_53[40]}
   );
   gpc1_1 gpc4244 (
      {stage1_53[71]},
      {stage2_53[41]}
   );
   gpc1_1 gpc4245 (
      {stage1_53[72]},
      {stage2_53[42]}
   );
   gpc1_1 gpc4246 (
      {stage1_53[73]},
      {stage2_53[43]}
   );
   gpc1_1 gpc4247 (
      {stage1_53[74]},
      {stage2_53[44]}
   );
   gpc1_1 gpc4248 (
      {stage1_53[75]},
      {stage2_53[45]}
   );
   gpc1_1 gpc4249 (
      {stage1_53[76]},
      {stage2_53[46]}
   );
   gpc1_1 gpc4250 (
      {stage1_53[77]},
      {stage2_53[47]}
   );
   gpc1_1 gpc4251 (
      {stage1_53[78]},
      {stage2_53[48]}
   );
   gpc1_1 gpc4252 (
      {stage1_53[79]},
      {stage2_53[49]}
   );
   gpc1_1 gpc4253 (
      {stage1_53[80]},
      {stage2_53[50]}
   );
   gpc1_1 gpc4254 (
      {stage1_53[81]},
      {stage2_53[51]}
   );
   gpc1_1 gpc4255 (
      {stage1_53[82]},
      {stage2_53[52]}
   );
   gpc1_1 gpc4256 (
      {stage1_53[83]},
      {stage2_53[53]}
   );
   gpc1_1 gpc4257 (
      {stage1_53[84]},
      {stage2_53[54]}
   );
   gpc1_1 gpc4258 (
      {stage1_53[85]},
      {stage2_53[55]}
   );
   gpc1_1 gpc4259 (
      {stage1_53[86]},
      {stage2_53[56]}
   );
   gpc1_1 gpc4260 (
      {stage1_53[87]},
      {stage2_53[57]}
   );
   gpc1_1 gpc4261 (
      {stage1_53[88]},
      {stage2_53[58]}
   );
   gpc1_1 gpc4262 (
      {stage1_53[89]},
      {stage2_53[59]}
   );
   gpc1_1 gpc4263 (
      {stage1_53[90]},
      {stage2_53[60]}
   );
   gpc1_1 gpc4264 (
      {stage1_53[91]},
      {stage2_53[61]}
   );
   gpc1_1 gpc4265 (
      {stage1_53[92]},
      {stage2_53[62]}
   );
   gpc1_1 gpc4266 (
      {stage1_53[93]},
      {stage2_53[63]}
   );
   gpc1_1 gpc4267 (
      {stage1_53[94]},
      {stage2_53[64]}
   );
   gpc1_1 gpc4268 (
      {stage1_53[95]},
      {stage2_53[65]}
   );
   gpc1_1 gpc4269 (
      {stage1_53[96]},
      {stage2_53[66]}
   );
   gpc1_1 gpc4270 (
      {stage1_53[97]},
      {stage2_53[67]}
   );
   gpc1_1 gpc4271 (
      {stage1_53[98]},
      {stage2_53[68]}
   );
   gpc1_1 gpc4272 (
      {stage1_53[99]},
      {stage2_53[69]}
   );
   gpc1_1 gpc4273 (
      {stage1_53[100]},
      {stage2_53[70]}
   );
   gpc1_1 gpc4274 (
      {stage1_53[101]},
      {stage2_53[71]}
   );
   gpc1_1 gpc4275 (
      {stage1_53[102]},
      {stage2_53[72]}
   );
   gpc1_1 gpc4276 (
      {stage1_53[103]},
      {stage2_53[73]}
   );
   gpc1_1 gpc4277 (
      {stage1_53[104]},
      {stage2_53[74]}
   );
   gpc1_1 gpc4278 (
      {stage1_53[105]},
      {stage2_53[75]}
   );
   gpc1_1 gpc4279 (
      {stage1_53[106]},
      {stage2_53[76]}
   );
   gpc1_1 gpc4280 (
      {stage1_53[107]},
      {stage2_53[77]}
   );
   gpc1_1 gpc4281 (
      {stage1_54[133]},
      {stage2_54[48]}
   );
   gpc1_1 gpc4282 (
      {stage1_54[134]},
      {stage2_54[49]}
   );
   gpc1_1 gpc4283 (
      {stage1_54[135]},
      {stage2_54[50]}
   );
   gpc1_1 gpc4284 (
      {stage1_54[136]},
      {stage2_54[51]}
   );
   gpc1_1 gpc4285 (
      {stage1_54[137]},
      {stage2_54[52]}
   );
   gpc1_1 gpc4286 (
      {stage1_54[138]},
      {stage2_54[53]}
   );
   gpc1_1 gpc4287 (
      {stage1_54[139]},
      {stage2_54[54]}
   );
   gpc1_1 gpc4288 (
      {stage1_54[140]},
      {stage2_54[55]}
   );
   gpc1_1 gpc4289 (
      {stage1_54[141]},
      {stage2_54[56]}
   );
   gpc1_1 gpc4290 (
      {stage1_54[142]},
      {stage2_54[57]}
   );
   gpc1_1 gpc4291 (
      {stage1_54[143]},
      {stage2_54[58]}
   );
   gpc1_1 gpc4292 (
      {stage1_54[144]},
      {stage2_54[59]}
   );
   gpc1_1 gpc4293 (
      {stage1_54[145]},
      {stage2_54[60]}
   );
   gpc1_1 gpc4294 (
      {stage1_54[146]},
      {stage2_54[61]}
   );
   gpc1_1 gpc4295 (
      {stage1_54[147]},
      {stage2_54[62]}
   );
   gpc1_1 gpc4296 (
      {stage1_54[148]},
      {stage2_54[63]}
   );
   gpc1_1 gpc4297 (
      {stage1_54[149]},
      {stage2_54[64]}
   );
   gpc1_1 gpc4298 (
      {stage1_54[150]},
      {stage2_54[65]}
   );
   gpc1_1 gpc4299 (
      {stage1_54[151]},
      {stage2_54[66]}
   );
   gpc1_1 gpc4300 (
      {stage1_54[152]},
      {stage2_54[67]}
   );
   gpc1_1 gpc4301 (
      {stage1_54[153]},
      {stage2_54[68]}
   );
   gpc1_1 gpc4302 (
      {stage1_54[154]},
      {stage2_54[69]}
   );
   gpc1_1 gpc4303 (
      {stage1_54[155]},
      {stage2_54[70]}
   );
   gpc1_1 gpc4304 (
      {stage1_54[156]},
      {stage2_54[71]}
   );
   gpc1_1 gpc4305 (
      {stage1_54[157]},
      {stage2_54[72]}
   );
   gpc1_1 gpc4306 (
      {stage1_54[158]},
      {stage2_54[73]}
   );
   gpc1_1 gpc4307 (
      {stage1_54[159]},
      {stage2_54[74]}
   );
   gpc1_1 gpc4308 (
      {stage1_56[150]},
      {stage2_56[45]}
   );
   gpc1_1 gpc4309 (
      {stage1_56[151]},
      {stage2_56[46]}
   );
   gpc1_1 gpc4310 (
      {stage1_56[152]},
      {stage2_56[47]}
   );
   gpc1_1 gpc4311 (
      {stage1_56[153]},
      {stage2_56[48]}
   );
   gpc1_1 gpc4312 (
      {stage1_56[154]},
      {stage2_56[49]}
   );
   gpc1_1 gpc4313 (
      {stage1_56[155]},
      {stage2_56[50]}
   );
   gpc1_1 gpc4314 (
      {stage1_56[156]},
      {stage2_56[51]}
   );
   gpc1_1 gpc4315 (
      {stage1_56[157]},
      {stage2_56[52]}
   );
   gpc1_1 gpc4316 (
      {stage1_56[158]},
      {stage2_56[53]}
   );
   gpc1_1 gpc4317 (
      {stage1_56[159]},
      {stage2_56[54]}
   );
   gpc1_1 gpc4318 (
      {stage1_56[160]},
      {stage2_56[55]}
   );
   gpc1_1 gpc4319 (
      {stage1_56[161]},
      {stage2_56[56]}
   );
   gpc1_1 gpc4320 (
      {stage1_56[162]},
      {stage2_56[57]}
   );
   gpc1_1 gpc4321 (
      {stage1_56[163]},
      {stage2_56[58]}
   );
   gpc1_1 gpc4322 (
      {stage1_56[164]},
      {stage2_56[59]}
   );
   gpc1_1 gpc4323 (
      {stage1_56[165]},
      {stage2_56[60]}
   );
   gpc1_1 gpc4324 (
      {stage1_56[166]},
      {stage2_56[61]}
   );
   gpc1_1 gpc4325 (
      {stage1_56[167]},
      {stage2_56[62]}
   );
   gpc1_1 gpc4326 (
      {stage1_56[168]},
      {stage2_56[63]}
   );
   gpc1_1 gpc4327 (
      {stage1_56[169]},
      {stage2_56[64]}
   );
   gpc1_1 gpc4328 (
      {stage1_56[170]},
      {stage2_56[65]}
   );
   gpc1_1 gpc4329 (
      {stage1_56[171]},
      {stage2_56[66]}
   );
   gpc1_1 gpc4330 (
      {stage1_56[172]},
      {stage2_56[67]}
   );
   gpc1_1 gpc4331 (
      {stage1_56[173]},
      {stage2_56[68]}
   );
   gpc1_1 gpc4332 (
      {stage1_56[174]},
      {stage2_56[69]}
   );
   gpc1_1 gpc4333 (
      {stage1_56[175]},
      {stage2_56[70]}
   );
   gpc1_1 gpc4334 (
      {stage1_56[176]},
      {stage2_56[71]}
   );
   gpc1_1 gpc4335 (
      {stage1_56[177]},
      {stage2_56[72]}
   );
   gpc1_1 gpc4336 (
      {stage1_57[72]},
      {stage2_57[50]}
   );
   gpc1_1 gpc4337 (
      {stage1_57[73]},
      {stage2_57[51]}
   );
   gpc1_1 gpc4338 (
      {stage1_57[74]},
      {stage2_57[52]}
   );
   gpc1_1 gpc4339 (
      {stage1_57[75]},
      {stage2_57[53]}
   );
   gpc1_1 gpc4340 (
      {stage1_57[76]},
      {stage2_57[54]}
   );
   gpc1_1 gpc4341 (
      {stage1_57[77]},
      {stage2_57[55]}
   );
   gpc1_1 gpc4342 (
      {stage1_57[78]},
      {stage2_57[56]}
   );
   gpc1_1 gpc4343 (
      {stage1_57[79]},
      {stage2_57[57]}
   );
   gpc1_1 gpc4344 (
      {stage1_57[80]},
      {stage2_57[58]}
   );
   gpc1_1 gpc4345 (
      {stage1_57[81]},
      {stage2_57[59]}
   );
   gpc1_1 gpc4346 (
      {stage1_57[82]},
      {stage2_57[60]}
   );
   gpc1_1 gpc4347 (
      {stage1_57[83]},
      {stage2_57[61]}
   );
   gpc1_1 gpc4348 (
      {stage1_57[84]},
      {stage2_57[62]}
   );
   gpc1_1 gpc4349 (
      {stage1_57[85]},
      {stage2_57[63]}
   );
   gpc1_1 gpc4350 (
      {stage1_57[86]},
      {stage2_57[64]}
   );
   gpc1_1 gpc4351 (
      {stage1_57[87]},
      {stage2_57[65]}
   );
   gpc1_1 gpc4352 (
      {stage1_57[88]},
      {stage2_57[66]}
   );
   gpc1_1 gpc4353 (
      {stage1_57[89]},
      {stage2_57[67]}
   );
   gpc1_1 gpc4354 (
      {stage1_57[90]},
      {stage2_57[68]}
   );
   gpc1_1 gpc4355 (
      {stage1_57[91]},
      {stage2_57[69]}
   );
   gpc1_1 gpc4356 (
      {stage1_57[92]},
      {stage2_57[70]}
   );
   gpc1_1 gpc4357 (
      {stage1_57[93]},
      {stage2_57[71]}
   );
   gpc1_1 gpc4358 (
      {stage1_57[94]},
      {stage2_57[72]}
   );
   gpc1_1 gpc4359 (
      {stage1_57[95]},
      {stage2_57[73]}
   );
   gpc1_1 gpc4360 (
      {stage1_57[96]},
      {stage2_57[74]}
   );
   gpc1_1 gpc4361 (
      {stage1_57[97]},
      {stage2_57[75]}
   );
   gpc1_1 gpc4362 (
      {stage1_57[98]},
      {stage2_57[76]}
   );
   gpc1_1 gpc4363 (
      {stage1_57[99]},
      {stage2_57[77]}
   );
   gpc1_1 gpc4364 (
      {stage1_57[100]},
      {stage2_57[78]}
   );
   gpc1_1 gpc4365 (
      {stage1_57[101]},
      {stage2_57[79]}
   );
   gpc1_1 gpc4366 (
      {stage1_57[102]},
      {stage2_57[80]}
   );
   gpc1_1 gpc4367 (
      {stage1_57[103]},
      {stage2_57[81]}
   );
   gpc1_1 gpc4368 (
      {stage1_57[104]},
      {stage2_57[82]}
   );
   gpc1_1 gpc4369 (
      {stage1_58[78]},
      {stage2_58[40]}
   );
   gpc1_1 gpc4370 (
      {stage1_58[79]},
      {stage2_58[41]}
   );
   gpc1_1 gpc4371 (
      {stage1_58[80]},
      {stage2_58[42]}
   );
   gpc1_1 gpc4372 (
      {stage1_58[81]},
      {stage2_58[43]}
   );
   gpc1_1 gpc4373 (
      {stage1_58[82]},
      {stage2_58[44]}
   );
   gpc1_1 gpc4374 (
      {stage1_58[83]},
      {stage2_58[45]}
   );
   gpc1_1 gpc4375 (
      {stage1_58[84]},
      {stage2_58[46]}
   );
   gpc1_1 gpc4376 (
      {stage1_58[85]},
      {stage2_58[47]}
   );
   gpc1_1 gpc4377 (
      {stage1_59[138]},
      {stage2_59[38]}
   );
   gpc1_1 gpc4378 (
      {stage1_59[139]},
      {stage2_59[39]}
   );
   gpc1_1 gpc4379 (
      {stage1_59[140]},
      {stage2_59[40]}
   );
   gpc1_1 gpc4380 (
      {stage1_59[141]},
      {stage2_59[41]}
   );
   gpc1_1 gpc4381 (
      {stage1_59[142]},
      {stage2_59[42]}
   );
   gpc1_1 gpc4382 (
      {stage1_59[143]},
      {stage2_59[43]}
   );
   gpc1_1 gpc4383 (
      {stage1_59[144]},
      {stage2_59[44]}
   );
   gpc1_1 gpc4384 (
      {stage1_59[145]},
      {stage2_59[45]}
   );
   gpc1_1 gpc4385 (
      {stage1_59[146]},
      {stage2_59[46]}
   );
   gpc1_1 gpc4386 (
      {stage1_59[147]},
      {stage2_59[47]}
   );
   gpc1_1 gpc4387 (
      {stage1_60[138]},
      {stage2_60[59]}
   );
   gpc1_1 gpc4388 (
      {stage1_60[139]},
      {stage2_60[60]}
   );
   gpc1_1 gpc4389 (
      {stage1_60[140]},
      {stage2_60[61]}
   );
   gpc1_1 gpc4390 (
      {stage1_60[141]},
      {stage2_60[62]}
   );
   gpc1_1 gpc4391 (
      {stage1_61[102]},
      {stage2_61[50]}
   );
   gpc1_1 gpc4392 (
      {stage1_61[103]},
      {stage2_61[51]}
   );
   gpc1_1 gpc4393 (
      {stage1_61[104]},
      {stage2_61[52]}
   );
   gpc1_1 gpc4394 (
      {stage1_61[105]},
      {stage2_61[53]}
   );
   gpc1_1 gpc4395 (
      {stage1_61[106]},
      {stage2_61[54]}
   );
   gpc1_1 gpc4396 (
      {stage1_61[107]},
      {stage2_61[55]}
   );
   gpc1_1 gpc4397 (
      {stage1_61[108]},
      {stage2_61[56]}
   );
   gpc1_1 gpc4398 (
      {stage1_62[198]},
      {stage2_62[50]}
   );
   gpc1_1 gpc4399 (
      {stage1_62[199]},
      {stage2_62[51]}
   );
   gpc1_1 gpc4400 (
      {stage1_62[200]},
      {stage2_62[52]}
   );
   gpc1_1 gpc4401 (
      {stage1_63[48]},
      {stage2_63[54]}
   );
   gpc1_1 gpc4402 (
      {stage1_63[49]},
      {stage2_63[55]}
   );
   gpc1_1 gpc4403 (
      {stage1_63[50]},
      {stage2_63[56]}
   );
   gpc1_1 gpc4404 (
      {stage1_63[51]},
      {stage2_63[57]}
   );
   gpc1_1 gpc4405 (
      {stage1_63[52]},
      {stage2_63[58]}
   );
   gpc1_1 gpc4406 (
      {stage1_63[53]},
      {stage2_63[59]}
   );
   gpc1_1 gpc4407 (
      {stage1_63[54]},
      {stage2_63[60]}
   );
   gpc1_1 gpc4408 (
      {stage1_63[55]},
      {stage2_63[61]}
   );
   gpc1_1 gpc4409 (
      {stage1_63[56]},
      {stage2_63[62]}
   );
   gpc1_1 gpc4410 (
      {stage1_63[57]},
      {stage2_63[63]}
   );
   gpc1_1 gpc4411 (
      {stage1_63[58]},
      {stage2_63[64]}
   );
   gpc1_1 gpc4412 (
      {stage1_63[59]},
      {stage2_63[65]}
   );
   gpc1_1 gpc4413 (
      {stage1_63[60]},
      {stage2_63[66]}
   );
   gpc1_1 gpc4414 (
      {stage1_63[61]},
      {stage2_63[67]}
   );
   gpc1_1 gpc4415 (
      {stage1_63[62]},
      {stage2_63[68]}
   );
   gpc1_1 gpc4416 (
      {stage1_63[63]},
      {stage2_63[69]}
   );
   gpc1_1 gpc4417 (
      {stage1_63[64]},
      {stage2_63[70]}
   );
   gpc1_1 gpc4418 (
      {stage1_63[65]},
      {stage2_63[71]}
   );
   gpc1_1 gpc4419 (
      {stage1_63[66]},
      {stage2_63[72]}
   );
   gpc1_1 gpc4420 (
      {stage1_63[67]},
      {stage2_63[73]}
   );
   gpc1_1 gpc4421 (
      {stage1_63[68]},
      {stage2_63[74]}
   );
   gpc1_1 gpc4422 (
      {stage1_64[60]},
      {stage2_64[41]}
   );
   gpc1_1 gpc4423 (
      {stage1_64[61]},
      {stage2_64[42]}
   );
   gpc1_1 gpc4424 (
      {stage1_64[62]},
      {stage2_64[43]}
   );
   gpc1_1 gpc4425 (
      {stage1_64[63]},
      {stage2_64[44]}
   );
   gpc615_5 gpc4426 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc4427 (
      {stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9]},
      {stage2_1[1]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc4428 (
      {stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_1[2]},
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc4429 (
      {stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19]},
      {stage2_1[3]},
      {stage2_2[18], stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc7_3 gpc4430 (
      {stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10]},
      {stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc606_5 gpc4431 (
      {stage2_1[11], stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[4],stage3_3[5],stage3_2[5],stage3_1[5]}
   );
   gpc606_5 gpc4432 (
      {stage2_1[17], stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[1],stage3_4[5],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc4433 (
      {stage2_1[23], stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28]},
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17]},
      {stage3_5[2],stage3_4[6],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc4434 (
      {stage2_1[29], stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34]},
      {stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage3_5[3],stage3_4[7],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc615_5 gpc4435 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28]},
      {stage2_3[24]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[4],stage3_4[8],stage3_3[9],stage3_2[9]}
   );
   gpc1163_5 gpc4436 (
      {stage2_3[25], stage2_3[26], stage2_3[27]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_5[0]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[1],stage3_5[5],stage3_4[9],stage3_3[10]}
   );
   gpc606_5 gpc4437 (
      {stage2_3[28], stage2_3[29], stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33]},
      {stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6]},
      {stage3_7[1],stage3_6[2],stage3_5[6],stage3_4[10],stage3_3[11]}
   );
   gpc606_5 gpc4438 (
      {stage2_3[34], stage2_3[35], stage2_3[36], stage2_3[37], stage2_3[38], stage2_3[39]},
      {stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12]},
      {stage3_7[2],stage3_6[3],stage3_5[7],stage3_4[11],stage3_3[12]}
   );
   gpc615_5 gpc4439 (
      {stage2_3[40], stage2_3[41], stage2_3[42], stage2_3[43], stage2_3[44]},
      {stage2_4[12]},
      {stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17], stage2_5[18]},
      {stage3_7[3],stage3_6[4],stage3_5[8],stage3_4[12],stage3_3[13]}
   );
   gpc615_5 gpc4440 (
      {stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48], stage2_3[49]},
      {stage2_4[13]},
      {stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23], stage2_5[24]},
      {stage3_7[4],stage3_6[5],stage3_5[9],stage3_4[13],stage3_3[14]}
   );
   gpc606_5 gpc4441 (
      {stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19]},
      {stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6]},
      {stage3_8[0],stage3_7[5],stage3_6[6],stage3_5[10],stage3_4[14]}
   );
   gpc606_5 gpc4442 (
      {stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11], stage2_6[12]},
      {stage3_8[1],stage3_7[6],stage3_6[7],stage3_5[11],stage3_4[15]}
   );
   gpc606_5 gpc4443 (
      {stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30], stage2_4[31]},
      {stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17], stage2_6[18]},
      {stage3_8[2],stage3_7[7],stage3_6[8],stage3_5[12],stage3_4[16]}
   );
   gpc606_5 gpc4444 (
      {stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36], stage2_4[37]},
      {stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23], stage2_6[24]},
      {stage3_8[3],stage3_7[8],stage3_6[9],stage3_5[13],stage3_4[17]}
   );
   gpc615_5 gpc4445 (
      {stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41], stage2_4[42]},
      {stage2_5[25]},
      {stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29], stage2_6[30]},
      {stage3_8[4],stage3_7[9],stage3_6[10],stage3_5[14],stage3_4[18]}
   );
   gpc606_5 gpc4446 (
      {stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35], stage2_6[36]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[0],stage3_8[5],stage3_7[10],stage3_6[11]}
   );
   gpc606_5 gpc4447 (
      {stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41], stage2_6[42]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[1],stage3_8[6],stage3_7[11],stage3_6[12]}
   );
   gpc606_5 gpc4448 (
      {stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47], stage2_6[48]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[2],stage3_8[7],stage3_7[12],stage3_6[13]}
   );
   gpc615_5 gpc4449 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[18]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[3],stage3_9[3],stage3_8[8],stage3_7[13]}
   );
   gpc615_5 gpc4450 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[19]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[4],stage3_9[4],stage3_8[9],stage3_7[14]}
   );
   gpc615_5 gpc4451 (
      {stage2_7[10], stage2_7[11], stage2_7[12], stage2_7[13], stage2_7[14]},
      {stage2_8[20]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[5],stage3_9[5],stage3_8[10],stage3_7[15]}
   );
   gpc615_5 gpc4452 (
      {stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18], stage2_7[19]},
      {stage2_8[21]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[6],stage3_9[6],stage3_8[11],stage3_7[16]}
   );
   gpc615_5 gpc4453 (
      {stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23], stage2_7[24]},
      {stage2_8[22]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[7],stage3_9[7],stage3_8[12],stage3_7[17]}
   );
   gpc615_5 gpc4454 (
      {stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage2_8[23]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[8],stage3_9[8],stage3_8[13],stage3_7[18]}
   );
   gpc615_5 gpc4455 (
      {stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34]},
      {stage2_8[24]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[9],stage3_9[9],stage3_8[14],stage3_7[19]}
   );
   gpc606_5 gpc4456 (
      {stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[7],stage3_10[10],stage3_9[10],stage3_8[15]}
   );
   gpc606_5 gpc4457 (
      {stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35], stage2_8[36]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[8],stage3_10[11],stage3_9[11],stage3_8[16]}
   );
   gpc606_5 gpc4458 (
      {stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41], stage2_8[42]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[9],stage3_10[12],stage3_9[12],stage3_8[17]}
   );
   gpc606_5 gpc4459 (
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[3],stage3_11[10],stage3_10[13],stage3_9[13]}
   );
   gpc606_5 gpc4460 (
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[4],stage3_11[11],stage3_10[14],stage3_9[14]}
   );
   gpc606_5 gpc4461 (
      {stage2_9[54], stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[5],stage3_11[12],stage3_10[15],stage3_9[15]}
   );
   gpc606_5 gpc4462 (
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[3],stage3_12[6],stage3_11[13],stage3_10[16]}
   );
   gpc606_5 gpc4463 (
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[4],stage3_12[7],stage3_11[14],stage3_10[17]}
   );
   gpc606_5 gpc4464 (
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[5],stage3_12[8],stage3_11[15],stage3_10[18]}
   );
   gpc606_5 gpc4465 (
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[3],stage3_13[6],stage3_12[9],stage3_11[16],stage3_10[19]}
   );
   gpc606_5 gpc4466 (
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[4],stage3_13[7],stage3_12[10],stage3_11[17],stage3_10[20]}
   );
   gpc606_5 gpc4467 (
      {stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53]},
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage3_14[5],stage3_13[8],stage3_12[11],stage3_11[18],stage3_10[21]}
   );
   gpc606_5 gpc4468 (
      {stage2_10[54], stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59]},
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage3_14[6],stage3_13[9],stage3_12[12],stage3_11[19],stage3_10[22]}
   );
   gpc615_5 gpc4469 (
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22]},
      {stage2_12[42]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[7],stage3_13[10],stage3_12[13],stage3_11[20]}
   );
   gpc615_5 gpc4470 (
      {stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27]},
      {stage2_12[43]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[8],stage3_13[11],stage3_12[14],stage3_11[21]}
   );
   gpc615_5 gpc4471 (
      {stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32]},
      {stage2_12[44]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[9],stage3_13[12],stage3_12[15],stage3_11[22]}
   );
   gpc615_5 gpc4472 (
      {stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37]},
      {stage2_12[45]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[10],stage3_13[13],stage3_12[16],stage3_11[23]}
   );
   gpc615_5 gpc4473 (
      {stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42]},
      {stage2_12[46]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[11],stage3_13[14],stage3_12[17],stage3_11[24]}
   );
   gpc606_5 gpc4474 (
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[0],stage3_15[5],stage3_14[12],stage3_13[15]}
   );
   gpc606_5 gpc4475 (
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[1],stage3_15[6],stage3_14[13],stage3_13[16]}
   );
   gpc606_5 gpc4476 (
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[2],stage3_15[7],stage3_14[14],stage3_13[17]}
   );
   gpc606_5 gpc4477 (
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[3],stage3_15[8],stage3_14[15],stage3_13[18]}
   );
   gpc606_5 gpc4478 (
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[4],stage3_15[9],stage3_14[16],stage3_13[19]}
   );
   gpc606_5 gpc4479 (
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[5],stage3_16[5],stage3_15[10],stage3_14[17]}
   );
   gpc606_5 gpc4480 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[6],stage3_16[6],stage3_15[11],stage3_14[18]}
   );
   gpc606_5 gpc4481 (
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[7],stage3_16[7],stage3_15[12],stage3_14[19]}
   );
   gpc606_5 gpc4482 (
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[8],stage3_16[8],stage3_15[13],stage3_14[20]}
   );
   gpc606_5 gpc4483 (
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[9],stage3_16[9],stage3_15[14],stage3_14[21]}
   );
   gpc606_5 gpc4484 (
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[10],stage3_16[10],stage3_15[15],stage3_14[22]}
   );
   gpc606_5 gpc4485 (
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[11],stage3_16[11],stage3_15[16],stage3_14[23]}
   );
   gpc615_5 gpc4486 (
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34]},
      {stage2_16[42]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[7],stage3_17[12],stage3_16[12],stage3_15[17]}
   );
   gpc615_5 gpc4487 (
      {stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39]},
      {stage2_16[43]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[8],stage3_17[13],stage3_16[13],stage3_15[18]}
   );
   gpc615_5 gpc4488 (
      {stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44]},
      {stage2_16[44]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[9],stage3_17[14],stage3_16[14],stage3_15[19]}
   );
   gpc615_5 gpc4489 (
      {stage2_15[45], stage2_15[46], stage2_15[47], stage2_15[48], stage2_15[49]},
      {stage2_16[45]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[10],stage3_17[15],stage3_16[15],stage3_15[20]}
   );
   gpc615_5 gpc4490 (
      {stage2_15[50], stage2_15[51], stage2_15[52], stage2_15[53], stage2_15[54]},
      {stage2_16[46]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[11],stage3_17[16],stage3_16[16],stage3_15[21]}
   );
   gpc606_5 gpc4491 (
      {stage2_16[47], stage2_16[48], stage2_16[49], stage2_16[50], stage2_16[51], stage2_16[52]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[5],stage3_18[12],stage3_17[17],stage3_16[17]}
   );
   gpc606_5 gpc4492 (
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[1],stage3_19[6],stage3_18[13],stage3_17[18]}
   );
   gpc606_5 gpc4493 (
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[2],stage3_19[7],stage3_18[14],stage3_17[19]}
   );
   gpc606_5 gpc4494 (
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage3_21[2],stage3_20[3],stage3_19[8],stage3_18[15],stage3_17[20]}
   );
   gpc615_5 gpc4495 (
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10]},
      {stage2_19[18]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[3],stage3_20[4],stage3_19[9],stage3_18[16]}
   );
   gpc615_5 gpc4496 (
      {stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15]},
      {stage2_19[19]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[4],stage3_20[5],stage3_19[10],stage3_18[17]}
   );
   gpc615_5 gpc4497 (
      {stage2_18[16], stage2_18[17], stage2_18[18], stage2_18[19], stage2_18[20]},
      {stage2_19[20]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[5],stage3_20[6],stage3_19[11],stage3_18[18]}
   );
   gpc615_5 gpc4498 (
      {stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24], stage2_18[25]},
      {stage2_19[21]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[6],stage3_20[7],stage3_19[12],stage3_18[19]}
   );
   gpc615_5 gpc4499 (
      {stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29], stage2_18[30]},
      {stage2_19[22]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[7],stage3_20[8],stage3_19[13],stage3_18[20]}
   );
   gpc615_5 gpc4500 (
      {stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34], stage2_18[35]},
      {stage2_19[23]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[8],stage3_20[9],stage3_19[14],stage3_18[21]}
   );
   gpc615_5 gpc4501 (
      {stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39], stage2_18[40]},
      {stage2_19[24]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[9],stage3_20[10],stage3_19[15],stage3_18[22]}
   );
   gpc615_5 gpc4502 (
      {stage2_18[41], stage2_18[42], stage2_18[43], stage2_18[44], stage2_18[45]},
      {stage2_19[25]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[7],stage3_21[10],stage3_20[11],stage3_19[16],stage3_18[23]}
   );
   gpc615_5 gpc4503 (
      {stage2_18[46], stage2_18[47], stage2_18[48], stage2_18[49], stage2_18[50]},
      {stage2_19[26]},
      {stage2_20[48], stage2_20[49], stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53]},
      {stage3_22[8],stage3_21[11],stage3_20[12],stage3_19[17],stage3_18[24]}
   );
   gpc615_5 gpc4504 (
      {stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54], stage2_18[55]},
      {stage2_19[27]},
      {stage2_20[54], stage2_20[55], stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59]},
      {stage3_22[9],stage3_21[12],stage3_20[13],stage3_19[18],stage3_18[25]}
   );
   gpc615_5 gpc4505 (
      {stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59], stage2_18[60]},
      {stage2_19[28]},
      {stage2_20[60], stage2_20[61], stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65]},
      {stage3_22[10],stage3_21[13],stage3_20[14],stage3_19[19],stage3_18[26]}
   );
   gpc615_5 gpc4506 (
      {stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64], stage2_18[65]},
      {stage2_19[29]},
      {stage2_20[66], stage2_20[67], stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71]},
      {stage3_22[11],stage3_21[14],stage3_20[15],stage3_19[20],stage3_18[27]}
   );
   gpc606_5 gpc4507 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[12],stage3_21[15]}
   );
   gpc606_5 gpc4508 (
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[13],stage3_21[16]}
   );
   gpc606_5 gpc4509 (
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16], stage2_21[17]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[14],stage3_21[17]}
   );
   gpc606_5 gpc4510 (
      {stage2_21[18], stage2_21[19], stage2_21[20], stage2_21[21], stage2_21[22], stage2_21[23]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[15],stage3_21[18]}
   );
   gpc615_5 gpc4511 (
      {stage2_21[24], stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28]},
      {stage2_22[0]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[4],stage3_24[4],stage3_23[4],stage3_22[16],stage3_21[19]}
   );
   gpc615_5 gpc4512 (
      {stage2_21[29], stage2_21[30], stage2_21[31], stage2_21[32], stage2_21[33]},
      {stage2_22[1]},
      {stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35]},
      {stage3_25[5],stage3_24[5],stage3_23[5],stage3_22[17],stage3_21[20]}
   );
   gpc615_5 gpc4513 (
      {stage2_21[34], stage2_21[35], stage2_21[36], stage2_21[37], stage2_21[38]},
      {stage2_22[2]},
      {stage2_23[36], stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40], stage2_23[41]},
      {stage3_25[6],stage3_24[6],stage3_23[6],stage3_22[18],stage3_21[21]}
   );
   gpc615_5 gpc4514 (
      {stage2_21[39], stage2_21[40], stage2_21[41], stage2_21[42], stage2_21[43]},
      {stage2_22[3]},
      {stage2_23[42], stage2_23[43], stage2_23[44], stage2_23[45], stage2_23[46], stage2_23[47]},
      {stage3_25[7],stage3_24[7],stage3_23[7],stage3_22[19],stage3_21[22]}
   );
   gpc615_5 gpc4515 (
      {stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47], stage2_21[48]},
      {stage2_22[4]},
      {stage2_23[48], stage2_23[49], stage2_23[50], stage2_23[51], stage2_23[52], stage2_23[53]},
      {stage3_25[8],stage3_24[8],stage3_23[8],stage3_22[20],stage3_21[23]}
   );
   gpc615_5 gpc4516 (
      {stage2_22[5], stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9]},
      {stage2_23[54]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[9],stage3_24[9],stage3_23[9],stage3_22[21]}
   );
   gpc615_5 gpc4517 (
      {stage2_22[10], stage2_22[11], stage2_22[12], stage2_22[13], stage2_22[14]},
      {stage2_23[55]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[10],stage3_24[10],stage3_23[10],stage3_22[22]}
   );
   gpc615_5 gpc4518 (
      {stage2_22[15], stage2_22[16], stage2_22[17], stage2_22[18], stage2_22[19]},
      {stage2_23[56]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[11],stage3_24[11],stage3_23[11],stage3_22[23]}
   );
   gpc615_5 gpc4519 (
      {stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23], stage2_22[24]},
      {stage2_23[57]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[12],stage3_24[12],stage3_23[12],stage3_22[24]}
   );
   gpc615_5 gpc4520 (
      {stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage2_23[58]},
      {stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29]},
      {stage3_26[4],stage3_25[13],stage3_24[13],stage3_23[13],stage3_22[25]}
   );
   gpc615_5 gpc4521 (
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34]},
      {stage2_23[59]},
      {stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34], stage2_24[35]},
      {stage3_26[5],stage3_25[14],stage3_24[14],stage3_23[14],stage3_22[26]}
   );
   gpc615_5 gpc4522 (
      {stage2_22[35], stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39]},
      {stage2_23[60]},
      {stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40], stage2_24[41]},
      {stage3_26[6],stage3_25[15],stage3_24[15],stage3_23[15],stage3_22[27]}
   );
   gpc606_5 gpc4523 (
      {stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46], stage2_24[47]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[0],stage3_26[7],stage3_25[16],stage3_24[16]}
   );
   gpc606_5 gpc4524 (
      {stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52], stage2_24[53]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[1],stage3_26[8],stage3_25[17],stage3_24[17]}
   );
   gpc606_5 gpc4525 (
      {stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58], stage2_24[59]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[2],stage3_26[9],stage3_25[18],stage3_24[18]}
   );
   gpc606_5 gpc4526 (
      {stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64], stage2_24[65]},
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23]},
      {stage3_28[3],stage3_27[3],stage3_26[10],stage3_25[19],stage3_24[19]}
   );
   gpc606_5 gpc4527 (
      {stage2_24[66], stage2_24[67], stage2_24[68], stage2_24[69], stage2_24[70], stage2_24[71]},
      {stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29]},
      {stage3_28[4],stage3_27[4],stage3_26[11],stage3_25[20],stage3_24[20]}
   );
   gpc2135_5 gpc4528 (
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4]},
      {stage2_26[30], stage2_26[31], stage2_26[32]},
      {stage2_27[0]},
      {stage2_28[0], stage2_28[1]},
      {stage3_29[0],stage3_28[5],stage3_27[5],stage3_26[12],stage3_25[21]}
   );
   gpc606_5 gpc4529 (
      {stage2_25[5], stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10]},
      {stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5], stage2_27[6]},
      {stage3_29[1],stage3_28[6],stage3_27[6],stage3_26[13],stage3_25[22]}
   );
   gpc606_5 gpc4530 (
      {stage2_25[11], stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16]},
      {stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11], stage2_27[12]},
      {stage3_29[2],stage3_28[7],stage3_27[7],stage3_26[14],stage3_25[23]}
   );
   gpc606_5 gpc4531 (
      {stage2_25[17], stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22]},
      {stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17], stage2_27[18]},
      {stage3_29[3],stage3_28[8],stage3_27[8],stage3_26[15],stage3_25[24]}
   );
   gpc606_5 gpc4532 (
      {stage2_25[23], stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28]},
      {stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23], stage2_27[24]},
      {stage3_29[4],stage3_28[9],stage3_27[9],stage3_26[16],stage3_25[25]}
   );
   gpc606_5 gpc4533 (
      {stage2_25[29], stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34]},
      {stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29], stage2_27[30]},
      {stage3_29[5],stage3_28[10],stage3_27[10],stage3_26[17],stage3_25[26]}
   );
   gpc606_5 gpc4534 (
      {stage2_25[35], stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40]},
      {stage2_27[31], stage2_27[32], stage2_27[33], stage2_27[34], stage2_27[35], stage2_27[36]},
      {stage3_29[6],stage3_28[11],stage3_27[11],stage3_26[18],stage3_25[27]}
   );
   gpc615_5 gpc4535 (
      {stage2_25[41], stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45]},
      {stage2_26[33]},
      {stage2_27[37], stage2_27[38], stage2_27[39], stage2_27[40], stage2_27[41], stage2_27[42]},
      {stage3_29[7],stage3_28[12],stage3_27[12],stage3_26[19],stage3_25[28]}
   );
   gpc615_5 gpc4536 (
      {stage2_26[34], stage2_26[35], stage2_26[36], stage2_26[37], stage2_26[38]},
      {stage2_27[43]},
      {stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5], stage2_28[6], stage2_28[7]},
      {stage3_30[0],stage3_29[8],stage3_28[13],stage3_27[13],stage3_26[20]}
   );
   gpc615_5 gpc4537 (
      {stage2_26[39], stage2_26[40], stage2_26[41], stage2_26[42], stage2_26[43]},
      {stage2_27[44]},
      {stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13]},
      {stage3_30[1],stage3_29[9],stage3_28[14],stage3_27[14],stage3_26[21]}
   );
   gpc615_5 gpc4538 (
      {stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47], stage2_26[48]},
      {stage2_27[45]},
      {stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17], stage2_28[18], stage2_28[19]},
      {stage3_30[2],stage3_29[10],stage3_28[15],stage3_27[15],stage3_26[22]}
   );
   gpc615_5 gpc4539 (
      {stage2_26[49], stage2_26[50], stage2_26[51], 1'b0, 1'b0},
      {stage2_27[46]},
      {stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23], stage2_28[24], stage2_28[25]},
      {stage3_30[3],stage3_29[11],stage3_28[16],stage3_27[16],stage3_26[23]}
   );
   gpc615_5 gpc4540 (
      {stage2_27[47], stage2_27[48], stage2_27[49], stage2_27[50], stage2_27[51]},
      {stage2_28[26]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[4],stage3_29[12],stage3_28[17],stage3_27[17]}
   );
   gpc615_5 gpc4541 (
      {stage2_27[52], stage2_27[53], stage2_27[54], stage2_27[55], stage2_27[56]},
      {stage2_28[27]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[5],stage3_29[13],stage3_28[18],stage3_27[18]}
   );
   gpc615_5 gpc4542 (
      {stage2_27[57], stage2_27[58], stage2_27[59], stage2_27[60], stage2_27[61]},
      {stage2_28[28]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[6],stage3_29[14],stage3_28[19],stage3_27[19]}
   );
   gpc615_5 gpc4543 (
      {stage2_27[62], stage2_27[63], stage2_27[64], stage2_27[65], stage2_27[66]},
      {stage2_28[29]},
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage3_31[3],stage3_30[7],stage3_29[15],stage3_28[20],stage3_27[20]}
   );
   gpc615_5 gpc4544 (
      {stage2_27[67], stage2_27[68], stage2_27[69], stage2_27[70], stage2_27[71]},
      {stage2_28[30]},
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage3_31[4],stage3_30[8],stage3_29[16],stage3_28[21],stage3_27[21]}
   );
   gpc606_5 gpc4545 (
      {stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34], stage2_28[35], stage2_28[36]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[5],stage3_30[9],stage3_29[17],stage3_28[22]}
   );
   gpc606_5 gpc4546 (
      {stage2_28[37], stage2_28[38], stage2_28[39], stage2_28[40], stage2_28[41], stage2_28[42]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[6],stage3_30[10],stage3_29[18],stage3_28[23]}
   );
   gpc606_5 gpc4547 (
      {stage2_28[43], stage2_28[44], stage2_28[45], stage2_28[46], stage2_28[47], stage2_28[48]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[7],stage3_30[11],stage3_29[19],stage3_28[24]}
   );
   gpc606_5 gpc4548 (
      {stage2_28[49], stage2_28[50], stage2_28[51], stage2_28[52], stage2_28[53], stage2_28[54]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[8],stage3_30[12],stage3_29[20],stage3_28[25]}
   );
   gpc606_5 gpc4549 (
      {stage2_28[55], stage2_28[56], stage2_28[57], stage2_28[58], stage2_28[59], stage2_28[60]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[9],stage3_30[13],stage3_29[21],stage3_28[26]}
   );
   gpc606_5 gpc4550 (
      {stage2_28[61], stage2_28[62], stage2_28[63], stage2_28[64], stage2_28[65], stage2_28[66]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage3_32[5],stage3_31[10],stage3_30[14],stage3_29[22],stage3_28[27]}
   );
   gpc606_5 gpc4551 (
      {stage2_28[67], stage2_28[68], stage2_28[69], stage2_28[70], stage2_28[71], stage2_28[72]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage3_32[6],stage3_31[11],stage3_30[15],stage3_29[23],stage3_28[28]}
   );
   gpc606_5 gpc4552 (
      {stage2_29[30], stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[7],stage3_31[12],stage3_30[16],stage3_29[24]}
   );
   gpc615_5 gpc4553 (
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46]},
      {stage2_31[6]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[1],stage3_32[8],stage3_31[13],stage3_30[17]}
   );
   gpc615_5 gpc4554 (
      {stage2_30[47], stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51]},
      {stage2_31[7]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[2],stage3_32[9],stage3_31[14],stage3_30[18]}
   );
   gpc606_5 gpc4555 (
      {stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11], stage2_31[12], stage2_31[13]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[2],stage3_33[3],stage3_32[10],stage3_31[15]}
   );
   gpc606_5 gpc4556 (
      {stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17], stage2_31[18], stage2_31[19]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[3],stage3_33[4],stage3_32[11],stage3_31[16]}
   );
   gpc606_5 gpc4557 (
      {stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23], stage2_31[24], stage2_31[25]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[4],stage3_33[5],stage3_32[12],stage3_31[17]}
   );
   gpc606_5 gpc4558 (
      {stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29], stage2_31[30], stage2_31[31]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[5],stage3_33[6],stage3_32[13],stage3_31[18]}
   );
   gpc606_5 gpc4559 (
      {stage2_31[32], stage2_31[33], stage2_31[34], stage2_31[35], stage2_31[36], stage2_31[37]},
      {stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29]},
      {stage3_35[4],stage3_34[6],stage3_33[7],stage3_32[14],stage3_31[19]}
   );
   gpc615_5 gpc4560 (
      {stage2_31[38], stage2_31[39], stage2_31[40], stage2_31[41], stage2_31[42]},
      {stage2_32[12]},
      {stage2_33[30], stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35]},
      {stage3_35[5],stage3_34[7],stage3_33[8],stage3_32[15],stage3_31[20]}
   );
   gpc117_4 gpc4561 (
      {stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17], stage2_32[18], stage2_32[19]},
      {stage2_33[36]},
      {stage2_34[0]},
      {stage3_35[6],stage3_34[8],stage3_33[9],stage3_32[16]}
   );
   gpc117_4 gpc4562 (
      {stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23], stage2_32[24], stage2_32[25], stage2_32[26]},
      {stage2_33[37]},
      {stage2_34[1]},
      {stage3_35[7],stage3_34[9],stage3_33[10],stage3_32[17]}
   );
   gpc606_5 gpc4563 (
      {stage2_32[27], stage2_32[28], stage2_32[29], stage2_32[30], stage2_32[31], stage2_32[32]},
      {stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5], stage2_34[6], stage2_34[7]},
      {stage3_36[0],stage3_35[8],stage3_34[10],stage3_33[11],stage3_32[18]}
   );
   gpc606_5 gpc4564 (
      {stage2_32[33], stage2_32[34], stage2_32[35], stage2_32[36], stage2_32[37], stage2_32[38]},
      {stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11], stage2_34[12], stage2_34[13]},
      {stage3_36[1],stage3_35[9],stage3_34[11],stage3_33[12],stage3_32[19]}
   );
   gpc615_5 gpc4565 (
      {stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17], stage2_34[18]},
      {stage2_35[0]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[0],stage3_36[2],stage3_35[10],stage3_34[12]}
   );
   gpc615_5 gpc4566 (
      {stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23]},
      {stage2_35[1]},
      {stage2_36[6], stage2_36[7], stage2_36[8], stage2_36[9], stage2_36[10], stage2_36[11]},
      {stage3_38[1],stage3_37[1],stage3_36[3],stage3_35[11],stage3_34[13]}
   );
   gpc615_5 gpc4567 (
      {stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5], stage2_35[6]},
      {stage2_36[12]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[2],stage3_37[2],stage3_36[4],stage3_35[12]}
   );
   gpc615_5 gpc4568 (
      {stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage2_36[13]},
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage3_39[1],stage3_38[3],stage3_37[3],stage3_36[5],stage3_35[13]}
   );
   gpc615_5 gpc4569 (
      {stage2_35[12], stage2_35[13], stage2_35[14], stage2_35[15], stage2_35[16]},
      {stage2_36[14]},
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage3_39[2],stage3_38[4],stage3_37[4],stage3_36[6],stage3_35[14]}
   );
   gpc615_5 gpc4570 (
      {stage2_35[17], stage2_35[18], stage2_35[19], stage2_35[20], stage2_35[21]},
      {stage2_36[15]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage3_39[3],stage3_38[5],stage3_37[5],stage3_36[7],stage3_35[15]}
   );
   gpc615_5 gpc4571 (
      {stage2_35[22], stage2_35[23], stage2_35[24], stage2_35[25], stage2_35[26]},
      {stage2_36[16]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage3_39[4],stage3_38[6],stage3_37[6],stage3_36[8],stage3_35[16]}
   );
   gpc615_5 gpc4572 (
      {stage2_35[27], stage2_35[28], stage2_35[29], stage2_35[30], stage2_35[31]},
      {stage2_36[17]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage3_39[5],stage3_38[7],stage3_37[7],stage3_36[9],stage3_35[17]}
   );
   gpc615_5 gpc4573 (
      {stage2_35[32], stage2_35[33], stage2_35[34], stage2_35[35], stage2_35[36]},
      {stage2_36[18]},
      {stage2_37[36], stage2_37[37], stage2_37[38], stage2_37[39], stage2_37[40], stage2_37[41]},
      {stage3_39[6],stage3_38[8],stage3_37[8],stage3_36[10],stage3_35[18]}
   );
   gpc615_5 gpc4574 (
      {stage2_35[37], stage2_35[38], stage2_35[39], stage2_35[40], stage2_35[41]},
      {stage2_36[19]},
      {stage2_37[42], stage2_37[43], stage2_37[44], stage2_37[45], stage2_37[46], stage2_37[47]},
      {stage3_39[7],stage3_38[9],stage3_37[9],stage3_36[11],stage3_35[19]}
   );
   gpc615_5 gpc4575 (
      {stage2_35[42], stage2_35[43], stage2_35[44], stage2_35[45], stage2_35[46]},
      {stage2_36[20]},
      {stage2_37[48], stage2_37[49], stage2_37[50], stage2_37[51], stage2_37[52], stage2_37[53]},
      {stage3_39[8],stage3_38[10],stage3_37[10],stage3_36[12],stage3_35[20]}
   );
   gpc606_5 gpc4576 (
      {stage2_36[21], stage2_36[22], stage2_36[23], stage2_36[24], stage2_36[25], stage2_36[26]},
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage3_40[0],stage3_39[9],stage3_38[11],stage3_37[11],stage3_36[13]}
   );
   gpc606_5 gpc4577 (
      {stage2_36[27], stage2_36[28], stage2_36[29], stage2_36[30], stage2_36[31], stage2_36[32]},
      {stage2_38[6], stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11]},
      {stage3_40[1],stage3_39[10],stage3_38[12],stage3_37[12],stage3_36[14]}
   );
   gpc606_5 gpc4578 (
      {stage2_36[33], stage2_36[34], stage2_36[35], stage2_36[36], stage2_36[37], stage2_36[38]},
      {stage2_38[12], stage2_38[13], stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17]},
      {stage3_40[2],stage3_39[11],stage3_38[13],stage3_37[13],stage3_36[15]}
   );
   gpc606_5 gpc4579 (
      {stage2_36[39], stage2_36[40], stage2_36[41], stage2_36[42], stage2_36[43], stage2_36[44]},
      {stage2_38[18], stage2_38[19], stage2_38[20], stage2_38[21], stage2_38[22], stage2_38[23]},
      {stage3_40[3],stage3_39[12],stage3_38[14],stage3_37[14],stage3_36[16]}
   );
   gpc606_5 gpc4580 (
      {stage2_36[45], stage2_36[46], stage2_36[47], stage2_36[48], stage2_36[49], stage2_36[50]},
      {stage2_38[24], stage2_38[25], stage2_38[26], stage2_38[27], stage2_38[28], stage2_38[29]},
      {stage3_40[4],stage3_39[13],stage3_38[15],stage3_37[15],stage3_36[17]}
   );
   gpc606_5 gpc4581 (
      {stage2_36[51], stage2_36[52], stage2_36[53], stage2_36[54], stage2_36[55], stage2_36[56]},
      {stage2_38[30], stage2_38[31], stage2_38[32], stage2_38[33], stage2_38[34], stage2_38[35]},
      {stage3_40[5],stage3_39[14],stage3_38[16],stage3_37[16],stage3_36[18]}
   );
   gpc606_5 gpc4582 (
      {stage2_36[57], stage2_36[58], stage2_36[59], stage2_36[60], stage2_36[61], stage2_36[62]},
      {stage2_38[36], stage2_38[37], stage2_38[38], stage2_38[39], stage2_38[40], stage2_38[41]},
      {stage3_40[6],stage3_39[15],stage3_38[17],stage3_37[17],stage3_36[19]}
   );
   gpc2135_5 gpc4583 (
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4]},
      {stage2_40[0], stage2_40[1], stage2_40[2]},
      {stage2_41[0]},
      {stage2_42[0], stage2_42[1]},
      {stage3_43[0],stage3_42[0],stage3_41[0],stage3_40[7],stage3_39[16]}
   );
   gpc2135_5 gpc4584 (
      {stage2_39[5], stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9]},
      {stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage2_41[1]},
      {stage2_42[2], stage2_42[3]},
      {stage3_43[1],stage3_42[1],stage3_41[1],stage3_40[8],stage3_39[17]}
   );
   gpc2135_5 gpc4585 (
      {stage2_39[10], stage2_39[11], stage2_39[12], stage2_39[13], stage2_39[14]},
      {stage2_40[6], stage2_40[7], stage2_40[8]},
      {stage2_41[2]},
      {stage2_42[4], stage2_42[5]},
      {stage3_43[2],stage3_42[2],stage3_41[2],stage3_40[9],stage3_39[18]}
   );
   gpc2135_5 gpc4586 (
      {stage2_39[15], stage2_39[16], stage2_39[17], stage2_39[18], stage2_39[19]},
      {stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage2_41[3]},
      {stage2_42[6], stage2_42[7]},
      {stage3_43[3],stage3_42[3],stage3_41[3],stage3_40[10],stage3_39[19]}
   );
   gpc2135_5 gpc4587 (
      {stage2_39[20], stage2_39[21], stage2_39[22], stage2_39[23], stage2_39[24]},
      {stage2_40[12], stage2_40[13], stage2_40[14]},
      {stage2_41[4]},
      {stage2_42[8], stage2_42[9]},
      {stage3_43[4],stage3_42[4],stage3_41[4],stage3_40[11],stage3_39[20]}
   );
   gpc2135_5 gpc4588 (
      {stage2_39[25], stage2_39[26], stage2_39[27], stage2_39[28], stage2_39[29]},
      {stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage2_41[5]},
      {stage2_42[10], stage2_42[11]},
      {stage3_43[5],stage3_42[5],stage3_41[5],stage3_40[12],stage3_39[21]}
   );
   gpc2135_5 gpc4589 (
      {stage2_39[30], stage2_39[31], stage2_39[32], stage2_39[33], stage2_39[34]},
      {stage2_40[18], stage2_40[19], stage2_40[20]},
      {stage2_41[6]},
      {stage2_42[12], stage2_42[13]},
      {stage3_43[6],stage3_42[6],stage3_41[6],stage3_40[13],stage3_39[22]}
   );
   gpc2135_5 gpc4590 (
      {stage2_39[35], stage2_39[36], stage2_39[37], stage2_39[38], stage2_39[39]},
      {stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage2_41[7]},
      {stage2_42[14], stage2_42[15]},
      {stage3_43[7],stage3_42[7],stage3_41[7],stage3_40[14],stage3_39[23]}
   );
   gpc2135_5 gpc4591 (
      {stage2_39[40], stage2_39[41], stage2_39[42], stage2_39[43], stage2_39[44]},
      {stage2_40[24], stage2_40[25], stage2_40[26]},
      {stage2_41[8]},
      {stage2_42[16], stage2_42[17]},
      {stage3_43[8],stage3_42[8],stage3_41[8],stage3_40[15],stage3_39[24]}
   );
   gpc606_5 gpc4592 (
      {stage2_39[45], stage2_39[46], stage2_39[47], stage2_39[48], stage2_39[49], stage2_39[50]},
      {stage2_41[9], stage2_41[10], stage2_41[11], stage2_41[12], stage2_41[13], stage2_41[14]},
      {stage3_43[9],stage3_42[9],stage3_41[9],stage3_40[16],stage3_39[25]}
   );
   gpc606_5 gpc4593 (
      {stage2_39[51], stage2_39[52], stage2_39[53], stage2_39[54], stage2_39[55], stage2_39[56]},
      {stage2_41[15], stage2_41[16], stage2_41[17], stage2_41[18], stage2_41[19], stage2_41[20]},
      {stage3_43[10],stage3_42[10],stage3_41[10],stage3_40[17],stage3_39[26]}
   );
   gpc606_5 gpc4594 (
      {stage2_39[57], stage2_39[58], stage2_39[59], stage2_39[60], stage2_39[61], stage2_39[62]},
      {stage2_41[21], stage2_41[22], stage2_41[23], stage2_41[24], stage2_41[25], stage2_41[26]},
      {stage3_43[11],stage3_42[11],stage3_41[11],stage3_40[18],stage3_39[27]}
   );
   gpc606_5 gpc4595 (
      {stage2_39[63], stage2_39[64], stage2_39[65], stage2_39[66], stage2_39[67], stage2_39[68]},
      {stage2_41[27], stage2_41[28], stage2_41[29], stage2_41[30], stage2_41[31], stage2_41[32]},
      {stage3_43[12],stage3_42[12],stage3_41[12],stage3_40[19],stage3_39[28]}
   );
   gpc606_5 gpc4596 (
      {stage2_39[69], stage2_39[70], stage2_39[71], stage2_39[72], stage2_39[73], stage2_39[74]},
      {stage2_41[33], stage2_41[34], stage2_41[35], stage2_41[36], stage2_41[37], stage2_41[38]},
      {stage3_43[13],stage3_42[13],stage3_41[13],stage3_40[20],stage3_39[29]}
   );
   gpc606_5 gpc4597 (
      {stage2_39[75], stage2_39[76], stage2_39[77], stage2_39[78], stage2_39[79], stage2_39[80]},
      {stage2_41[39], stage2_41[40], stage2_41[41], stage2_41[42], stage2_41[43], stage2_41[44]},
      {stage3_43[14],stage3_42[14],stage3_41[14],stage3_40[21],stage3_39[30]}
   );
   gpc606_5 gpc4598 (
      {stage2_40[27], stage2_40[28], stage2_40[29], stage2_40[30], stage2_40[31], stage2_40[32]},
      {stage2_42[18], stage2_42[19], stage2_42[20], stage2_42[21], stage2_42[22], stage2_42[23]},
      {stage3_44[0],stage3_43[15],stage3_42[15],stage3_41[15],stage3_40[22]}
   );
   gpc606_5 gpc4599 (
      {stage2_40[33], stage2_40[34], stage2_40[35], stage2_40[36], stage2_40[37], stage2_40[38]},
      {stage2_42[24], stage2_42[25], stage2_42[26], stage2_42[27], stage2_42[28], stage2_42[29]},
      {stage3_44[1],stage3_43[16],stage3_42[16],stage3_41[16],stage3_40[23]}
   );
   gpc2135_5 gpc4600 (
      {stage2_41[45], stage2_41[46], stage2_41[47], stage2_41[48], stage2_41[49]},
      {stage2_42[30], stage2_42[31], stage2_42[32]},
      {stage2_43[0]},
      {stage2_44[0], stage2_44[1]},
      {stage3_45[0],stage3_44[2],stage3_43[17],stage3_42[17],stage3_41[17]}
   );
   gpc1163_5 gpc4601 (
      {stage2_41[50], stage2_41[51], stage2_41[52]},
      {stage2_42[33], stage2_42[34], stage2_42[35], stage2_42[36], stage2_42[37], stage2_42[38]},
      {stage2_43[1]},
      {stage2_44[2]},
      {stage3_45[1],stage3_44[3],stage3_43[18],stage3_42[18],stage3_41[18]}
   );
   gpc1163_5 gpc4602 (
      {stage2_41[53], stage2_41[54], stage2_41[55]},
      {stage2_42[39], stage2_42[40], stage2_42[41], stage2_42[42], stage2_42[43], stage2_42[44]},
      {stage2_43[2]},
      {stage2_44[3]},
      {stage3_45[2],stage3_44[4],stage3_43[19],stage3_42[19],stage3_41[19]}
   );
   gpc1163_5 gpc4603 (
      {stage2_41[56], stage2_41[57], stage2_41[58]},
      {stage2_42[45], stage2_42[46], stage2_42[47], stage2_42[48], stage2_42[49], stage2_42[50]},
      {stage2_43[3]},
      {stage2_44[4]},
      {stage3_45[3],stage3_44[5],stage3_43[20],stage3_42[20],stage3_41[20]}
   );
   gpc606_5 gpc4604 (
      {stage2_41[59], stage2_41[60], stage2_41[61], stage2_41[62], stage2_41[63], stage2_41[64]},
      {stage2_43[4], stage2_43[5], stage2_43[6], stage2_43[7], stage2_43[8], stage2_43[9]},
      {stage3_45[4],stage3_44[6],stage3_43[21],stage3_42[21],stage3_41[21]}
   );
   gpc615_5 gpc4605 (
      {stage2_41[65], stage2_41[66], stage2_41[67], stage2_41[68], stage2_41[69]},
      {stage2_42[51]},
      {stage2_43[10], stage2_43[11], stage2_43[12], stage2_43[13], stage2_43[14], stage2_43[15]},
      {stage3_45[5],stage3_44[7],stage3_43[22],stage3_42[22],stage3_41[22]}
   );
   gpc615_5 gpc4606 (
      {stage2_41[70], stage2_41[71], stage2_41[72], stage2_41[73], stage2_41[74]},
      {stage2_42[52]},
      {stage2_43[16], stage2_43[17], stage2_43[18], stage2_43[19], stage2_43[20], stage2_43[21]},
      {stage3_45[6],stage3_44[8],stage3_43[23],stage3_42[23],stage3_41[23]}
   );
   gpc615_5 gpc4607 (
      {stage2_42[53], stage2_42[54], stage2_42[55], stage2_42[56], stage2_42[57]},
      {stage2_43[22]},
      {stage2_44[5], stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10]},
      {stage3_46[0],stage3_45[7],stage3_44[9],stage3_43[24],stage3_42[24]}
   );
   gpc606_5 gpc4608 (
      {stage2_43[23], stage2_43[24], stage2_43[25], stage2_43[26], stage2_43[27], stage2_43[28]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[1],stage3_45[8],stage3_44[10],stage3_43[25]}
   );
   gpc615_5 gpc4609 (
      {stage2_43[29], stage2_43[30], stage2_43[31], stage2_43[32], stage2_43[33]},
      {stage2_44[11]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[2],stage3_45[9],stage3_44[11],stage3_43[26]}
   );
   gpc615_5 gpc4610 (
      {stage2_43[34], stage2_43[35], stage2_43[36], stage2_43[37], stage2_43[38]},
      {stage2_44[12]},
      {stage2_45[12], stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage3_47[2],stage3_46[3],stage3_45[10],stage3_44[12],stage3_43[27]}
   );
   gpc615_5 gpc4611 (
      {stage2_43[39], stage2_43[40], stage2_43[41], stage2_43[42], stage2_43[43]},
      {stage2_44[13]},
      {stage2_45[18], stage2_45[19], stage2_45[20], stage2_45[21], stage2_45[22], stage2_45[23]},
      {stage3_47[3],stage3_46[4],stage3_45[11],stage3_44[13],stage3_43[28]}
   );
   gpc615_5 gpc4612 (
      {stage2_43[44], stage2_43[45], stage2_43[46], stage2_43[47], stage2_43[48]},
      {stage2_44[14]},
      {stage2_45[24], stage2_45[25], stage2_45[26], stage2_45[27], stage2_45[28], stage2_45[29]},
      {stage3_47[4],stage3_46[5],stage3_45[12],stage3_44[14],stage3_43[29]}
   );
   gpc615_5 gpc4613 (
      {stage2_43[49], stage2_43[50], stage2_43[51], stage2_43[52], stage2_43[53]},
      {stage2_44[15]},
      {stage2_45[30], stage2_45[31], stage2_45[32], stage2_45[33], stage2_45[34], stage2_45[35]},
      {stage3_47[5],stage3_46[6],stage3_45[13],stage3_44[15],stage3_43[30]}
   );
   gpc606_5 gpc4614 (
      {stage2_44[16], stage2_44[17], stage2_44[18], stage2_44[19], stage2_44[20], stage2_44[21]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[6],stage3_46[7],stage3_45[14],stage3_44[16]}
   );
   gpc606_5 gpc4615 (
      {stage2_44[22], stage2_44[23], stage2_44[24], stage2_44[25], stage2_44[26], stage2_44[27]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[7],stage3_46[8],stage3_45[15],stage3_44[17]}
   );
   gpc606_5 gpc4616 (
      {stage2_44[28], stage2_44[29], stage2_44[30], stage2_44[31], stage2_44[32], stage2_44[33]},
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage3_48[2],stage3_47[8],stage3_46[9],stage3_45[16],stage3_44[18]}
   );
   gpc606_5 gpc4617 (
      {stage2_44[34], stage2_44[35], stage2_44[36], stage2_44[37], stage2_44[38], stage2_44[39]},
      {stage2_46[18], stage2_46[19], stage2_46[20], stage2_46[21], stage2_46[22], stage2_46[23]},
      {stage3_48[3],stage3_47[9],stage3_46[10],stage3_45[17],stage3_44[19]}
   );
   gpc606_5 gpc4618 (
      {stage2_44[40], stage2_44[41], stage2_44[42], stage2_44[43], stage2_44[44], stage2_44[45]},
      {stage2_46[24], stage2_46[25], stage2_46[26], stage2_46[27], stage2_46[28], stage2_46[29]},
      {stage3_48[4],stage3_47[10],stage3_46[11],stage3_45[18],stage3_44[20]}
   );
   gpc606_5 gpc4619 (
      {stage2_44[46], stage2_44[47], stage2_44[48], stage2_44[49], stage2_44[50], stage2_44[51]},
      {stage2_46[30], stage2_46[31], stage2_46[32], stage2_46[33], stage2_46[34], stage2_46[35]},
      {stage3_48[5],stage3_47[11],stage3_46[12],stage3_45[19],stage3_44[21]}
   );
   gpc615_5 gpc4620 (
      {stage2_45[36], stage2_45[37], stage2_45[38], stage2_45[39], stage2_45[40]},
      {stage2_46[36]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[6],stage3_47[12],stage3_46[13],stage3_45[20]}
   );
   gpc615_5 gpc4621 (
      {stage2_45[41], stage2_45[42], stage2_45[43], stage2_45[44], stage2_45[45]},
      {stage2_46[37]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[7],stage3_47[13],stage3_46[14],stage3_45[21]}
   );
   gpc615_5 gpc4622 (
      {stage2_45[46], stage2_45[47], stage2_45[48], stage2_45[49], stage2_45[50]},
      {stage2_46[38]},
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17]},
      {stage3_49[2],stage3_48[8],stage3_47[14],stage3_46[15],stage3_45[22]}
   );
   gpc615_5 gpc4623 (
      {stage2_45[51], stage2_45[52], stage2_45[53], stage2_45[54], stage2_45[55]},
      {stage2_46[39]},
      {stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21], stage2_47[22], stage2_47[23]},
      {stage3_49[3],stage3_48[9],stage3_47[15],stage3_46[16],stage3_45[23]}
   );
   gpc615_5 gpc4624 (
      {stage2_45[56], stage2_45[57], stage2_45[58], stage2_45[59], stage2_45[60]},
      {stage2_46[40]},
      {stage2_47[24], stage2_47[25], stage2_47[26], stage2_47[27], stage2_47[28], stage2_47[29]},
      {stage3_49[4],stage3_48[10],stage3_47[16],stage3_46[17],stage3_45[24]}
   );
   gpc615_5 gpc4625 (
      {stage2_45[61], stage2_45[62], stage2_45[63], stage2_45[64], stage2_45[65]},
      {stage2_46[41]},
      {stage2_47[30], stage2_47[31], stage2_47[32], stage2_47[33], stage2_47[34], stage2_47[35]},
      {stage3_49[5],stage3_48[11],stage3_47[17],stage3_46[18],stage3_45[25]}
   );
   gpc615_5 gpc4626 (
      {stage2_47[36], stage2_47[37], stage2_47[38], stage2_47[39], stage2_47[40]},
      {stage2_48[0]},
      {stage2_49[0], stage2_49[1], stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5]},
      {stage3_51[0],stage3_50[0],stage3_49[6],stage3_48[12],stage3_47[18]}
   );
   gpc615_5 gpc4627 (
      {stage2_47[41], stage2_47[42], stage2_47[43], stage2_47[44], stage2_47[45]},
      {stage2_48[1]},
      {stage2_49[6], stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11]},
      {stage3_51[1],stage3_50[1],stage3_49[7],stage3_48[13],stage3_47[19]}
   );
   gpc615_5 gpc4628 (
      {stage2_47[46], stage2_47[47], stage2_47[48], stage2_47[49], stage2_47[50]},
      {stage2_48[2]},
      {stage2_49[12], stage2_49[13], stage2_49[14], stage2_49[15], stage2_49[16], stage2_49[17]},
      {stage3_51[2],stage3_50[2],stage3_49[8],stage3_48[14],stage3_47[20]}
   );
   gpc615_5 gpc4629 (
      {stage2_47[51], stage2_47[52], stage2_47[53], stage2_47[54], stage2_47[55]},
      {stage2_48[3]},
      {stage2_49[18], stage2_49[19], stage2_49[20], stage2_49[21], stage2_49[22], stage2_49[23]},
      {stage3_51[3],stage3_50[3],stage3_49[9],stage3_48[15],stage3_47[21]}
   );
   gpc615_5 gpc4630 (
      {stage2_47[56], stage2_47[57], stage2_47[58], stage2_47[59], stage2_47[60]},
      {stage2_48[4]},
      {stage2_49[24], stage2_49[25], stage2_49[26], stage2_49[27], stage2_49[28], stage2_49[29]},
      {stage3_51[4],stage3_50[4],stage3_49[10],stage3_48[16],stage3_47[22]}
   );
   gpc606_5 gpc4631 (
      {stage2_48[5], stage2_48[6], stage2_48[7], stage2_48[8], stage2_48[9], stage2_48[10]},
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage3_52[0],stage3_51[5],stage3_50[5],stage3_49[11],stage3_48[17]}
   );
   gpc606_5 gpc4632 (
      {stage2_48[11], stage2_48[12], stage2_48[13], stage2_48[14], stage2_48[15], stage2_48[16]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage3_52[1],stage3_51[6],stage3_50[6],stage3_49[12],stage3_48[18]}
   );
   gpc615_5 gpc4633 (
      {stage2_48[17], stage2_48[18], stage2_48[19], stage2_48[20], stage2_48[21]},
      {stage2_49[30]},
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16], stage2_50[17]},
      {stage3_52[2],stage3_51[7],stage3_50[7],stage3_49[13],stage3_48[19]}
   );
   gpc615_5 gpc4634 (
      {stage2_48[22], stage2_48[23], stage2_48[24], stage2_48[25], stage2_48[26]},
      {stage2_49[31]},
      {stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21], stage2_50[22], stage2_50[23]},
      {stage3_52[3],stage3_51[8],stage3_50[8],stage3_49[14],stage3_48[20]}
   );
   gpc615_5 gpc4635 (
      {stage2_48[27], stage2_48[28], stage2_48[29], stage2_48[30], stage2_48[31]},
      {stage2_49[32]},
      {stage2_50[24], stage2_50[25], stage2_50[26], stage2_50[27], stage2_50[28], stage2_50[29]},
      {stage3_52[4],stage3_51[9],stage3_50[9],stage3_49[15],stage3_48[21]}
   );
   gpc615_5 gpc4636 (
      {stage2_48[32], stage2_48[33], stage2_48[34], stage2_48[35], stage2_48[36]},
      {stage2_49[33]},
      {stage2_50[30], stage2_50[31], stage2_50[32], stage2_50[33], stage2_50[34], stage2_50[35]},
      {stage3_52[5],stage3_51[10],stage3_50[10],stage3_49[16],stage3_48[22]}
   );
   gpc615_5 gpc4637 (
      {stage2_48[37], stage2_48[38], stage2_48[39], stage2_48[40], stage2_48[41]},
      {stage2_49[34]},
      {stage2_50[36], stage2_50[37], stage2_50[38], stage2_50[39], stage2_50[40], stage2_50[41]},
      {stage3_52[6],stage3_51[11],stage3_50[11],stage3_49[17],stage3_48[23]}
   );
   gpc117_4 gpc4638 (
      {stage2_49[35], stage2_49[36], stage2_49[37], stage2_49[38], stage2_49[39], stage2_49[40], stage2_49[41]},
      {stage2_50[42]},
      {stage2_51[0]},
      {stage3_52[7],stage3_51[12],stage3_50[12],stage3_49[18]}
   );
   gpc117_4 gpc4639 (
      {stage2_49[42], stage2_49[43], stage2_49[44], stage2_49[45], stage2_49[46], stage2_49[47], stage2_49[48]},
      {stage2_50[43]},
      {stage2_51[1]},
      {stage3_52[8],stage3_51[13],stage3_50[13],stage3_49[19]}
   );
   gpc117_4 gpc4640 (
      {stage2_49[49], stage2_49[50], stage2_49[51], stage2_49[52], stage2_49[53], stage2_49[54], stage2_49[55]},
      {stage2_50[44]},
      {stage2_51[2]},
      {stage3_52[9],stage3_51[14],stage3_50[14],stage3_49[20]}
   );
   gpc117_4 gpc4641 (
      {stage2_49[56], stage2_49[57], stage2_49[58], stage2_49[59], stage2_49[60], stage2_49[61], stage2_49[62]},
      {stage2_50[45]},
      {stage2_51[3]},
      {stage3_52[10],stage3_51[15],stage3_50[15],stage3_49[21]}
   );
   gpc117_4 gpc4642 (
      {stage2_49[63], stage2_49[64], stage2_49[65], stage2_49[66], stage2_49[67], stage2_49[68], stage2_49[69]},
      {stage2_50[46]},
      {stage2_51[4]},
      {stage3_52[11],stage3_51[16],stage3_50[16],stage3_49[22]}
   );
   gpc615_5 gpc4643 (
      {stage2_50[47], stage2_50[48], stage2_50[49], stage2_50[50], stage2_50[51]},
      {stage2_51[5]},
      {stage2_52[0], stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage3_54[0],stage3_53[0],stage3_52[12],stage3_51[17],stage3_50[17]}
   );
   gpc615_5 gpc4644 (
      {stage2_50[52], stage2_50[53], stage2_50[54], stage2_50[55], stage2_50[56]},
      {stage2_51[6]},
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10], stage2_52[11]},
      {stage3_54[1],stage3_53[1],stage3_52[13],stage3_51[18],stage3_50[18]}
   );
   gpc606_5 gpc4645 (
      {stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11], stage2_51[12]},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[2],stage3_53[2],stage3_52[14],stage3_51[19]}
   );
   gpc606_5 gpc4646 (
      {stage2_51[13], stage2_51[14], stage2_51[15], stage2_51[16], stage2_51[17], stage2_51[18]},
      {stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11]},
      {stage3_55[1],stage3_54[3],stage3_53[3],stage3_52[15],stage3_51[20]}
   );
   gpc606_5 gpc4647 (
      {stage2_51[19], stage2_51[20], stage2_51[21], stage2_51[22], stage2_51[23], stage2_51[24]},
      {stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16], stage2_53[17]},
      {stage3_55[2],stage3_54[4],stage3_53[4],stage3_52[16],stage3_51[21]}
   );
   gpc606_5 gpc4648 (
      {stage2_51[25], stage2_51[26], stage2_51[27], stage2_51[28], stage2_51[29], stage2_51[30]},
      {stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21], stage2_53[22], stage2_53[23]},
      {stage3_55[3],stage3_54[5],stage3_53[5],stage3_52[17],stage3_51[22]}
   );
   gpc606_5 gpc4649 (
      {stage2_51[31], stage2_51[32], stage2_51[33], stage2_51[34], stage2_51[35], stage2_51[36]},
      {stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27], stage2_53[28], stage2_53[29]},
      {stage3_55[4],stage3_54[6],stage3_53[6],stage3_52[18],stage3_51[23]}
   );
   gpc615_5 gpc4650 (
      {stage2_51[37], stage2_51[38], stage2_51[39], stage2_51[40], stage2_51[41]},
      {stage2_52[12]},
      {stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33], stage2_53[34], stage2_53[35]},
      {stage3_55[5],stage3_54[7],stage3_53[7],stage3_52[19],stage3_51[24]}
   );
   gpc615_5 gpc4651 (
      {stage2_51[42], stage2_51[43], stage2_51[44], stage2_51[45], stage2_51[46]},
      {stage2_52[13]},
      {stage2_53[36], stage2_53[37], stage2_53[38], stage2_53[39], stage2_53[40], stage2_53[41]},
      {stage3_55[6],stage3_54[8],stage3_53[8],stage3_52[20],stage3_51[25]}
   );
   gpc615_5 gpc4652 (
      {stage2_51[47], stage2_51[48], stage2_51[49], stage2_51[50], stage2_51[51]},
      {stage2_52[14]},
      {stage2_53[42], stage2_53[43], stage2_53[44], stage2_53[45], stage2_53[46], stage2_53[47]},
      {stage3_55[7],stage3_54[9],stage3_53[9],stage3_52[21],stage3_51[26]}
   );
   gpc623_5 gpc4653 (
      {stage2_51[52], stage2_51[53], stage2_51[54]},
      {stage2_52[15], stage2_52[16]},
      {stage2_53[48], stage2_53[49], stage2_53[50], stage2_53[51], stage2_53[52], stage2_53[53]},
      {stage3_55[8],stage3_54[10],stage3_53[10],stage3_52[22],stage3_51[27]}
   );
   gpc623_5 gpc4654 (
      {stage2_51[55], stage2_51[56], stage2_51[57]},
      {stage2_52[17], stage2_52[18]},
      {stage2_53[54], stage2_53[55], stage2_53[56], stage2_53[57], stage2_53[58], stage2_53[59]},
      {stage3_55[9],stage3_54[11],stage3_53[11],stage3_52[23],stage3_51[28]}
   );
   gpc623_5 gpc4655 (
      {stage2_51[58], stage2_51[59], stage2_51[60]},
      {stage2_52[19], stage2_52[20]},
      {stage2_53[60], stage2_53[61], stage2_53[62], stage2_53[63], stage2_53[64], stage2_53[65]},
      {stage3_55[10],stage3_54[12],stage3_53[12],stage3_52[24],stage3_51[29]}
   );
   gpc606_5 gpc4656 (
      {stage2_52[21], stage2_52[22], stage2_52[23], stage2_52[24], stage2_52[25], stage2_52[26]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[11],stage3_54[13],stage3_53[13],stage3_52[25]}
   );
   gpc606_5 gpc4657 (
      {stage2_52[27], stage2_52[28], stage2_52[29], stage2_52[30], stage2_52[31], stage2_52[32]},
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage3_56[1],stage3_55[12],stage3_54[14],stage3_53[14],stage3_52[26]}
   );
   gpc606_5 gpc4658 (
      {stage2_52[33], stage2_52[34], stage2_52[35], stage2_52[36], stage2_52[37], stage2_52[38]},
      {stage2_54[12], stage2_54[13], stage2_54[14], stage2_54[15], stage2_54[16], stage2_54[17]},
      {stage3_56[2],stage3_55[13],stage3_54[15],stage3_53[15],stage3_52[27]}
   );
   gpc606_5 gpc4659 (
      {stage2_54[18], stage2_54[19], stage2_54[20], stage2_54[21], stage2_54[22], stage2_54[23]},
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5]},
      {stage3_58[0],stage3_57[0],stage3_56[3],stage3_55[14],stage3_54[16]}
   );
   gpc606_5 gpc4660 (
      {stage2_54[24], stage2_54[25], stage2_54[26], stage2_54[27], stage2_54[28], stage2_54[29]},
      {stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9], stage2_56[10], stage2_56[11]},
      {stage3_58[1],stage3_57[1],stage3_56[4],stage3_55[15],stage3_54[17]}
   );
   gpc606_5 gpc4661 (
      {stage2_54[30], stage2_54[31], stage2_54[32], stage2_54[33], stage2_54[34], stage2_54[35]},
      {stage2_56[12], stage2_56[13], stage2_56[14], stage2_56[15], stage2_56[16], stage2_56[17]},
      {stage3_58[2],stage3_57[2],stage3_56[5],stage3_55[16],stage3_54[18]}
   );
   gpc606_5 gpc4662 (
      {stage2_54[36], stage2_54[37], stage2_54[38], stage2_54[39], stage2_54[40], stage2_54[41]},
      {stage2_56[18], stage2_56[19], stage2_56[20], stage2_56[21], stage2_56[22], stage2_56[23]},
      {stage3_58[3],stage3_57[3],stage3_56[6],stage3_55[17],stage3_54[19]}
   );
   gpc606_5 gpc4663 (
      {stage2_54[42], stage2_54[43], stage2_54[44], stage2_54[45], stage2_54[46], stage2_54[47]},
      {stage2_56[24], stage2_56[25], stage2_56[26], stage2_56[27], stage2_56[28], stage2_56[29]},
      {stage3_58[4],stage3_57[4],stage3_56[7],stage3_55[18],stage3_54[20]}
   );
   gpc606_5 gpc4664 (
      {stage2_54[48], stage2_54[49], stage2_54[50], stage2_54[51], stage2_54[52], stage2_54[53]},
      {stage2_56[30], stage2_56[31], stage2_56[32], stage2_56[33], stage2_56[34], stage2_56[35]},
      {stage3_58[5],stage3_57[5],stage3_56[8],stage3_55[19],stage3_54[21]}
   );
   gpc606_5 gpc4665 (
      {stage2_54[54], stage2_54[55], stage2_54[56], stage2_54[57], stage2_54[58], stage2_54[59]},
      {stage2_56[36], stage2_56[37], stage2_56[38], stage2_56[39], stage2_56[40], stage2_56[41]},
      {stage3_58[6],stage3_57[6],stage3_56[9],stage3_55[20],stage3_54[22]}
   );
   gpc606_5 gpc4666 (
      {stage2_54[60], stage2_54[61], stage2_54[62], stage2_54[63], stage2_54[64], stage2_54[65]},
      {stage2_56[42], stage2_56[43], stage2_56[44], stage2_56[45], stage2_56[46], stage2_56[47]},
      {stage3_58[7],stage3_57[7],stage3_56[10],stage3_55[21],stage3_54[23]}
   );
   gpc606_5 gpc4667 (
      {stage2_54[66], stage2_54[67], stage2_54[68], stage2_54[69], stage2_54[70], stage2_54[71]},
      {stage2_56[48], stage2_56[49], stage2_56[50], stage2_56[51], stage2_56[52], stage2_56[53]},
      {stage3_58[8],stage3_57[8],stage3_56[11],stage3_55[22],stage3_54[24]}
   );
   gpc615_5 gpc4668 (
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4]},
      {stage2_56[54]},
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5]},
      {stage3_59[0],stage3_58[9],stage3_57[9],stage3_56[12],stage3_55[23]}
   );
   gpc615_5 gpc4669 (
      {stage2_55[5], stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9]},
      {stage2_56[55]},
      {stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10], stage2_57[11]},
      {stage3_59[1],stage3_58[10],stage3_57[10],stage3_56[13],stage3_55[24]}
   );
   gpc615_5 gpc4670 (
      {stage2_55[10], stage2_55[11], stage2_55[12], stage2_55[13], stage2_55[14]},
      {stage2_56[56]},
      {stage2_57[12], stage2_57[13], stage2_57[14], stage2_57[15], stage2_57[16], stage2_57[17]},
      {stage3_59[2],stage3_58[11],stage3_57[11],stage3_56[14],stage3_55[25]}
   );
   gpc615_5 gpc4671 (
      {stage2_55[15], stage2_55[16], stage2_55[17], stage2_55[18], stage2_55[19]},
      {stage2_56[57]},
      {stage2_57[18], stage2_57[19], stage2_57[20], stage2_57[21], stage2_57[22], stage2_57[23]},
      {stage3_59[3],stage3_58[12],stage3_57[12],stage3_56[15],stage3_55[26]}
   );
   gpc615_5 gpc4672 (
      {stage2_55[20], stage2_55[21], stage2_55[22], stage2_55[23], stage2_55[24]},
      {stage2_56[58]},
      {stage2_57[24], stage2_57[25], stage2_57[26], stage2_57[27], stage2_57[28], stage2_57[29]},
      {stage3_59[4],stage3_58[13],stage3_57[13],stage3_56[16],stage3_55[27]}
   );
   gpc615_5 gpc4673 (
      {stage2_55[25], stage2_55[26], stage2_55[27], stage2_55[28], stage2_55[29]},
      {stage2_56[59]},
      {stage2_57[30], stage2_57[31], stage2_57[32], stage2_57[33], stage2_57[34], stage2_57[35]},
      {stage3_59[5],stage3_58[14],stage3_57[14],stage3_56[17],stage3_55[28]}
   );
   gpc615_5 gpc4674 (
      {stage2_55[30], stage2_55[31], stage2_55[32], stage2_55[33], stage2_55[34]},
      {stage2_56[60]},
      {stage2_57[36], stage2_57[37], stage2_57[38], stage2_57[39], stage2_57[40], stage2_57[41]},
      {stage3_59[6],stage3_58[15],stage3_57[15],stage3_56[18],stage3_55[29]}
   );
   gpc606_5 gpc4675 (
      {stage2_56[61], stage2_56[62], stage2_56[63], stage2_56[64], stage2_56[65], stage2_56[66]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[7],stage3_58[16],stage3_57[16],stage3_56[19]}
   );
   gpc606_5 gpc4676 (
      {stage2_57[42], stage2_57[43], stage2_57[44], stage2_57[45], stage2_57[46], stage2_57[47]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[1],stage3_59[8],stage3_58[17],stage3_57[17]}
   );
   gpc606_5 gpc4677 (
      {stage2_57[48], stage2_57[49], stage2_57[50], stage2_57[51], stage2_57[52], stage2_57[53]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[2],stage3_59[9],stage3_58[18],stage3_57[18]}
   );
   gpc606_5 gpc4678 (
      {stage2_57[54], stage2_57[55], stage2_57[56], stage2_57[57], stage2_57[58], stage2_57[59]},
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17]},
      {stage3_61[2],stage3_60[3],stage3_59[10],stage3_58[19],stage3_57[19]}
   );
   gpc606_5 gpc4679 (
      {stage2_57[60], stage2_57[61], stage2_57[62], stage2_57[63], stage2_57[64], stage2_57[65]},
      {stage2_59[18], stage2_59[19], stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23]},
      {stage3_61[3],stage3_60[4],stage3_59[11],stage3_58[20],stage3_57[20]}
   );
   gpc606_5 gpc4680 (
      {stage2_57[66], stage2_57[67], stage2_57[68], stage2_57[69], stage2_57[70], stage2_57[71]},
      {stage2_59[24], stage2_59[25], stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29]},
      {stage3_61[4],stage3_60[5],stage3_59[12],stage3_58[21],stage3_57[21]}
   );
   gpc606_5 gpc4681 (
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage2_60[0], stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5]},
      {stage3_62[0],stage3_61[5],stage3_60[6],stage3_59[13],stage3_58[22]}
   );
   gpc606_5 gpc4682 (
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage2_60[6], stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11]},
      {stage3_62[1],stage3_61[6],stage3_60[7],stage3_59[14],stage3_58[23]}
   );
   gpc606_5 gpc4683 (
      {stage2_58[18], stage2_58[19], stage2_58[20], stage2_58[21], stage2_58[22], stage2_58[23]},
      {stage2_60[12], stage2_60[13], stage2_60[14], stage2_60[15], stage2_60[16], stage2_60[17]},
      {stage3_62[2],stage3_61[7],stage3_60[8],stage3_59[15],stage3_58[24]}
   );
   gpc606_5 gpc4684 (
      {stage2_58[24], stage2_58[25], stage2_58[26], stage2_58[27], stage2_58[28], stage2_58[29]},
      {stage2_60[18], stage2_60[19], stage2_60[20], stage2_60[21], stage2_60[22], stage2_60[23]},
      {stage3_62[3],stage3_61[8],stage3_60[9],stage3_59[16],stage3_58[25]}
   );
   gpc606_5 gpc4685 (
      {stage2_58[30], stage2_58[31], stage2_58[32], stage2_58[33], stage2_58[34], stage2_58[35]},
      {stage2_60[24], stage2_60[25], stage2_60[26], stage2_60[27], stage2_60[28], stage2_60[29]},
      {stage3_62[4],stage3_61[9],stage3_60[10],stage3_59[17],stage3_58[26]}
   );
   gpc606_5 gpc4686 (
      {stage2_58[36], stage2_58[37], stage2_58[38], stage2_58[39], stage2_58[40], stage2_58[41]},
      {stage2_60[30], stage2_60[31], stage2_60[32], stage2_60[33], stage2_60[34], stage2_60[35]},
      {stage3_62[5],stage3_61[10],stage3_60[11],stage3_59[18],stage3_58[27]}
   );
   gpc606_5 gpc4687 (
      {stage2_58[42], stage2_58[43], stage2_58[44], stage2_58[45], stage2_58[46], stage2_58[47]},
      {stage2_60[36], stage2_60[37], stage2_60[38], stage2_60[39], stage2_60[40], stage2_60[41]},
      {stage3_62[6],stage3_61[11],stage3_60[12],stage3_59[19],stage3_58[28]}
   );
   gpc606_5 gpc4688 (
      {stage2_59[30], stage2_59[31], stage2_59[32], stage2_59[33], stage2_59[34], stage2_59[35]},
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage3_63[0],stage3_62[7],stage3_61[12],stage3_60[13],stage3_59[20]}
   );
   gpc606_5 gpc4689 (
      {stage2_61[6], stage2_61[7], stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[0],stage3_63[1],stage3_62[8],stage3_61[13]}
   );
   gpc606_5 gpc4690 (
      {stage2_61[12], stage2_61[13], stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17]},
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11]},
      {stage3_65[1],stage3_64[1],stage3_63[2],stage3_62[9],stage3_61[14]}
   );
   gpc606_5 gpc4691 (
      {stage2_61[18], stage2_61[19], stage2_61[20], stage2_61[21], stage2_61[22], stage2_61[23]},
      {stage2_63[12], stage2_63[13], stage2_63[14], stage2_63[15], stage2_63[16], stage2_63[17]},
      {stage3_65[2],stage3_64[2],stage3_63[3],stage3_62[10],stage3_61[15]}
   );
   gpc606_5 gpc4692 (
      {stage2_61[24], stage2_61[25], stage2_61[26], stage2_61[27], stage2_61[28], stage2_61[29]},
      {stage2_63[18], stage2_63[19], stage2_63[20], stage2_63[21], stage2_63[22], stage2_63[23]},
      {stage3_65[3],stage3_64[3],stage3_63[4],stage3_62[11],stage3_61[16]}
   );
   gpc606_5 gpc4693 (
      {stage2_61[30], stage2_61[31], stage2_61[32], stage2_61[33], stage2_61[34], stage2_61[35]},
      {stage2_63[24], stage2_63[25], stage2_63[26], stage2_63[27], stage2_63[28], stage2_63[29]},
      {stage3_65[4],stage3_64[4],stage3_63[5],stage3_62[12],stage3_61[17]}
   );
   gpc606_5 gpc4694 (
      {stage2_61[36], stage2_61[37], stage2_61[38], stage2_61[39], stage2_61[40], stage2_61[41]},
      {stage2_63[30], stage2_63[31], stage2_63[32], stage2_63[33], stage2_63[34], stage2_63[35]},
      {stage3_65[5],stage3_64[5],stage3_63[6],stage3_62[13],stage3_61[18]}
   );
   gpc606_5 gpc4695 (
      {stage2_61[42], stage2_61[43], stage2_61[44], stage2_61[45], stage2_61[46], stage2_61[47]},
      {stage2_63[36], stage2_63[37], stage2_63[38], stage2_63[39], stage2_63[40], stage2_63[41]},
      {stage3_65[6],stage3_64[6],stage3_63[7],stage3_62[14],stage3_61[19]}
   );
   gpc606_5 gpc4696 (
      {stage2_61[48], stage2_61[49], stage2_61[50], stage2_61[51], stage2_61[52], stage2_61[53]},
      {stage2_63[42], stage2_63[43], stage2_63[44], stage2_63[45], stage2_63[46], stage2_63[47]},
      {stage3_65[7],stage3_64[7],stage3_63[8],stage3_62[15],stage3_61[20]}
   );
   gpc1163_5 gpc4697 (
      {stage2_62[0], stage2_62[1], stage2_62[2]},
      {stage2_63[48], stage2_63[49], stage2_63[50], stage2_63[51], stage2_63[52], stage2_63[53]},
      {stage2_64[0]},
      {stage2_65[0]},
      {stage3_66[0],stage3_65[8],stage3_64[8],stage3_63[9],stage3_62[16]}
   );
   gpc1163_5 gpc4698 (
      {stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage2_63[54], stage2_63[55], stage2_63[56], stage2_63[57], stage2_63[58], stage2_63[59]},
      {stage2_64[1]},
      {stage2_65[1]},
      {stage3_66[1],stage3_65[9],stage3_64[9],stage3_63[10],stage3_62[17]}
   );
   gpc1163_5 gpc4699 (
      {stage2_62[6], stage2_62[7], stage2_62[8]},
      {stage2_63[60], stage2_63[61], stage2_63[62], stage2_63[63], stage2_63[64], stage2_63[65]},
      {stage2_64[2]},
      {stage2_65[2]},
      {stage3_66[2],stage3_65[10],stage3_64[10],stage3_63[11],stage3_62[18]}
   );
   gpc606_5 gpc4700 (
      {stage2_62[9], stage2_62[10], stage2_62[11], stage2_62[12], stage2_62[13], stage2_62[14]},
      {stage2_64[3], stage2_64[4], stage2_64[5], stage2_64[6], stage2_64[7], stage2_64[8]},
      {stage3_66[3],stage3_65[11],stage3_64[11],stage3_63[12],stage3_62[19]}
   );
   gpc606_5 gpc4701 (
      {stage2_62[15], stage2_62[16], stage2_62[17], stage2_62[18], stage2_62[19], stage2_62[20]},
      {stage2_64[9], stage2_64[10], stage2_64[11], stage2_64[12], stage2_64[13], stage2_64[14]},
      {stage3_66[4],stage3_65[12],stage3_64[12],stage3_63[13],stage3_62[20]}
   );
   gpc606_5 gpc4702 (
      {stage2_62[21], stage2_62[22], stage2_62[23], stage2_62[24], stage2_62[25], stage2_62[26]},
      {stage2_64[15], stage2_64[16], stage2_64[17], stage2_64[18], stage2_64[19], stage2_64[20]},
      {stage3_66[5],stage3_65[13],stage3_64[13],stage3_63[14],stage3_62[21]}
   );
   gpc606_5 gpc4703 (
      {stage2_62[27], stage2_62[28], stage2_62[29], stage2_62[30], stage2_62[31], stage2_62[32]},
      {stage2_64[21], stage2_64[22], stage2_64[23], stage2_64[24], stage2_64[25], stage2_64[26]},
      {stage3_66[6],stage3_65[14],stage3_64[14],stage3_63[15],stage3_62[22]}
   );
   gpc606_5 gpc4704 (
      {stage2_62[33], stage2_62[34], stage2_62[35], stage2_62[36], stage2_62[37], stage2_62[38]},
      {stage2_64[27], stage2_64[28], stage2_64[29], stage2_64[30], stage2_64[31], stage2_64[32]},
      {stage3_66[7],stage3_65[15],stage3_64[15],stage3_63[16],stage3_62[23]}
   );
   gpc606_5 gpc4705 (
      {stage2_62[39], stage2_62[40], stage2_62[41], stage2_62[42], stage2_62[43], stage2_62[44]},
      {stage2_64[33], stage2_64[34], stage2_64[35], stage2_64[36], stage2_64[37], stage2_64[38]},
      {stage3_66[8],stage3_65[16],stage3_64[16],stage3_63[17],stage3_62[24]}
   );
   gpc606_5 gpc4706 (
      {stage2_62[45], stage2_62[46], stage2_62[47], stage2_62[48], stage2_62[49], stage2_62[50]},
      {stage2_64[39], stage2_64[40], stage2_64[41], stage2_64[42], stage2_64[43], stage2_64[44]},
      {stage3_66[9],stage3_65[17],stage3_64[17],stage3_63[18],stage3_62[25]}
   );
   gpc606_5 gpc4707 (
      {stage2_65[3], stage2_65[4], stage2_65[5], stage2_65[6], stage2_65[7], stage2_65[8]},
      {stage2_67[0], stage2_67[1], stage2_67[2], stage2_67[3], stage2_67[4], stage2_67[5]},
      {stage3_69[0],stage3_68[0],stage3_67[0],stage3_66[10],stage3_65[18]}
   );
   gpc1_1 gpc4708 (
      {stage2_0[20]},
      {stage3_0[4]}
   );
   gpc1_1 gpc4709 (
      {stage2_0[21]},
      {stage3_0[5]}
   );
   gpc1_1 gpc4710 (
      {stage2_0[22]},
      {stage3_0[6]}
   );
   gpc1_1 gpc4711 (
      {stage2_0[23]},
      {stage3_0[7]}
   );
   gpc1_1 gpc4712 (
      {stage2_0[24]},
      {stage3_0[8]}
   );
   gpc1_1 gpc4713 (
      {stage2_0[25]},
      {stage3_0[9]}
   );
   gpc1_1 gpc4714 (
      {stage2_0[26]},
      {stage3_0[10]}
   );
   gpc1_1 gpc4715 (
      {stage2_0[27]},
      {stage3_0[11]}
   );
   gpc1_1 gpc4716 (
      {stage2_0[28]},
      {stage3_0[12]}
   );
   gpc1_1 gpc4717 (
      {stage2_0[29]},
      {stage3_0[13]}
   );
   gpc1_1 gpc4718 (
      {stage2_1[35]},
      {stage3_1[9]}
   );
   gpc1_1 gpc4719 (
      {stage2_1[36]},
      {stage3_1[10]}
   );
   gpc1_1 gpc4720 (
      {stage2_2[29]},
      {stage3_2[10]}
   );
   gpc1_1 gpc4721 (
      {stage2_2[30]},
      {stage3_2[11]}
   );
   gpc1_1 gpc4722 (
      {stage2_2[31]},
      {stage3_2[12]}
   );
   gpc1_1 gpc4723 (
      {stage2_2[32]},
      {stage3_2[13]}
   );
   gpc1_1 gpc4724 (
      {stage2_2[33]},
      {stage3_2[14]}
   );
   gpc1_1 gpc4725 (
      {stage2_2[34]},
      {stage3_2[15]}
   );
   gpc1_1 gpc4726 (
      {stage2_2[35]},
      {stage3_2[16]}
   );
   gpc1_1 gpc4727 (
      {stage2_2[36]},
      {stage3_2[17]}
   );
   gpc1_1 gpc4728 (
      {stage2_3[50]},
      {stage3_3[15]}
   );
   gpc1_1 gpc4729 (
      {stage2_3[51]},
      {stage3_3[16]}
   );
   gpc1_1 gpc4730 (
      {stage2_3[52]},
      {stage3_3[17]}
   );
   gpc1_1 gpc4731 (
      {stage2_3[53]},
      {stage3_3[18]}
   );
   gpc1_1 gpc4732 (
      {stage2_4[43]},
      {stage3_4[19]}
   );
   gpc1_1 gpc4733 (
      {stage2_4[44]},
      {stage3_4[20]}
   );
   gpc1_1 gpc4734 (
      {stage2_5[26]},
      {stage3_5[15]}
   );
   gpc1_1 gpc4735 (
      {stage2_5[27]},
      {stage3_5[16]}
   );
   gpc1_1 gpc4736 (
      {stage2_5[28]},
      {stage3_5[17]}
   );
   gpc1_1 gpc4737 (
      {stage2_5[29]},
      {stage3_5[18]}
   );
   gpc1_1 gpc4738 (
      {stage2_5[30]},
      {stage3_5[19]}
   );
   gpc1_1 gpc4739 (
      {stage2_5[31]},
      {stage3_5[20]}
   );
   gpc1_1 gpc4740 (
      {stage2_5[32]},
      {stage3_5[21]}
   );
   gpc1_1 gpc4741 (
      {stage2_5[33]},
      {stage3_5[22]}
   );
   gpc1_1 gpc4742 (
      {stage2_5[34]},
      {stage3_5[23]}
   );
   gpc1_1 gpc4743 (
      {stage2_5[35]},
      {stage3_5[24]}
   );
   gpc1_1 gpc4744 (
      {stage2_5[36]},
      {stage3_5[25]}
   );
   gpc1_1 gpc4745 (
      {stage2_5[37]},
      {stage3_5[26]}
   );
   gpc1_1 gpc4746 (
      {stage2_5[38]},
      {stage3_5[27]}
   );
   gpc1_1 gpc4747 (
      {stage2_5[39]},
      {stage3_5[28]}
   );
   gpc1_1 gpc4748 (
      {stage2_5[40]},
      {stage3_5[29]}
   );
   gpc1_1 gpc4749 (
      {stage2_5[41]},
      {stage3_5[30]}
   );
   gpc1_1 gpc4750 (
      {stage2_5[42]},
      {stage3_5[31]}
   );
   gpc1_1 gpc4751 (
      {stage2_5[43]},
      {stage3_5[32]}
   );
   gpc1_1 gpc4752 (
      {stage2_5[44]},
      {stage3_5[33]}
   );
   gpc1_1 gpc4753 (
      {stage2_5[45]},
      {stage3_5[34]}
   );
   gpc1_1 gpc4754 (
      {stage2_6[49]},
      {stage3_6[14]}
   );
   gpc1_1 gpc4755 (
      {stage2_6[50]},
      {stage3_6[15]}
   );
   gpc1_1 gpc4756 (
      {stage2_6[51]},
      {stage3_6[16]}
   );
   gpc1_1 gpc4757 (
      {stage2_7[35]},
      {stage3_7[20]}
   );
   gpc1_1 gpc4758 (
      {stage2_7[36]},
      {stage3_7[21]}
   );
   gpc1_1 gpc4759 (
      {stage2_7[37]},
      {stage3_7[22]}
   );
   gpc1_1 gpc4760 (
      {stage2_7[38]},
      {stage3_7[23]}
   );
   gpc1_1 gpc4761 (
      {stage2_7[39]},
      {stage3_7[24]}
   );
   gpc1_1 gpc4762 (
      {stage2_7[40]},
      {stage3_7[25]}
   );
   gpc1_1 gpc4763 (
      {stage2_7[41]},
      {stage3_7[26]}
   );
   gpc1_1 gpc4764 (
      {stage2_7[42]},
      {stage3_7[27]}
   );
   gpc1_1 gpc4765 (
      {stage2_10[60]},
      {stage3_10[23]}
   );
   gpc1_1 gpc4766 (
      {stage2_10[61]},
      {stage3_10[24]}
   );
   gpc1_1 gpc4767 (
      {stage2_10[62]},
      {stage3_10[25]}
   );
   gpc1_1 gpc4768 (
      {stage2_10[63]},
      {stage3_10[26]}
   );
   gpc1_1 gpc4769 (
      {stage2_10[64]},
      {stage3_10[27]}
   );
   gpc1_1 gpc4770 (
      {stage2_10[65]},
      {stage3_10[28]}
   );
   gpc1_1 gpc4771 (
      {stage2_10[66]},
      {stage3_10[29]}
   );
   gpc1_1 gpc4772 (
      {stage2_10[67]},
      {stage3_10[30]}
   );
   gpc1_1 gpc4773 (
      {stage2_10[68]},
      {stage3_10[31]}
   );
   gpc1_1 gpc4774 (
      {stage2_10[69]},
      {stage3_10[32]}
   );
   gpc1_1 gpc4775 (
      {stage2_11[43]},
      {stage3_11[25]}
   );
   gpc1_1 gpc4776 (
      {stage2_11[44]},
      {stage3_11[26]}
   );
   gpc1_1 gpc4777 (
      {stage2_11[45]},
      {stage3_11[27]}
   );
   gpc1_1 gpc4778 (
      {stage2_11[46]},
      {stage3_11[28]}
   );
   gpc1_1 gpc4779 (
      {stage2_11[47]},
      {stage3_11[29]}
   );
   gpc1_1 gpc4780 (
      {stage2_11[48]},
      {stage3_11[30]}
   );
   gpc1_1 gpc4781 (
      {stage2_12[47]},
      {stage3_12[18]}
   );
   gpc1_1 gpc4782 (
      {stage2_12[48]},
      {stage3_12[19]}
   );
   gpc1_1 gpc4783 (
      {stage2_12[49]},
      {stage3_12[20]}
   );
   gpc1_1 gpc4784 (
      {stage2_12[50]},
      {stage3_12[21]}
   );
   gpc1_1 gpc4785 (
      {stage2_12[51]},
      {stage3_12[22]}
   );
   gpc1_1 gpc4786 (
      {stage2_12[52]},
      {stage3_12[23]}
   );
   gpc1_1 gpc4787 (
      {stage2_12[53]},
      {stage3_12[24]}
   );
   gpc1_1 gpc4788 (
      {stage2_13[60]},
      {stage3_13[20]}
   );
   gpc1_1 gpc4789 (
      {stage2_13[61]},
      {stage3_13[21]}
   );
   gpc1_1 gpc4790 (
      {stage2_13[62]},
      {stage3_13[22]}
   );
   gpc1_1 gpc4791 (
      {stage2_13[63]},
      {stage3_13[23]}
   );
   gpc1_1 gpc4792 (
      {stage2_14[42]},
      {stage3_14[24]}
   );
   gpc1_1 gpc4793 (
      {stage2_14[43]},
      {stage3_14[25]}
   );
   gpc1_1 gpc4794 (
      {stage2_14[44]},
      {stage3_14[26]}
   );
   gpc1_1 gpc4795 (
      {stage2_15[55]},
      {stage3_15[22]}
   );
   gpc1_1 gpc4796 (
      {stage2_15[56]},
      {stage3_15[23]}
   );
   gpc1_1 gpc4797 (
      {stage2_15[57]},
      {stage3_15[24]}
   );
   gpc1_1 gpc4798 (
      {stage2_15[58]},
      {stage3_15[25]}
   );
   gpc1_1 gpc4799 (
      {stage2_15[59]},
      {stage3_15[26]}
   );
   gpc1_1 gpc4800 (
      {stage2_15[60]},
      {stage3_15[27]}
   );
   gpc1_1 gpc4801 (
      {stage2_15[61]},
      {stage3_15[28]}
   );
   gpc1_1 gpc4802 (
      {stage2_15[62]},
      {stage3_15[29]}
   );
   gpc1_1 gpc4803 (
      {stage2_15[63]},
      {stage3_15[30]}
   );
   gpc1_1 gpc4804 (
      {stage2_15[64]},
      {stage3_15[31]}
   );
   gpc1_1 gpc4805 (
      {stage2_15[65]},
      {stage3_15[32]}
   );
   gpc1_1 gpc4806 (
      {stage2_15[66]},
      {stage3_15[33]}
   );
   gpc1_1 gpc4807 (
      {stage2_15[67]},
      {stage3_15[34]}
   );
   gpc1_1 gpc4808 (
      {stage2_15[68]},
      {stage3_15[35]}
   );
   gpc1_1 gpc4809 (
      {stage2_15[69]},
      {stage3_15[36]}
   );
   gpc1_1 gpc4810 (
      {stage2_15[70]},
      {stage3_15[37]}
   );
   gpc1_1 gpc4811 (
      {stage2_15[71]},
      {stage3_15[38]}
   );
   gpc1_1 gpc4812 (
      {stage2_15[72]},
      {stage3_15[39]}
   );
   gpc1_1 gpc4813 (
      {stage2_15[73]},
      {stage3_15[40]}
   );
   gpc1_1 gpc4814 (
      {stage2_16[53]},
      {stage3_16[18]}
   );
   gpc1_1 gpc4815 (
      {stage2_16[54]},
      {stage3_16[19]}
   );
   gpc1_1 gpc4816 (
      {stage2_17[48]},
      {stage3_17[21]}
   );
   gpc1_1 gpc4817 (
      {stage2_17[49]},
      {stage3_17[22]}
   );
   gpc1_1 gpc4818 (
      {stage2_17[50]},
      {stage3_17[23]}
   );
   gpc1_1 gpc4819 (
      {stage2_17[51]},
      {stage3_17[24]}
   );
   gpc1_1 gpc4820 (
      {stage2_17[52]},
      {stage3_17[25]}
   );
   gpc1_1 gpc4821 (
      {stage2_17[53]},
      {stage3_17[26]}
   );
   gpc1_1 gpc4822 (
      {stage2_17[54]},
      {stage3_17[27]}
   );
   gpc1_1 gpc4823 (
      {stage2_17[55]},
      {stage3_17[28]}
   );
   gpc1_1 gpc4824 (
      {stage2_17[56]},
      {stage3_17[29]}
   );
   gpc1_1 gpc4825 (
      {stage2_19[30]},
      {stage3_19[21]}
   );
   gpc1_1 gpc4826 (
      {stage2_19[31]},
      {stage3_19[22]}
   );
   gpc1_1 gpc4827 (
      {stage2_19[32]},
      {stage3_19[23]}
   );
   gpc1_1 gpc4828 (
      {stage2_19[33]},
      {stage3_19[24]}
   );
   gpc1_1 gpc4829 (
      {stage2_19[34]},
      {stage3_19[25]}
   );
   gpc1_1 gpc4830 (
      {stage2_19[35]},
      {stage3_19[26]}
   );
   gpc1_1 gpc4831 (
      {stage2_19[36]},
      {stage3_19[27]}
   );
   gpc1_1 gpc4832 (
      {stage2_20[72]},
      {stage3_20[16]}
   );
   gpc1_1 gpc4833 (
      {stage2_20[73]},
      {stage3_20[17]}
   );
   gpc1_1 gpc4834 (
      {stage2_20[74]},
      {stage3_20[18]}
   );
   gpc1_1 gpc4835 (
      {stage2_20[75]},
      {stage3_20[19]}
   );
   gpc1_1 gpc4836 (
      {stage2_20[76]},
      {stage3_20[20]}
   );
   gpc1_1 gpc4837 (
      {stage2_20[77]},
      {stage3_20[21]}
   );
   gpc1_1 gpc4838 (
      {stage2_20[78]},
      {stage3_20[22]}
   );
   gpc1_1 gpc4839 (
      {stage2_20[79]},
      {stage3_20[23]}
   );
   gpc1_1 gpc4840 (
      {stage2_22[40]},
      {stage3_22[28]}
   );
   gpc1_1 gpc4841 (
      {stage2_24[72]},
      {stage3_24[21]}
   );
   gpc1_1 gpc4842 (
      {stage2_24[73]},
      {stage3_24[22]}
   );
   gpc1_1 gpc4843 (
      {stage2_24[74]},
      {stage3_24[23]}
   );
   gpc1_1 gpc4844 (
      {stage2_24[75]},
      {stage3_24[24]}
   );
   gpc1_1 gpc4845 (
      {stage2_24[76]},
      {stage3_24[25]}
   );
   gpc1_1 gpc4846 (
      {stage2_24[77]},
      {stage3_24[26]}
   );
   gpc1_1 gpc4847 (
      {stage2_24[78]},
      {stage3_24[27]}
   );
   gpc1_1 gpc4848 (
      {stage2_24[79]},
      {stage3_24[28]}
   );
   gpc1_1 gpc4849 (
      {stage2_24[80]},
      {stage3_24[29]}
   );
   gpc1_1 gpc4850 (
      {stage2_24[81]},
      {stage3_24[30]}
   );
   gpc1_1 gpc4851 (
      {stage2_25[46]},
      {stage3_25[29]}
   );
   gpc1_1 gpc4852 (
      {stage2_25[47]},
      {stage3_25[30]}
   );
   gpc1_1 gpc4853 (
      {stage2_25[48]},
      {stage3_25[31]}
   );
   gpc1_1 gpc4854 (
      {stage2_25[49]},
      {stage3_25[32]}
   );
   gpc1_1 gpc4855 (
      {stage2_25[50]},
      {stage3_25[33]}
   );
   gpc1_1 gpc4856 (
      {stage2_29[36]},
      {stage3_29[25]}
   );
   gpc1_1 gpc4857 (
      {stage2_29[37]},
      {stage3_29[26]}
   );
   gpc1_1 gpc4858 (
      {stage2_29[38]},
      {stage3_29[27]}
   );
   gpc1_1 gpc4859 (
      {stage2_29[39]},
      {stage3_29[28]}
   );
   gpc1_1 gpc4860 (
      {stage2_29[40]},
      {stage3_29[29]}
   );
   gpc1_1 gpc4861 (
      {stage2_29[41]},
      {stage3_29[30]}
   );
   gpc1_1 gpc4862 (
      {stage2_29[42]},
      {stage3_29[31]}
   );
   gpc1_1 gpc4863 (
      {stage2_29[43]},
      {stage3_29[32]}
   );
   gpc1_1 gpc4864 (
      {stage2_29[44]},
      {stage3_29[33]}
   );
   gpc1_1 gpc4865 (
      {stage2_29[45]},
      {stage3_29[34]}
   );
   gpc1_1 gpc4866 (
      {stage2_30[52]},
      {stage3_30[19]}
   );
   gpc1_1 gpc4867 (
      {stage2_30[53]},
      {stage3_30[20]}
   );
   gpc1_1 gpc4868 (
      {stage2_30[54]},
      {stage3_30[21]}
   );
   gpc1_1 gpc4869 (
      {stage2_30[55]},
      {stage3_30[22]}
   );
   gpc1_1 gpc4870 (
      {stage2_30[56]},
      {stage3_30[23]}
   );
   gpc1_1 gpc4871 (
      {stage2_30[57]},
      {stage3_30[24]}
   );
   gpc1_1 gpc4872 (
      {stage2_30[58]},
      {stage3_30[25]}
   );
   gpc1_1 gpc4873 (
      {stage2_31[43]},
      {stage3_31[21]}
   );
   gpc1_1 gpc4874 (
      {stage2_31[44]},
      {stage3_31[22]}
   );
   gpc1_1 gpc4875 (
      {stage2_31[45]},
      {stage3_31[23]}
   );
   gpc1_1 gpc4876 (
      {stage2_31[46]},
      {stage3_31[24]}
   );
   gpc1_1 gpc4877 (
      {stage2_31[47]},
      {stage3_31[25]}
   );
   gpc1_1 gpc4878 (
      {stage2_31[48]},
      {stage3_31[26]}
   );
   gpc1_1 gpc4879 (
      {stage2_31[49]},
      {stage3_31[27]}
   );
   gpc1_1 gpc4880 (
      {stage2_31[50]},
      {stage3_31[28]}
   );
   gpc1_1 gpc4881 (
      {stage2_31[51]},
      {stage3_31[29]}
   );
   gpc1_1 gpc4882 (
      {stage2_31[52]},
      {stage3_31[30]}
   );
   gpc1_1 gpc4883 (
      {stage2_31[53]},
      {stage3_31[31]}
   );
   gpc1_1 gpc4884 (
      {stage2_32[39]},
      {stage3_32[20]}
   );
   gpc1_1 gpc4885 (
      {stage2_32[40]},
      {stage3_32[21]}
   );
   gpc1_1 gpc4886 (
      {stage2_32[41]},
      {stage3_32[22]}
   );
   gpc1_1 gpc4887 (
      {stage2_32[42]},
      {stage3_32[23]}
   );
   gpc1_1 gpc4888 (
      {stage2_32[43]},
      {stage3_32[24]}
   );
   gpc1_1 gpc4889 (
      {stage2_32[44]},
      {stage3_32[25]}
   );
   gpc1_1 gpc4890 (
      {stage2_32[45]},
      {stage3_32[26]}
   );
   gpc1_1 gpc4891 (
      {stage2_32[46]},
      {stage3_32[27]}
   );
   gpc1_1 gpc4892 (
      {stage2_33[38]},
      {stage3_33[13]}
   );
   gpc1_1 gpc4893 (
      {stage2_33[39]},
      {stage3_33[14]}
   );
   gpc1_1 gpc4894 (
      {stage2_33[40]},
      {stage3_33[15]}
   );
   gpc1_1 gpc4895 (
      {stage2_33[41]},
      {stage3_33[16]}
   );
   gpc1_1 gpc4896 (
      {stage2_33[42]},
      {stage3_33[17]}
   );
   gpc1_1 gpc4897 (
      {stage2_33[43]},
      {stage3_33[18]}
   );
   gpc1_1 gpc4898 (
      {stage2_33[44]},
      {stage3_33[19]}
   );
   gpc1_1 gpc4899 (
      {stage2_33[45]},
      {stage3_33[20]}
   );
   gpc1_1 gpc4900 (
      {stage2_33[46]},
      {stage3_33[21]}
   );
   gpc1_1 gpc4901 (
      {stage2_33[47]},
      {stage3_33[22]}
   );
   gpc1_1 gpc4902 (
      {stage2_33[48]},
      {stage3_33[23]}
   );
   gpc1_1 gpc4903 (
      {stage2_33[49]},
      {stage3_33[24]}
   );
   gpc1_1 gpc4904 (
      {stage2_33[50]},
      {stage3_33[25]}
   );
   gpc1_1 gpc4905 (
      {stage2_33[51]},
      {stage3_33[26]}
   );
   gpc1_1 gpc4906 (
      {stage2_34[24]},
      {stage3_34[14]}
   );
   gpc1_1 gpc4907 (
      {stage2_34[25]},
      {stage3_34[15]}
   );
   gpc1_1 gpc4908 (
      {stage2_34[26]},
      {stage3_34[16]}
   );
   gpc1_1 gpc4909 (
      {stage2_34[27]},
      {stage3_34[17]}
   );
   gpc1_1 gpc4910 (
      {stage2_34[28]},
      {stage3_34[18]}
   );
   gpc1_1 gpc4911 (
      {stage2_34[29]},
      {stage3_34[19]}
   );
   gpc1_1 gpc4912 (
      {stage2_34[30]},
      {stage3_34[20]}
   );
   gpc1_1 gpc4913 (
      {stage2_34[31]},
      {stage3_34[21]}
   );
   gpc1_1 gpc4914 (
      {stage2_34[32]},
      {stage3_34[22]}
   );
   gpc1_1 gpc4915 (
      {stage2_34[33]},
      {stage3_34[23]}
   );
   gpc1_1 gpc4916 (
      {stage2_34[34]},
      {stage3_34[24]}
   );
   gpc1_1 gpc4917 (
      {stage2_34[35]},
      {stage3_34[25]}
   );
   gpc1_1 gpc4918 (
      {stage2_34[36]},
      {stage3_34[26]}
   );
   gpc1_1 gpc4919 (
      {stage2_35[47]},
      {stage3_35[21]}
   );
   gpc1_1 gpc4920 (
      {stage2_35[48]},
      {stage3_35[22]}
   );
   gpc1_1 gpc4921 (
      {stage2_35[49]},
      {stage3_35[23]}
   );
   gpc1_1 gpc4922 (
      {stage2_35[50]},
      {stage3_35[24]}
   );
   gpc1_1 gpc4923 (
      {stage2_35[51]},
      {stage3_35[25]}
   );
   gpc1_1 gpc4924 (
      {stage2_35[52]},
      {stage3_35[26]}
   );
   gpc1_1 gpc4925 (
      {stage2_35[53]},
      {stage3_35[27]}
   );
   gpc1_1 gpc4926 (
      {stage2_35[54]},
      {stage3_35[28]}
   );
   gpc1_1 gpc4927 (
      {stage2_35[55]},
      {stage3_35[29]}
   );
   gpc1_1 gpc4928 (
      {stage2_35[56]},
      {stage3_35[30]}
   );
   gpc1_1 gpc4929 (
      {stage2_35[57]},
      {stage3_35[31]}
   );
   gpc1_1 gpc4930 (
      {stage2_35[58]},
      {stage3_35[32]}
   );
   gpc1_1 gpc4931 (
      {stage2_37[54]},
      {stage3_37[18]}
   );
   gpc1_1 gpc4932 (
      {stage2_38[42]},
      {stage3_38[18]}
   );
   gpc1_1 gpc4933 (
      {stage2_38[43]},
      {stage3_38[19]}
   );
   gpc1_1 gpc4934 (
      {stage2_38[44]},
      {stage3_38[20]}
   );
   gpc1_1 gpc4935 (
      {stage2_38[45]},
      {stage3_38[21]}
   );
   gpc1_1 gpc4936 (
      {stage2_38[46]},
      {stage3_38[22]}
   );
   gpc1_1 gpc4937 (
      {stage2_40[39]},
      {stage3_40[24]}
   );
   gpc1_1 gpc4938 (
      {stage2_40[40]},
      {stage3_40[25]}
   );
   gpc1_1 gpc4939 (
      {stage2_40[41]},
      {stage3_40[26]}
   );
   gpc1_1 gpc4940 (
      {stage2_40[42]},
      {stage3_40[27]}
   );
   gpc1_1 gpc4941 (
      {stage2_40[43]},
      {stage3_40[28]}
   );
   gpc1_1 gpc4942 (
      {stage2_40[44]},
      {stage3_40[29]}
   );
   gpc1_1 gpc4943 (
      {stage2_42[58]},
      {stage3_42[25]}
   );
   gpc1_1 gpc4944 (
      {stage2_42[59]},
      {stage3_42[26]}
   );
   gpc1_1 gpc4945 (
      {stage2_42[60]},
      {stage3_42[27]}
   );
   gpc1_1 gpc4946 (
      {stage2_42[61]},
      {stage3_42[28]}
   );
   gpc1_1 gpc4947 (
      {stage2_42[62]},
      {stage3_42[29]}
   );
   gpc1_1 gpc4948 (
      {stage2_43[54]},
      {stage3_43[31]}
   );
   gpc1_1 gpc4949 (
      {stage2_43[55]},
      {stage3_43[32]}
   );
   gpc1_1 gpc4950 (
      {stage2_43[56]},
      {stage3_43[33]}
   );
   gpc1_1 gpc4951 (
      {stage2_43[57]},
      {stage3_43[34]}
   );
   gpc1_1 gpc4952 (
      {stage2_43[58]},
      {stage3_43[35]}
   );
   gpc1_1 gpc4953 (
      {stage2_43[59]},
      {stage3_43[36]}
   );
   gpc1_1 gpc4954 (
      {stage2_43[60]},
      {stage3_43[37]}
   );
   gpc1_1 gpc4955 (
      {stage2_43[61]},
      {stage3_43[38]}
   );
   gpc1_1 gpc4956 (
      {stage2_45[66]},
      {stage3_45[26]}
   );
   gpc1_1 gpc4957 (
      {stage2_45[67]},
      {stage3_45[27]}
   );
   gpc1_1 gpc4958 (
      {stage2_45[68]},
      {stage3_45[28]}
   );
   gpc1_1 gpc4959 (
      {stage2_45[69]},
      {stage3_45[29]}
   );
   gpc1_1 gpc4960 (
      {stage2_45[70]},
      {stage3_45[30]}
   );
   gpc1_1 gpc4961 (
      {stage2_45[71]},
      {stage3_45[31]}
   );
   gpc1_1 gpc4962 (
      {stage2_45[72]},
      {stage3_45[32]}
   );
   gpc1_1 gpc4963 (
      {stage2_45[73]},
      {stage3_45[33]}
   );
   gpc1_1 gpc4964 (
      {stage2_45[74]},
      {stage3_45[34]}
   );
   gpc1_1 gpc4965 (
      {stage2_45[75]},
      {stage3_45[35]}
   );
   gpc1_1 gpc4966 (
      {stage2_45[76]},
      {stage3_45[36]}
   );
   gpc1_1 gpc4967 (
      {stage2_45[77]},
      {stage3_45[37]}
   );
   gpc1_1 gpc4968 (
      {stage2_45[78]},
      {stage3_45[38]}
   );
   gpc1_1 gpc4969 (
      {stage2_46[42]},
      {stage3_46[19]}
   );
   gpc1_1 gpc4970 (
      {stage2_46[43]},
      {stage3_46[20]}
   );
   gpc1_1 gpc4971 (
      {stage2_46[44]},
      {stage3_46[21]}
   );
   gpc1_1 gpc4972 (
      {stage2_46[45]},
      {stage3_46[22]}
   );
   gpc1_1 gpc4973 (
      {stage2_46[46]},
      {stage3_46[23]}
   );
   gpc1_1 gpc4974 (
      {stage2_46[47]},
      {stage3_46[24]}
   );
   gpc1_1 gpc4975 (
      {stage2_46[48]},
      {stage3_46[25]}
   );
   gpc1_1 gpc4976 (
      {stage2_46[49]},
      {stage3_46[26]}
   );
   gpc1_1 gpc4977 (
      {stage2_46[50]},
      {stage3_46[27]}
   );
   gpc1_1 gpc4978 (
      {stage2_46[51]},
      {stage3_46[28]}
   );
   gpc1_1 gpc4979 (
      {stage2_46[52]},
      {stage3_46[29]}
   );
   gpc1_1 gpc4980 (
      {stage2_46[53]},
      {stage3_46[30]}
   );
   gpc1_1 gpc4981 (
      {stage2_46[54]},
      {stage3_46[31]}
   );
   gpc1_1 gpc4982 (
      {stage2_46[55]},
      {stage3_46[32]}
   );
   gpc1_1 gpc4983 (
      {stage2_46[56]},
      {stage3_46[33]}
   );
   gpc1_1 gpc4984 (
      {stage2_46[57]},
      {stage3_46[34]}
   );
   gpc1_1 gpc4985 (
      {stage2_46[58]},
      {stage3_46[35]}
   );
   gpc1_1 gpc4986 (
      {stage2_46[59]},
      {stage3_46[36]}
   );
   gpc1_1 gpc4987 (
      {stage2_46[60]},
      {stage3_46[37]}
   );
   gpc1_1 gpc4988 (
      {stage2_46[61]},
      {stage3_46[38]}
   );
   gpc1_1 gpc4989 (
      {stage2_46[62]},
      {stage3_46[39]}
   );
   gpc1_1 gpc4990 (
      {stage2_47[61]},
      {stage3_47[23]}
   );
   gpc1_1 gpc4991 (
      {stage2_47[62]},
      {stage3_47[24]}
   );
   gpc1_1 gpc4992 (
      {stage2_47[63]},
      {stage3_47[25]}
   );
   gpc1_1 gpc4993 (
      {stage2_47[64]},
      {stage3_47[26]}
   );
   gpc1_1 gpc4994 (
      {stage2_47[65]},
      {stage3_47[27]}
   );
   gpc1_1 gpc4995 (
      {stage2_47[66]},
      {stage3_47[28]}
   );
   gpc1_1 gpc4996 (
      {stage2_47[67]},
      {stage3_47[29]}
   );
   gpc1_1 gpc4997 (
      {stage2_47[68]},
      {stage3_47[30]}
   );
   gpc1_1 gpc4998 (
      {stage2_47[69]},
      {stage3_47[31]}
   );
   gpc1_1 gpc4999 (
      {stage2_47[70]},
      {stage3_47[32]}
   );
   gpc1_1 gpc5000 (
      {stage2_49[70]},
      {stage3_49[23]}
   );
   gpc1_1 gpc5001 (
      {stage2_49[71]},
      {stage3_49[24]}
   );
   gpc1_1 gpc5002 (
      {stage2_49[72]},
      {stage3_49[25]}
   );
   gpc1_1 gpc5003 (
      {stage2_49[73]},
      {stage3_49[26]}
   );
   gpc1_1 gpc5004 (
      {stage2_49[74]},
      {stage3_49[27]}
   );
   gpc1_1 gpc5005 (
      {stage2_49[75]},
      {stage3_49[28]}
   );
   gpc1_1 gpc5006 (
      {stage2_49[76]},
      {stage3_49[29]}
   );
   gpc1_1 gpc5007 (
      {stage2_49[77]},
      {stage3_49[30]}
   );
   gpc1_1 gpc5008 (
      {stage2_49[78]},
      {stage3_49[31]}
   );
   gpc1_1 gpc5009 (
      {stage2_49[79]},
      {stage3_49[32]}
   );
   gpc1_1 gpc5010 (
      {stage2_49[80]},
      {stage3_49[33]}
   );
   gpc1_1 gpc5011 (
      {stage2_49[81]},
      {stage3_49[34]}
   );
   gpc1_1 gpc5012 (
      {stage2_49[82]},
      {stage3_49[35]}
   );
   gpc1_1 gpc5013 (
      {stage2_49[83]},
      {stage3_49[36]}
   );
   gpc1_1 gpc5014 (
      {stage2_49[84]},
      {stage3_49[37]}
   );
   gpc1_1 gpc5015 (
      {stage2_49[85]},
      {stage3_49[38]}
   );
   gpc1_1 gpc5016 (
      {stage2_49[86]},
      {stage3_49[39]}
   );
   gpc1_1 gpc5017 (
      {stage2_49[87]},
      {stage3_49[40]}
   );
   gpc1_1 gpc5018 (
      {stage2_49[88]},
      {stage3_49[41]}
   );
   gpc1_1 gpc5019 (
      {stage2_49[89]},
      {stage3_49[42]}
   );
   gpc1_1 gpc5020 (
      {stage2_49[90]},
      {stage3_49[43]}
   );
   gpc1_1 gpc5021 (
      {stage2_49[91]},
      {stage3_49[44]}
   );
   gpc1_1 gpc5022 (
      {stage2_49[92]},
      {stage3_49[45]}
   );
   gpc1_1 gpc5023 (
      {stage2_49[93]},
      {stage3_49[46]}
   );
   gpc1_1 gpc5024 (
      {stage2_49[94]},
      {stage3_49[47]}
   );
   gpc1_1 gpc5025 (
      {stage2_49[95]},
      {stage3_49[48]}
   );
   gpc1_1 gpc5026 (
      {stage2_49[96]},
      {stage3_49[49]}
   );
   gpc1_1 gpc5027 (
      {stage2_49[97]},
      {stage3_49[50]}
   );
   gpc1_1 gpc5028 (
      {stage2_49[98]},
      {stage3_49[51]}
   );
   gpc1_1 gpc5029 (
      {stage2_49[99]},
      {stage3_49[52]}
   );
   gpc1_1 gpc5030 (
      {stage2_49[100]},
      {stage3_49[53]}
   );
   gpc1_1 gpc5031 (
      {stage2_49[101]},
      {stage3_49[54]}
   );
   gpc1_1 gpc5032 (
      {stage2_49[102]},
      {stage3_49[55]}
   );
   gpc1_1 gpc5033 (
      {stage2_49[103]},
      {stage3_49[56]}
   );
   gpc1_1 gpc5034 (
      {stage2_49[104]},
      {stage3_49[57]}
   );
   gpc1_1 gpc5035 (
      {stage2_49[105]},
      {stage3_49[58]}
   );
   gpc1_1 gpc5036 (
      {stage2_49[106]},
      {stage3_49[59]}
   );
   gpc1_1 gpc5037 (
      {stage2_49[107]},
      {stage3_49[60]}
   );
   gpc1_1 gpc5038 (
      {stage2_49[108]},
      {stage3_49[61]}
   );
   gpc1_1 gpc5039 (
      {stage2_49[109]},
      {stage3_49[62]}
   );
   gpc1_1 gpc5040 (
      {stage2_49[110]},
      {stage3_49[63]}
   );
   gpc1_1 gpc5041 (
      {stage2_49[111]},
      {stage3_49[64]}
   );
   gpc1_1 gpc5042 (
      {stage2_49[112]},
      {stage3_49[65]}
   );
   gpc1_1 gpc5043 (
      {stage2_49[113]},
      {stage3_49[66]}
   );
   gpc1_1 gpc5044 (
      {stage2_49[114]},
      {stage3_49[67]}
   );
   gpc1_1 gpc5045 (
      {stage2_50[57]},
      {stage3_50[19]}
   );
   gpc1_1 gpc5046 (
      {stage2_50[58]},
      {stage3_50[20]}
   );
   gpc1_1 gpc5047 (
      {stage2_50[59]},
      {stage3_50[21]}
   );
   gpc1_1 gpc5048 (
      {stage2_50[60]},
      {stage3_50[22]}
   );
   gpc1_1 gpc5049 (
      {stage2_50[61]},
      {stage3_50[23]}
   );
   gpc1_1 gpc5050 (
      {stage2_50[62]},
      {stage3_50[24]}
   );
   gpc1_1 gpc5051 (
      {stage2_50[63]},
      {stage3_50[25]}
   );
   gpc1_1 gpc5052 (
      {stage2_50[64]},
      {stage3_50[26]}
   );
   gpc1_1 gpc5053 (
      {stage2_50[65]},
      {stage3_50[27]}
   );
   gpc1_1 gpc5054 (
      {stage2_50[66]},
      {stage3_50[28]}
   );
   gpc1_1 gpc5055 (
      {stage2_50[67]},
      {stage3_50[29]}
   );
   gpc1_1 gpc5056 (
      {stage2_51[61]},
      {stage3_51[30]}
   );
   gpc1_1 gpc5057 (
      {stage2_51[62]},
      {stage3_51[31]}
   );
   gpc1_1 gpc5058 (
      {stage2_51[63]},
      {stage3_51[32]}
   );
   gpc1_1 gpc5059 (
      {stage2_51[64]},
      {stage3_51[33]}
   );
   gpc1_1 gpc5060 (
      {stage2_51[65]},
      {stage3_51[34]}
   );
   gpc1_1 gpc5061 (
      {stage2_51[66]},
      {stage3_51[35]}
   );
   gpc1_1 gpc5062 (
      {stage2_51[67]},
      {stage3_51[36]}
   );
   gpc1_1 gpc5063 (
      {stage2_51[68]},
      {stage3_51[37]}
   );
   gpc1_1 gpc5064 (
      {stage2_51[69]},
      {stage3_51[38]}
   );
   gpc1_1 gpc5065 (
      {stage2_51[70]},
      {stage3_51[39]}
   );
   gpc1_1 gpc5066 (
      {stage2_51[71]},
      {stage3_51[40]}
   );
   gpc1_1 gpc5067 (
      {stage2_51[72]},
      {stage3_51[41]}
   );
   gpc1_1 gpc5068 (
      {stage2_51[73]},
      {stage3_51[42]}
   );
   gpc1_1 gpc5069 (
      {stage2_51[74]},
      {stage3_51[43]}
   );
   gpc1_1 gpc5070 (
      {stage2_51[75]},
      {stage3_51[44]}
   );
   gpc1_1 gpc5071 (
      {stage2_51[76]},
      {stage3_51[45]}
   );
   gpc1_1 gpc5072 (
      {stage2_51[77]},
      {stage3_51[46]}
   );
   gpc1_1 gpc5073 (
      {stage2_51[78]},
      {stage3_51[47]}
   );
   gpc1_1 gpc5074 (
      {stage2_52[39]},
      {stage3_52[28]}
   );
   gpc1_1 gpc5075 (
      {stage2_52[40]},
      {stage3_52[29]}
   );
   gpc1_1 gpc5076 (
      {stage2_52[41]},
      {stage3_52[30]}
   );
   gpc1_1 gpc5077 (
      {stage2_52[42]},
      {stage3_52[31]}
   );
   gpc1_1 gpc5078 (
      {stage2_52[43]},
      {stage3_52[32]}
   );
   gpc1_1 gpc5079 (
      {stage2_52[44]},
      {stage3_52[33]}
   );
   gpc1_1 gpc5080 (
      {stage2_52[45]},
      {stage3_52[34]}
   );
   gpc1_1 gpc5081 (
      {stage2_52[46]},
      {stage3_52[35]}
   );
   gpc1_1 gpc5082 (
      {stage2_52[47]},
      {stage3_52[36]}
   );
   gpc1_1 gpc5083 (
      {stage2_52[48]},
      {stage3_52[37]}
   );
   gpc1_1 gpc5084 (
      {stage2_52[49]},
      {stage3_52[38]}
   );
   gpc1_1 gpc5085 (
      {stage2_52[50]},
      {stage3_52[39]}
   );
   gpc1_1 gpc5086 (
      {stage2_53[66]},
      {stage3_53[16]}
   );
   gpc1_1 gpc5087 (
      {stage2_53[67]},
      {stage3_53[17]}
   );
   gpc1_1 gpc5088 (
      {stage2_53[68]},
      {stage3_53[18]}
   );
   gpc1_1 gpc5089 (
      {stage2_53[69]},
      {stage3_53[19]}
   );
   gpc1_1 gpc5090 (
      {stage2_53[70]},
      {stage3_53[20]}
   );
   gpc1_1 gpc5091 (
      {stage2_53[71]},
      {stage3_53[21]}
   );
   gpc1_1 gpc5092 (
      {stage2_53[72]},
      {stage3_53[22]}
   );
   gpc1_1 gpc5093 (
      {stage2_53[73]},
      {stage3_53[23]}
   );
   gpc1_1 gpc5094 (
      {stage2_53[74]},
      {stage3_53[24]}
   );
   gpc1_1 gpc5095 (
      {stage2_53[75]},
      {stage3_53[25]}
   );
   gpc1_1 gpc5096 (
      {stage2_53[76]},
      {stage3_53[26]}
   );
   gpc1_1 gpc5097 (
      {stage2_53[77]},
      {stage3_53[27]}
   );
   gpc1_1 gpc5098 (
      {stage2_54[72]},
      {stage3_54[25]}
   );
   gpc1_1 gpc5099 (
      {stage2_54[73]},
      {stage3_54[26]}
   );
   gpc1_1 gpc5100 (
      {stage2_54[74]},
      {stage3_54[27]}
   );
   gpc1_1 gpc5101 (
      {stage2_56[67]},
      {stage3_56[20]}
   );
   gpc1_1 gpc5102 (
      {stage2_56[68]},
      {stage3_56[21]}
   );
   gpc1_1 gpc5103 (
      {stage2_56[69]},
      {stage3_56[22]}
   );
   gpc1_1 gpc5104 (
      {stage2_56[70]},
      {stage3_56[23]}
   );
   gpc1_1 gpc5105 (
      {stage2_56[71]},
      {stage3_56[24]}
   );
   gpc1_1 gpc5106 (
      {stage2_56[72]},
      {stage3_56[25]}
   );
   gpc1_1 gpc5107 (
      {stage2_57[72]},
      {stage3_57[22]}
   );
   gpc1_1 gpc5108 (
      {stage2_57[73]},
      {stage3_57[23]}
   );
   gpc1_1 gpc5109 (
      {stage2_57[74]},
      {stage3_57[24]}
   );
   gpc1_1 gpc5110 (
      {stage2_57[75]},
      {stage3_57[25]}
   );
   gpc1_1 gpc5111 (
      {stage2_57[76]},
      {stage3_57[26]}
   );
   gpc1_1 gpc5112 (
      {stage2_57[77]},
      {stage3_57[27]}
   );
   gpc1_1 gpc5113 (
      {stage2_57[78]},
      {stage3_57[28]}
   );
   gpc1_1 gpc5114 (
      {stage2_57[79]},
      {stage3_57[29]}
   );
   gpc1_1 gpc5115 (
      {stage2_57[80]},
      {stage3_57[30]}
   );
   gpc1_1 gpc5116 (
      {stage2_57[81]},
      {stage3_57[31]}
   );
   gpc1_1 gpc5117 (
      {stage2_57[82]},
      {stage3_57[32]}
   );
   gpc1_1 gpc5118 (
      {stage2_59[36]},
      {stage3_59[21]}
   );
   gpc1_1 gpc5119 (
      {stage2_59[37]},
      {stage3_59[22]}
   );
   gpc1_1 gpc5120 (
      {stage2_59[38]},
      {stage3_59[23]}
   );
   gpc1_1 gpc5121 (
      {stage2_59[39]},
      {stage3_59[24]}
   );
   gpc1_1 gpc5122 (
      {stage2_59[40]},
      {stage3_59[25]}
   );
   gpc1_1 gpc5123 (
      {stage2_59[41]},
      {stage3_59[26]}
   );
   gpc1_1 gpc5124 (
      {stage2_59[42]},
      {stage3_59[27]}
   );
   gpc1_1 gpc5125 (
      {stage2_59[43]},
      {stage3_59[28]}
   );
   gpc1_1 gpc5126 (
      {stage2_59[44]},
      {stage3_59[29]}
   );
   gpc1_1 gpc5127 (
      {stage2_59[45]},
      {stage3_59[30]}
   );
   gpc1_1 gpc5128 (
      {stage2_59[46]},
      {stage3_59[31]}
   );
   gpc1_1 gpc5129 (
      {stage2_59[47]},
      {stage3_59[32]}
   );
   gpc1_1 gpc5130 (
      {stage2_60[42]},
      {stage3_60[14]}
   );
   gpc1_1 gpc5131 (
      {stage2_60[43]},
      {stage3_60[15]}
   );
   gpc1_1 gpc5132 (
      {stage2_60[44]},
      {stage3_60[16]}
   );
   gpc1_1 gpc5133 (
      {stage2_60[45]},
      {stage3_60[17]}
   );
   gpc1_1 gpc5134 (
      {stage2_60[46]},
      {stage3_60[18]}
   );
   gpc1_1 gpc5135 (
      {stage2_60[47]},
      {stage3_60[19]}
   );
   gpc1_1 gpc5136 (
      {stage2_60[48]},
      {stage3_60[20]}
   );
   gpc1_1 gpc5137 (
      {stage2_60[49]},
      {stage3_60[21]}
   );
   gpc1_1 gpc5138 (
      {stage2_60[50]},
      {stage3_60[22]}
   );
   gpc1_1 gpc5139 (
      {stage2_60[51]},
      {stage3_60[23]}
   );
   gpc1_1 gpc5140 (
      {stage2_60[52]},
      {stage3_60[24]}
   );
   gpc1_1 gpc5141 (
      {stage2_60[53]},
      {stage3_60[25]}
   );
   gpc1_1 gpc5142 (
      {stage2_60[54]},
      {stage3_60[26]}
   );
   gpc1_1 gpc5143 (
      {stage2_60[55]},
      {stage3_60[27]}
   );
   gpc1_1 gpc5144 (
      {stage2_60[56]},
      {stage3_60[28]}
   );
   gpc1_1 gpc5145 (
      {stage2_60[57]},
      {stage3_60[29]}
   );
   gpc1_1 gpc5146 (
      {stage2_60[58]},
      {stage3_60[30]}
   );
   gpc1_1 gpc5147 (
      {stage2_60[59]},
      {stage3_60[31]}
   );
   gpc1_1 gpc5148 (
      {stage2_60[60]},
      {stage3_60[32]}
   );
   gpc1_1 gpc5149 (
      {stage2_60[61]},
      {stage3_60[33]}
   );
   gpc1_1 gpc5150 (
      {stage2_60[62]},
      {stage3_60[34]}
   );
   gpc1_1 gpc5151 (
      {stage2_61[54]},
      {stage3_61[21]}
   );
   gpc1_1 gpc5152 (
      {stage2_61[55]},
      {stage3_61[22]}
   );
   gpc1_1 gpc5153 (
      {stage2_61[56]},
      {stage3_61[23]}
   );
   gpc1_1 gpc5154 (
      {stage2_62[51]},
      {stage3_62[26]}
   );
   gpc1_1 gpc5155 (
      {stage2_62[52]},
      {stage3_62[27]}
   );
   gpc1_1 gpc5156 (
      {stage2_63[66]},
      {stage3_63[19]}
   );
   gpc1_1 gpc5157 (
      {stage2_63[67]},
      {stage3_63[20]}
   );
   gpc1_1 gpc5158 (
      {stage2_63[68]},
      {stage3_63[21]}
   );
   gpc1_1 gpc5159 (
      {stage2_63[69]},
      {stage3_63[22]}
   );
   gpc1_1 gpc5160 (
      {stage2_63[70]},
      {stage3_63[23]}
   );
   gpc1_1 gpc5161 (
      {stage2_63[71]},
      {stage3_63[24]}
   );
   gpc1_1 gpc5162 (
      {stage2_63[72]},
      {stage3_63[25]}
   );
   gpc1_1 gpc5163 (
      {stage2_63[73]},
      {stage3_63[26]}
   );
   gpc1_1 gpc5164 (
      {stage2_63[74]},
      {stage3_63[27]}
   );
   gpc1_1 gpc5165 (
      {stage2_65[9]},
      {stage3_65[19]}
   );
   gpc1_1 gpc5166 (
      {stage2_65[10]},
      {stage3_65[20]}
   );
   gpc1_1 gpc5167 (
      {stage2_65[11]},
      {stage3_65[21]}
   );
   gpc1_1 gpc5168 (
      {stage2_65[12]},
      {stage3_65[22]}
   );
   gpc1_1 gpc5169 (
      {stage2_65[13]},
      {stage3_65[23]}
   );
   gpc1_1 gpc5170 (
      {stage2_65[14]},
      {stage3_65[24]}
   );
   gpc1_1 gpc5171 (
      {stage2_65[15]},
      {stage3_65[25]}
   );
   gpc1_1 gpc5172 (
      {stage2_65[16]},
      {stage3_65[26]}
   );
   gpc1_1 gpc5173 (
      {stage2_65[17]},
      {stage3_65[27]}
   );
   gpc1_1 gpc5174 (
      {stage2_66[0]},
      {stage3_66[11]}
   );
   gpc1_1 gpc5175 (
      {stage2_66[1]},
      {stage3_66[12]}
   );
   gpc1_1 gpc5176 (
      {stage2_66[2]},
      {stage3_66[13]}
   );
   gpc1_1 gpc5177 (
      {stage2_66[3]},
      {stage3_66[14]}
   );
   gpc1_1 gpc5178 (
      {stage2_66[4]},
      {stage3_66[15]}
   );
   gpc1_1 gpc5179 (
      {stage2_66[5]},
      {stage3_66[16]}
   );
   gpc1_1 gpc5180 (
      {stage2_66[6]},
      {stage3_66[17]}
   );
   gpc1_1 gpc5181 (
      {stage2_66[7]},
      {stage3_66[18]}
   );
   gpc1_1 gpc5182 (
      {stage2_66[8]},
      {stage3_66[19]}
   );
   gpc1_1 gpc5183 (
      {stage2_66[9]},
      {stage3_66[20]}
   );
   gpc1_1 gpc5184 (
      {stage2_66[10]},
      {stage3_66[21]}
   );
   gpc1_1 gpc5185 (
      {stage2_66[11]},
      {stage3_66[22]}
   );
   gpc1_1 gpc5186 (
      {stage2_66[12]},
      {stage3_66[23]}
   );
   gpc1_1 gpc5187 (
      {stage2_66[13]},
      {stage3_66[24]}
   );
   gpc1_1 gpc5188 (
      {stage2_66[14]},
      {stage3_66[25]}
   );
   gpc1_1 gpc5189 (
      {stage2_66[15]},
      {stage3_66[26]}
   );
   gpc1_1 gpc5190 (
      {stage2_66[16]},
      {stage3_66[27]}
   );
   gpc1_1 gpc5191 (
      {stage2_67[6]},
      {stage3_67[1]}
   );
   gpc2135_5 gpc5192 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4]},
      {stage3_2[0], stage3_2[1], stage3_2[2]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc1163_5 gpc5193 (
      {stage3_1[5], stage3_1[6], stage3_1[7]},
      {stage3_2[3], stage3_2[4], stage3_2[5], stage3_2[6], stage3_2[7], stage3_2[8]},
      {stage3_3[1]},
      {stage3_4[2]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc5194 (
      {stage3_2[9], stage3_2[10], stage3_2[11], stage3_2[12], stage3_2[13]},
      {stage3_3[2]},
      {stage3_4[3], stage3_4[4], stage3_4[5], stage3_4[6], stage3_4[7], stage3_4[8]},
      {stage4_6[0],stage4_5[2],stage4_4[2],stage4_3[2],stage4_2[2]}
   );
   gpc606_5 gpc5195 (
      {stage3_4[9], stage3_4[10], stage3_4[11], stage3_4[12], stage3_4[13], stage3_4[14]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[3],stage4_4[3]}
   );
   gpc1343_5 gpc5196 (
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage3_7[0], stage3_7[1], stage3_7[2]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[2],stage4_5[4]}
   );
   gpc1343_5 gpc5197 (
      {stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_6[10], stage3_6[11], stage3_6[12], stage3_6[13]},
      {stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[1]},
      {stage4_9[1],stage4_8[2],stage4_7[2],stage4_6[3],stage4_5[5]}
   );
   gpc606_5 gpc5198 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[2],stage4_8[3],stage4_7[3],stage4_6[4],stage4_5[6]}
   );
   gpc606_5 gpc5199 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[3],stage4_8[4],stage4_7[4],stage4_6[5],stage4_5[7]}
   );
   gpc606_5 gpc5200 (
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23]},
      {stage4_9[4],stage4_8[5],stage4_7[5],stage4_6[6],stage4_5[8]}
   );
   gpc606_5 gpc5201 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[5]}
   );
   gpc615_5 gpc5202 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10]},
      {stage3_10[0]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[1],stage4_10[1],stage4_9[6]}
   );
   gpc615_5 gpc5203 (
      {stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15]},
      {stage3_10[1]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[2],stage4_11[2],stage4_10[2],stage4_9[7]}
   );
   gpc2135_5 gpc5204 (
      {stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage3_11[18], stage3_11[19], stage3_11[20]},
      {stage3_12[0]},
      {stage3_13[0], stage3_13[1]},
      {stage4_14[0],stage4_13[3],stage4_12[3],stage4_11[3],stage4_10[3]}
   );
   gpc2135_5 gpc5205 (
      {stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage3_12[1]},
      {stage3_13[2], stage3_13[3]},
      {stage4_14[1],stage4_13[4],stage4_12[4],stage4_11[4],stage4_10[4]}
   );
   gpc117_4 gpc5206 (
      {stage3_10[12], stage3_10[13], stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18]},
      {stage3_11[24]},
      {stage3_12[2]},
      {stage4_13[5],stage4_12[5],stage4_11[5],stage4_10[5]}
   );
   gpc117_4 gpc5207 (
      {stage3_10[19], stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24], stage3_10[25]},
      {stage3_11[25]},
      {stage3_12[3]},
      {stage4_13[6],stage4_12[6],stage4_11[6],stage4_10[6]}
   );
   gpc606_5 gpc5208 (
      {stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[2],stage4_13[7],stage4_12[7]}
   );
   gpc606_5 gpc5209 (
      {stage3_12[10], stage3_12[11], stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[1],stage4_14[3],stage4_13[8],stage4_12[8]}
   );
   gpc606_5 gpc5210 (
      {stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[2],stage4_15[2],stage4_14[4],stage4_13[9]}
   );
   gpc606_5 gpc5211 (
      {stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[3],stage4_15[3],stage4_14[5],stage4_13[10]}
   );
   gpc606_5 gpc5212 (
      {stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21]},
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17]},
      {stage4_17[2],stage4_16[4],stage4_15[4],stage4_14[6],stage4_13[11]}
   );
   gpc117_4 gpc5213 (
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17], stage3_14[18]},
      {stage3_15[18]},
      {stage3_16[0]},
      {stage4_17[3],stage4_16[5],stage4_15[5],stage4_14[7]}
   );
   gpc615_5 gpc5214 (
      {stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage3_15[19]},
      {stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5], stage3_16[6]},
      {stage4_18[0],stage4_17[4],stage4_16[6],stage4_15[6],stage4_14[8]}
   );
   gpc615_5 gpc5215 (
      {stage3_15[20], stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24]},
      {stage3_16[7]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[1],stage4_17[5],stage4_16[7],stage4_15[7]}
   );
   gpc615_5 gpc5216 (
      {stage3_15[25], stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29]},
      {stage3_16[8]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[2],stage4_17[6],stage4_16[8],stage4_15[8]}
   );
   gpc615_5 gpc5217 (
      {stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34]},
      {stage3_16[9]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[3],stage4_17[7],stage4_16[9],stage4_15[9]}
   );
   gpc615_5 gpc5218 (
      {stage3_15[35], stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39]},
      {stage3_16[10]},
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage4_19[3],stage4_18[4],stage4_17[8],stage4_16[10],stage4_15[10]}
   );
   gpc615_5 gpc5219 (
      {stage3_16[11], stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15]},
      {stage3_17[24]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[4],stage4_18[5],stage4_17[9],stage4_16[11]}
   );
   gpc615_5 gpc5220 (
      {stage3_16[16], stage3_16[17], stage3_16[18], stage3_16[19], 1'b0},
      {stage3_17[25]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[5],stage4_18[6],stage4_17[10],stage4_16[12]}
   );
   gpc615_5 gpc5221 (
      {stage3_18[12], stage3_18[13], stage3_18[14], stage3_18[15], stage3_18[16]},
      {stage3_19[0]},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage4_22[0],stage4_21[0],stage4_20[2],stage4_19[6],stage4_18[7]}
   );
   gpc615_5 gpc5222 (
      {stage3_18[17], stage3_18[18], stage3_18[19], stage3_18[20], stage3_18[21]},
      {stage3_19[1]},
      {stage3_20[6], stage3_20[7], stage3_20[8], stage3_20[9], stage3_20[10], stage3_20[11]},
      {stage4_22[1],stage4_21[1],stage4_20[3],stage4_19[7],stage4_18[8]}
   );
   gpc615_5 gpc5223 (
      {stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25], stage3_18[26]},
      {stage3_19[2]},
      {stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15], stage3_20[16], stage3_20[17]},
      {stage4_22[2],stage4_21[2],stage4_20[4],stage4_19[8],stage4_18[9]}
   );
   gpc215_4 gpc5224 (
      {stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6], stage3_19[7]},
      {stage3_20[18]},
      {stage3_21[0], stage3_21[1]},
      {stage4_22[3],stage4_21[3],stage4_20[5],stage4_19[9]}
   );
   gpc223_4 gpc5225 (
      {stage3_19[8], stage3_19[9], stage3_19[10]},
      {stage3_20[19], stage3_20[20]},
      {stage3_21[2], stage3_21[3]},
      {stage4_22[4],stage4_21[4],stage4_20[6],stage4_19[10]}
   );
   gpc207_4 gpc5226 (
      {stage3_19[11], stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17]},
      {stage3_21[4], stage3_21[5]},
      {stage4_22[5],stage4_21[5],stage4_20[7],stage4_19[11]}
   );
   gpc615_5 gpc5227 (
      {stage3_19[18], stage3_19[19], stage3_19[20], stage3_19[21], stage3_19[22]},
      {stage3_20[21]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[0],stage4_22[6],stage4_21[6],stage4_20[8],stage4_19[12]}
   );
   gpc615_5 gpc5228 (
      {stage3_19[23], stage3_19[24], stage3_19[25], stage3_19[26], stage3_19[27]},
      {stage3_20[22]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[1],stage4_22[7],stage4_21[7],stage4_20[9],stage4_19[13]}
   );
   gpc606_5 gpc5229 (
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[0],stage4_23[2],stage4_22[8],stage4_21[8]}
   );
   gpc2135_5 gpc5230 (
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4]},
      {stage3_23[6], stage3_23[7], stage3_23[8]},
      {stage3_24[0]},
      {stage3_25[0], stage3_25[1]},
      {stage4_26[0],stage4_25[1],stage4_24[1],stage4_23[3],stage4_22[9]}
   );
   gpc2135_5 gpc5231 (
      {stage3_22[5], stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9]},
      {stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage3_24[1]},
      {stage3_25[2], stage3_25[3]},
      {stage4_26[1],stage4_25[2],stage4_24[2],stage4_23[4],stage4_22[10]}
   );
   gpc615_5 gpc5232 (
      {stage3_22[10], stage3_22[11], stage3_22[12], stage3_22[13], stage3_22[14]},
      {stage3_23[12]},
      {stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6], stage3_24[7]},
      {stage4_26[2],stage4_25[3],stage4_24[3],stage4_23[5],stage4_22[11]}
   );
   gpc615_5 gpc5233 (
      {stage3_22[15], stage3_22[16], stage3_22[17], stage3_22[18], stage3_22[19]},
      {stage3_23[13]},
      {stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11], stage3_24[12], stage3_24[13]},
      {stage4_26[3],stage4_25[4],stage4_24[4],stage4_23[6],stage4_22[12]}
   );
   gpc615_5 gpc5234 (
      {stage3_22[20], stage3_22[21], stage3_22[22], stage3_22[23], stage3_22[24]},
      {stage3_23[14]},
      {stage3_24[14], stage3_24[15], stage3_24[16], stage3_24[17], stage3_24[18], stage3_24[19]},
      {stage4_26[4],stage4_25[5],stage4_24[5],stage4_23[7],stage4_22[13]}
   );
   gpc615_5 gpc5235 (
      {stage3_22[25], stage3_22[26], stage3_22[27], stage3_22[28], 1'b0},
      {stage3_23[15]},
      {stage3_24[20], stage3_24[21], stage3_24[22], stage3_24[23], stage3_24[24], stage3_24[25]},
      {stage4_26[5],stage4_25[6],stage4_24[6],stage4_23[8],stage4_22[14]}
   );
   gpc1163_5 gpc5236 (
      {stage3_25[4], stage3_25[5], stage3_25[6]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_27[0]},
      {stage3_28[0]},
      {stage4_29[0],stage4_28[0],stage4_27[0],stage4_26[6],stage4_25[7]}
   );
   gpc1163_5 gpc5237 (
      {stage3_25[7], stage3_25[8], stage3_25[9]},
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage3_27[1]},
      {stage3_28[1]},
      {stage4_29[1],stage4_28[1],stage4_27[1],stage4_26[7],stage4_25[8]}
   );
   gpc1163_5 gpc5238 (
      {stage3_25[10], stage3_25[11], stage3_25[12]},
      {stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15], stage3_26[16], stage3_26[17]},
      {stage3_27[2]},
      {stage3_28[2]},
      {stage4_29[2],stage4_28[2],stage4_27[2],stage4_26[8],stage4_25[9]}
   );
   gpc1163_5 gpc5239 (
      {stage3_25[13], stage3_25[14], stage3_25[15]},
      {stage3_26[18], stage3_26[19], stage3_26[20], stage3_26[21], stage3_26[22], stage3_26[23]},
      {stage3_27[3]},
      {stage3_28[3]},
      {stage4_29[3],stage4_28[3],stage4_27[3],stage4_26[9],stage4_25[10]}
   );
   gpc606_5 gpc5240 (
      {stage3_25[16], stage3_25[17], stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21]},
      {stage3_27[4], stage3_27[5], stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9]},
      {stage4_29[4],stage4_28[4],stage4_27[4],stage4_26[10],stage4_25[11]}
   );
   gpc606_5 gpc5241 (
      {stage3_25[22], stage3_25[23], stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27]},
      {stage3_27[10], stage3_27[11], stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15]},
      {stage4_29[5],stage4_28[5],stage4_27[5],stage4_26[11],stage4_25[12]}
   );
   gpc606_5 gpc5242 (
      {stage3_25[28], stage3_25[29], stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33]},
      {stage3_27[16], stage3_27[17], stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21]},
      {stage4_29[6],stage4_28[6],stage4_27[6],stage4_26[12],stage4_25[13]}
   );
   gpc606_5 gpc5243 (
      {stage3_28[4], stage3_28[5], stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[0],stage4_30[0],stage4_29[7],stage4_28[7]}
   );
   gpc606_5 gpc5244 (
      {stage3_28[10], stage3_28[11], stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[1],stage4_30[1],stage4_29[8],stage4_28[8]}
   );
   gpc606_5 gpc5245 (
      {stage3_28[16], stage3_28[17], stage3_28[18], stage3_28[19], stage3_28[20], stage3_28[21]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage4_32[2],stage4_31[2],stage4_30[2],stage4_29[9],stage4_28[9]}
   );
   gpc606_5 gpc5246 (
      {stage3_28[22], stage3_28[23], stage3_28[24], stage3_28[25], stage3_28[26], stage3_28[27]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage4_32[3],stage4_31[3],stage4_30[3],stage4_29[10],stage4_28[10]}
   );
   gpc606_5 gpc5247 (
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[4],stage4_31[4],stage4_30[4],stage4_29[11]}
   );
   gpc606_5 gpc5248 (
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11]},
      {stage4_33[1],stage4_32[5],stage4_31[5],stage4_30[5],stage4_29[12]}
   );
   gpc606_5 gpc5249 (
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17]},
      {stage4_33[2],stage4_32[6],stage4_31[6],stage4_30[6],stage4_29[13]}
   );
   gpc606_5 gpc5250 (
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21], stage3_31[22], stage3_31[23]},
      {stage4_33[3],stage4_32[7],stage4_31[7],stage4_30[7],stage4_29[14]}
   );
   gpc606_5 gpc5251 (
      {stage3_29[24], stage3_29[25], stage3_29[26], stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27], stage3_31[28], stage3_31[29]},
      {stage4_33[4],stage4_32[8],stage4_31[8],stage4_30[8],stage4_29[15]}
   );
   gpc606_5 gpc5252 (
      {stage3_29[30], stage3_29[31], stage3_29[32], stage3_29[33], stage3_29[34], 1'b0},
      {stage3_31[30], stage3_31[31], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage4_33[5],stage4_32[9],stage4_31[9],stage4_30[9],stage4_29[16]}
   );
   gpc606_5 gpc5253 (
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[0],stage4_34[0],stage4_33[6],stage4_32[10]}
   );
   gpc606_5 gpc5254 (
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage4_36[1],stage4_35[1],stage4_34[1],stage4_33[7],stage4_32[11]}
   );
   gpc606_5 gpc5255 (
      {stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15], stage3_32[16], stage3_32[17]},
      {stage3_34[12], stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage4_36[2],stage4_35[2],stage4_34[2],stage4_33[8],stage4_32[12]}
   );
   gpc606_5 gpc5256 (
      {stage3_32[18], stage3_32[19], stage3_32[20], stage3_32[21], stage3_32[22], stage3_32[23]},
      {stage3_34[18], stage3_34[19], stage3_34[20], stage3_34[21], stage3_34[22], stage3_34[23]},
      {stage4_36[3],stage4_35[3],stage4_34[3],stage4_33[9],stage4_32[13]}
   );
   gpc606_5 gpc5257 (
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[4],stage4_35[4],stage4_34[4],stage4_33[10]}
   );
   gpc606_5 gpc5258 (
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage3_35[6], stage3_35[7], stage3_35[8], stage3_35[9], stage3_35[10], stage3_35[11]},
      {stage4_37[1],stage4_36[5],stage4_35[5],stage4_34[5],stage4_33[11]}
   );
   gpc606_5 gpc5259 (
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage3_35[12], stage3_35[13], stage3_35[14], stage3_35[15], stage3_35[16], stage3_35[17]},
      {stage4_37[2],stage4_36[6],stage4_35[6],stage4_34[6],stage4_33[12]}
   );
   gpc606_5 gpc5260 (
      {stage3_33[18], stage3_33[19], stage3_33[20], stage3_33[21], stage3_33[22], stage3_33[23]},
      {stage3_35[18], stage3_35[19], stage3_35[20], stage3_35[21], stage3_35[22], stage3_35[23]},
      {stage4_37[3],stage4_36[7],stage4_35[7],stage4_34[7],stage4_33[13]}
   );
   gpc606_5 gpc5261 (
      {stage3_36[0], stage3_36[1], stage3_36[2], stage3_36[3], stage3_36[4], stage3_36[5]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5]},
      {stage4_40[0],stage4_39[0],stage4_38[0],stage4_37[4],stage4_36[8]}
   );
   gpc606_5 gpc5262 (
      {stage3_36[6], stage3_36[7], stage3_36[8], stage3_36[9], stage3_36[10], stage3_36[11]},
      {stage3_38[6], stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10], stage3_38[11]},
      {stage4_40[1],stage4_39[1],stage4_38[1],stage4_37[5],stage4_36[9]}
   );
   gpc606_5 gpc5263 (
      {stage3_36[12], stage3_36[13], stage3_36[14], stage3_36[15], stage3_36[16], stage3_36[17]},
      {stage3_38[12], stage3_38[13], stage3_38[14], stage3_38[15], stage3_38[16], stage3_38[17]},
      {stage4_40[2],stage4_39[2],stage4_38[2],stage4_37[6],stage4_36[10]}
   );
   gpc606_5 gpc5264 (
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[3],stage4_39[3],stage4_38[3],stage4_37[7]}
   );
   gpc606_5 gpc5265 (
      {stage3_37[6], stage3_37[7], stage3_37[8], stage3_37[9], stage3_37[10], stage3_37[11]},
      {stage3_39[6], stage3_39[7], stage3_39[8], stage3_39[9], stage3_39[10], stage3_39[11]},
      {stage4_41[1],stage4_40[4],stage4_39[4],stage4_38[4],stage4_37[8]}
   );
   gpc615_5 gpc5266 (
      {stage3_37[12], stage3_37[13], stage3_37[14], stage3_37[15], stage3_37[16]},
      {stage3_38[18]},
      {stage3_39[12], stage3_39[13], stage3_39[14], stage3_39[15], stage3_39[16], stage3_39[17]},
      {stage4_41[2],stage4_40[5],stage4_39[5],stage4_38[5],stage4_37[9]}
   );
   gpc615_5 gpc5267 (
      {stage3_38[19], stage3_38[20], stage3_38[21], stage3_38[22], 1'b0},
      {stage3_39[18]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[3],stage4_40[6],stage4_39[6],stage4_38[6]}
   );
   gpc606_5 gpc5268 (
      {stage3_39[19], stage3_39[20], stage3_39[21], stage3_39[22], stage3_39[23], stage3_39[24]},
      {stage3_41[0], stage3_41[1], stage3_41[2], stage3_41[3], stage3_41[4], stage3_41[5]},
      {stage4_43[0],stage4_42[1],stage4_41[4],stage4_40[7],stage4_39[7]}
   );
   gpc606_5 gpc5269 (
      {stage3_39[25], stage3_39[26], stage3_39[27], stage3_39[28], stage3_39[29], stage3_39[30]},
      {stage3_41[6], stage3_41[7], stage3_41[8], stage3_41[9], stage3_41[10], stage3_41[11]},
      {stage4_43[1],stage4_42[2],stage4_41[5],stage4_40[8],stage4_39[8]}
   );
   gpc606_5 gpc5270 (
      {stage3_40[6], stage3_40[7], stage3_40[8], stage3_40[9], stage3_40[10], stage3_40[11]},
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5]},
      {stage4_44[0],stage4_43[2],stage4_42[3],stage4_41[6],stage4_40[9]}
   );
   gpc606_5 gpc5271 (
      {stage3_40[12], stage3_40[13], stage3_40[14], stage3_40[15], stage3_40[16], stage3_40[17]},
      {stage3_42[6], stage3_42[7], stage3_42[8], stage3_42[9], stage3_42[10], stage3_42[11]},
      {stage4_44[1],stage4_43[3],stage4_42[4],stage4_41[7],stage4_40[10]}
   );
   gpc606_5 gpc5272 (
      {stage3_40[18], stage3_40[19], stage3_40[20], stage3_40[21], stage3_40[22], stage3_40[23]},
      {stage3_42[12], stage3_42[13], stage3_42[14], stage3_42[15], stage3_42[16], stage3_42[17]},
      {stage4_44[2],stage4_43[4],stage4_42[5],stage4_41[8],stage4_40[11]}
   );
   gpc606_5 gpc5273 (
      {stage3_40[24], stage3_40[25], stage3_40[26], stage3_40[27], stage3_40[28], stage3_40[29]},
      {stage3_42[18], stage3_42[19], stage3_42[20], stage3_42[21], stage3_42[22], stage3_42[23]},
      {stage4_44[3],stage4_43[5],stage4_42[6],stage4_41[9],stage4_40[12]}
   );
   gpc606_5 gpc5274 (
      {stage3_41[12], stage3_41[13], stage3_41[14], stage3_41[15], stage3_41[16], stage3_41[17]},
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4], stage3_43[5]},
      {stage4_45[0],stage4_44[4],stage4_43[6],stage4_42[7],stage4_41[10]}
   );
   gpc606_5 gpc5275 (
      {stage3_41[18], stage3_41[19], stage3_41[20], stage3_41[21], stage3_41[22], stage3_41[23]},
      {stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9], stage3_43[10], stage3_43[11]},
      {stage4_45[1],stage4_44[5],stage4_43[7],stage4_42[8],stage4_41[11]}
   );
   gpc606_5 gpc5276 (
      {stage3_43[12], stage3_43[13], stage3_43[14], stage3_43[15], stage3_43[16], stage3_43[17]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[0],stage4_45[2],stage4_44[6],stage4_43[8]}
   );
   gpc606_5 gpc5277 (
      {stage3_43[18], stage3_43[19], stage3_43[20], stage3_43[21], stage3_43[22], stage3_43[23]},
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9], stage3_45[10], stage3_45[11]},
      {stage4_47[1],stage4_46[1],stage4_45[3],stage4_44[7],stage4_43[9]}
   );
   gpc606_5 gpc5278 (
      {stage3_43[24], stage3_43[25], stage3_43[26], stage3_43[27], stage3_43[28], stage3_43[29]},
      {stage3_45[12], stage3_45[13], stage3_45[14], stage3_45[15], stage3_45[16], stage3_45[17]},
      {stage4_47[2],stage4_46[2],stage4_45[4],stage4_44[8],stage4_43[10]}
   );
   gpc606_5 gpc5279 (
      {stage3_44[0], stage3_44[1], stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5]},
      {stage3_46[0], stage3_46[1], stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage4_48[0],stage4_47[3],stage4_46[3],stage4_45[5],stage4_44[9]}
   );
   gpc615_5 gpc5280 (
      {stage3_44[6], stage3_44[7], stage3_44[8], stage3_44[9], stage3_44[10]},
      {stage3_45[18]},
      {stage3_46[6], stage3_46[7], stage3_46[8], stage3_46[9], stage3_46[10], stage3_46[11]},
      {stage4_48[1],stage4_47[4],stage4_46[4],stage4_45[6],stage4_44[10]}
   );
   gpc615_5 gpc5281 (
      {stage3_44[11], stage3_44[12], stage3_44[13], stage3_44[14], stage3_44[15]},
      {stage3_45[19]},
      {stage3_46[12], stage3_46[13], stage3_46[14], stage3_46[15], stage3_46[16], stage3_46[17]},
      {stage4_48[2],stage4_47[5],stage4_46[5],stage4_45[7],stage4_44[11]}
   );
   gpc615_5 gpc5282 (
      {stage3_44[16], stage3_44[17], stage3_44[18], stage3_44[19], stage3_44[20]},
      {stage3_45[20]},
      {stage3_46[18], stage3_46[19], stage3_46[20], stage3_46[21], stage3_46[22], stage3_46[23]},
      {stage4_48[3],stage4_47[6],stage4_46[6],stage4_45[8],stage4_44[12]}
   );
   gpc606_5 gpc5283 (
      {stage3_45[21], stage3_45[22], stage3_45[23], stage3_45[24], stage3_45[25], stage3_45[26]},
      {stage3_47[0], stage3_47[1], stage3_47[2], stage3_47[3], stage3_47[4], stage3_47[5]},
      {stage4_49[0],stage4_48[4],stage4_47[7],stage4_46[7],stage4_45[9]}
   );
   gpc606_5 gpc5284 (
      {stage3_45[27], stage3_45[28], stage3_45[29], stage3_45[30], stage3_45[31], stage3_45[32]},
      {stage3_47[6], stage3_47[7], stage3_47[8], stage3_47[9], stage3_47[10], stage3_47[11]},
      {stage4_49[1],stage4_48[5],stage4_47[8],stage4_46[8],stage4_45[10]}
   );
   gpc606_5 gpc5285 (
      {stage3_45[33], stage3_45[34], stage3_45[35], stage3_45[36], stage3_45[37], stage3_45[38]},
      {stage3_47[12], stage3_47[13], stage3_47[14], stage3_47[15], stage3_47[16], stage3_47[17]},
      {stage4_49[2],stage4_48[6],stage4_47[9],stage4_46[9],stage4_45[11]}
   );
   gpc1406_5 gpc5286 (
      {stage3_46[24], stage3_46[25], stage3_46[26], stage3_46[27], stage3_46[28], stage3_46[29]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3]},
      {stage3_49[0]},
      {stage4_50[0],stage4_49[3],stage4_48[7],stage4_47[10],stage4_46[10]}
   );
   gpc207_4 gpc5287 (
      {stage3_46[30], stage3_46[31], stage3_46[32], stage3_46[33], stage3_46[34], stage3_46[35], stage3_46[36]},
      {stage3_48[4], stage3_48[5]},
      {stage4_49[4],stage4_48[8],stage4_47[11],stage4_46[11]}
   );
   gpc615_5 gpc5288 (
      {stage3_47[18], stage3_47[19], stage3_47[20], stage3_47[21], stage3_47[22]},
      {stage3_48[6]},
      {stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5], stage3_49[6]},
      {stage4_51[0],stage4_50[1],stage4_49[5],stage4_48[9],stage4_47[12]}
   );
   gpc615_5 gpc5289 (
      {stage3_47[23], stage3_47[24], stage3_47[25], stage3_47[26], stage3_47[27]},
      {stage3_48[7]},
      {stage3_49[7], stage3_49[8], stage3_49[9], stage3_49[10], stage3_49[11], stage3_49[12]},
      {stage4_51[1],stage4_50[2],stage4_49[6],stage4_48[10],stage4_47[13]}
   );
   gpc615_5 gpc5290 (
      {stage3_47[28], stage3_47[29], stage3_47[30], stage3_47[31], stage3_47[32]},
      {stage3_48[8]},
      {stage3_49[13], stage3_49[14], stage3_49[15], stage3_49[16], stage3_49[17], stage3_49[18]},
      {stage4_51[2],stage4_50[3],stage4_49[7],stage4_48[11],stage4_47[14]}
   );
   gpc135_4 gpc5291 (
      {stage3_48[9], stage3_48[10], stage3_48[11], stage3_48[12], stage3_48[13]},
      {stage3_49[19], stage3_49[20], stage3_49[21]},
      {stage3_50[0]},
      {stage4_51[3],stage4_50[4],stage4_49[8],stage4_48[12]}
   );
   gpc135_4 gpc5292 (
      {stage3_48[14], stage3_48[15], stage3_48[16], stage3_48[17], stage3_48[18]},
      {stage3_49[22], stage3_49[23], stage3_49[24]},
      {stage3_50[1]},
      {stage4_51[4],stage4_50[5],stage4_49[9],stage4_48[13]}
   );
   gpc135_4 gpc5293 (
      {stage3_48[19], stage3_48[20], stage3_48[21], stage3_48[22], stage3_48[23]},
      {stage3_49[25], stage3_49[26], stage3_49[27]},
      {stage3_50[2]},
      {stage4_51[5],stage4_50[6],stage4_49[10],stage4_48[14]}
   );
   gpc606_5 gpc5294 (
      {stage3_49[28], stage3_49[29], stage3_49[30], stage3_49[31], stage3_49[32], stage3_49[33]},
      {stage3_51[0], stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage4_53[0],stage4_52[0],stage4_51[6],stage4_50[7],stage4_49[11]}
   );
   gpc606_5 gpc5295 (
      {stage3_49[34], stage3_49[35], stage3_49[36], stage3_49[37], stage3_49[38], stage3_49[39]},
      {stage3_51[6], stage3_51[7], stage3_51[8], stage3_51[9], stage3_51[10], stage3_51[11]},
      {stage4_53[1],stage4_52[1],stage4_51[7],stage4_50[8],stage4_49[12]}
   );
   gpc606_5 gpc5296 (
      {stage3_49[40], stage3_49[41], stage3_49[42], stage3_49[43], stage3_49[44], stage3_49[45]},
      {stage3_51[12], stage3_51[13], stage3_51[14], stage3_51[15], stage3_51[16], stage3_51[17]},
      {stage4_53[2],stage4_52[2],stage4_51[8],stage4_50[9],stage4_49[13]}
   );
   gpc615_5 gpc5297 (
      {stage3_50[3], stage3_50[4], stage3_50[5], stage3_50[6], stage3_50[7]},
      {stage3_51[18]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[3],stage4_52[3],stage4_51[9],stage4_50[10]}
   );
   gpc615_5 gpc5298 (
      {stage3_50[8], stage3_50[9], stage3_50[10], stage3_50[11], stage3_50[12]},
      {stage3_51[19]},
      {stage3_52[6], stage3_52[7], stage3_52[8], stage3_52[9], stage3_52[10], stage3_52[11]},
      {stage4_54[1],stage4_53[4],stage4_52[4],stage4_51[10],stage4_50[11]}
   );
   gpc615_5 gpc5299 (
      {stage3_50[13], stage3_50[14], stage3_50[15], stage3_50[16], stage3_50[17]},
      {stage3_51[20]},
      {stage3_52[12], stage3_52[13], stage3_52[14], stage3_52[15], stage3_52[16], stage3_52[17]},
      {stage4_54[2],stage4_53[5],stage4_52[5],stage4_51[11],stage4_50[12]}
   );
   gpc615_5 gpc5300 (
      {stage3_50[18], stage3_50[19], stage3_50[20], stage3_50[21], stage3_50[22]},
      {stage3_51[21]},
      {stage3_52[18], stage3_52[19], stage3_52[20], stage3_52[21], stage3_52[22], stage3_52[23]},
      {stage4_54[3],stage4_53[6],stage4_52[6],stage4_51[12],stage4_50[13]}
   );
   gpc615_5 gpc5301 (
      {stage3_50[23], stage3_50[24], stage3_50[25], stage3_50[26], stage3_50[27]},
      {stage3_51[22]},
      {stage3_52[24], stage3_52[25], stage3_52[26], stage3_52[27], stage3_52[28], stage3_52[29]},
      {stage4_54[4],stage4_53[7],stage4_52[7],stage4_51[13],stage4_50[14]}
   );
   gpc215_4 gpc5302 (
      {stage3_51[23], stage3_51[24], stage3_51[25], stage3_51[26], stage3_51[27]},
      {stage3_52[30]},
      {stage3_53[0], stage3_53[1]},
      {stage4_54[5],stage4_53[8],stage4_52[8],stage4_51[14]}
   );
   gpc215_4 gpc5303 (
      {stage3_51[28], stage3_51[29], stage3_51[30], stage3_51[31], stage3_51[32]},
      {stage3_52[31]},
      {stage3_53[2], stage3_53[3]},
      {stage4_54[6],stage4_53[9],stage4_52[9],stage4_51[15]}
   );
   gpc606_5 gpc5304 (
      {stage3_51[33], stage3_51[34], stage3_51[35], stage3_51[36], stage3_51[37], stage3_51[38]},
      {stage3_53[4], stage3_53[5], stage3_53[6], stage3_53[7], stage3_53[8], stage3_53[9]},
      {stage4_55[0],stage4_54[7],stage4_53[10],stage4_52[10],stage4_51[16]}
   );
   gpc615_5 gpc5305 (
      {stage3_51[39], stage3_51[40], stage3_51[41], stage3_51[42], stage3_51[43]},
      {stage3_52[32]},
      {stage3_53[10], stage3_53[11], stage3_53[12], stage3_53[13], stage3_53[14], stage3_53[15]},
      {stage4_55[1],stage4_54[8],stage4_53[11],stage4_52[11],stage4_51[17]}
   );
   gpc623_5 gpc5306 (
      {stage3_51[44], stage3_51[45], stage3_51[46]},
      {stage3_52[33], stage3_52[34]},
      {stage3_53[16], stage3_53[17], stage3_53[18], stage3_53[19], stage3_53[20], stage3_53[21]},
      {stage4_55[2],stage4_54[9],stage4_53[12],stage4_52[12],stage4_51[18]}
   );
   gpc606_5 gpc5307 (
      {stage3_52[35], stage3_52[36], stage3_52[37], stage3_52[38], stage3_52[39], 1'b0},
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage4_56[0],stage4_55[3],stage4_54[10],stage4_53[13],stage4_52[13]}
   );
   gpc606_5 gpc5308 (
      {stage3_53[22], stage3_53[23], stage3_53[24], stage3_53[25], stage3_53[26], stage3_53[27]},
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage4_57[0],stage4_56[1],stage4_55[4],stage4_54[11],stage4_53[14]}
   );
   gpc2135_5 gpc5309 (
      {stage3_54[6], stage3_54[7], stage3_54[8], stage3_54[9], stage3_54[10]},
      {stage3_55[6], stage3_55[7], stage3_55[8]},
      {stage3_56[0]},
      {stage3_57[0], stage3_57[1]},
      {stage4_58[0],stage4_57[1],stage4_56[2],stage4_55[5],stage4_54[12]}
   );
   gpc615_5 gpc5310 (
      {stage3_54[11], stage3_54[12], stage3_54[13], stage3_54[14], stage3_54[15]},
      {stage3_55[9]},
      {stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5], stage3_56[6]},
      {stage4_58[1],stage4_57[2],stage4_56[3],stage4_55[6],stage4_54[13]}
   );
   gpc615_5 gpc5311 (
      {stage3_54[16], stage3_54[17], stage3_54[18], stage3_54[19], stage3_54[20]},
      {stage3_55[10]},
      {stage3_56[7], stage3_56[8], stage3_56[9], stage3_56[10], stage3_56[11], stage3_56[12]},
      {stage4_58[2],stage4_57[3],stage4_56[4],stage4_55[7],stage4_54[14]}
   );
   gpc615_5 gpc5312 (
      {stage3_54[21], stage3_54[22], stage3_54[23], stage3_54[24], stage3_54[25]},
      {stage3_55[11]},
      {stage3_56[13], stage3_56[14], stage3_56[15], stage3_56[16], stage3_56[17], stage3_56[18]},
      {stage4_58[3],stage4_57[4],stage4_56[5],stage4_55[8],stage4_54[15]}
   );
   gpc615_5 gpc5313 (
      {stage3_55[12], stage3_55[13], stage3_55[14], stage3_55[15], stage3_55[16]},
      {stage3_56[19]},
      {stage3_57[2], stage3_57[3], stage3_57[4], stage3_57[5], stage3_57[6], stage3_57[7]},
      {stage4_59[0],stage4_58[4],stage4_57[5],stage4_56[6],stage4_55[9]}
   );
   gpc615_5 gpc5314 (
      {stage3_55[17], stage3_55[18], stage3_55[19], stage3_55[20], stage3_55[21]},
      {stage3_56[20]},
      {stage3_57[8], stage3_57[9], stage3_57[10], stage3_57[11], stage3_57[12], stage3_57[13]},
      {stage4_59[1],stage4_58[5],stage4_57[6],stage4_56[7],stage4_55[10]}
   );
   gpc615_5 gpc5315 (
      {stage3_55[22], stage3_55[23], stage3_55[24], stage3_55[25], stage3_55[26]},
      {stage3_56[21]},
      {stage3_57[14], stage3_57[15], stage3_57[16], stage3_57[17], stage3_57[18], stage3_57[19]},
      {stage4_59[2],stage4_58[6],stage4_57[7],stage4_56[8],stage4_55[11]}
   );
   gpc623_5 gpc5316 (
      {stage3_55[27], stage3_55[28], stage3_55[29]},
      {stage3_56[22], stage3_56[23]},
      {stage3_57[20], stage3_57[21], stage3_57[22], stage3_57[23], stage3_57[24], stage3_57[25]},
      {stage4_59[3],stage4_58[7],stage4_57[8],stage4_56[9],stage4_55[12]}
   );
   gpc615_5 gpc5317 (
      {stage3_57[26], stage3_57[27], stage3_57[28], stage3_57[29], stage3_57[30]},
      {stage3_58[0]},
      {stage3_59[0], stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5]},
      {stage4_61[0],stage4_60[0],stage4_59[4],stage4_58[8],stage4_57[9]}
   );
   gpc2135_5 gpc5318 (
      {stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5]},
      {stage3_59[6], stage3_59[7], stage3_59[8]},
      {stage3_60[0]},
      {stage3_61[0], stage3_61[1]},
      {stage4_62[0],stage4_61[1],stage4_60[1],stage4_59[5],stage4_58[9]}
   );
   gpc2135_5 gpc5319 (
      {stage3_58[6], stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10]},
      {stage3_59[9], stage3_59[10], stage3_59[11]},
      {stage3_60[1]},
      {stage3_61[2], stage3_61[3]},
      {stage4_62[1],stage4_61[2],stage4_60[2],stage4_59[6],stage4_58[10]}
   );
   gpc2135_5 gpc5320 (
      {stage3_58[11], stage3_58[12], stage3_58[13], stage3_58[14], stage3_58[15]},
      {stage3_59[12], stage3_59[13], stage3_59[14]},
      {stage3_60[2]},
      {stage3_61[4], stage3_61[5]},
      {stage4_62[2],stage4_61[3],stage4_60[3],stage4_59[7],stage4_58[11]}
   );
   gpc606_5 gpc5321 (
      {stage3_58[16], stage3_58[17], stage3_58[18], stage3_58[19], stage3_58[20], stage3_58[21]},
      {stage3_60[3], stage3_60[4], stage3_60[5], stage3_60[6], stage3_60[7], stage3_60[8]},
      {stage4_62[3],stage4_61[4],stage4_60[4],stage4_59[8],stage4_58[12]}
   );
   gpc606_5 gpc5322 (
      {stage3_59[15], stage3_59[16], stage3_59[17], stage3_59[18], stage3_59[19], stage3_59[20]},
      {stage3_61[6], stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11]},
      {stage4_63[0],stage4_62[4],stage4_61[5],stage4_60[5],stage4_59[9]}
   );
   gpc606_5 gpc5323 (
      {stage3_59[21], stage3_59[22], stage3_59[23], stage3_59[24], stage3_59[25], stage3_59[26]},
      {stage3_61[12], stage3_61[13], stage3_61[14], stage3_61[15], stage3_61[16], stage3_61[17]},
      {stage4_63[1],stage4_62[5],stage4_61[6],stage4_60[6],stage4_59[10]}
   );
   gpc606_5 gpc5324 (
      {stage3_59[27], stage3_59[28], stage3_59[29], stage3_59[30], stage3_59[31], stage3_59[32]},
      {stage3_61[18], stage3_61[19], stage3_61[20], stage3_61[21], stage3_61[22], stage3_61[23]},
      {stage4_63[2],stage4_62[6],stage4_61[7],stage4_60[7],stage4_59[11]}
   );
   gpc606_5 gpc5325 (
      {stage3_60[9], stage3_60[10], stage3_60[11], stage3_60[12], stage3_60[13], stage3_60[14]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], stage3_62[5]},
      {stage4_64[0],stage4_63[3],stage4_62[7],stage4_61[8],stage4_60[8]}
   );
   gpc606_5 gpc5326 (
      {stage3_60[15], stage3_60[16], stage3_60[17], stage3_60[18], stage3_60[19], stage3_60[20]},
      {stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9], stage3_62[10], stage3_62[11]},
      {stage4_64[1],stage4_63[4],stage4_62[8],stage4_61[9],stage4_60[9]}
   );
   gpc606_5 gpc5327 (
      {stage3_60[21], stage3_60[22], stage3_60[23], stage3_60[24], stage3_60[25], stage3_60[26]},
      {stage3_62[12], stage3_62[13], stage3_62[14], stage3_62[15], stage3_62[16], stage3_62[17]},
      {stage4_64[2],stage4_63[5],stage4_62[9],stage4_61[10],stage4_60[10]}
   );
   gpc606_5 gpc5328 (
      {stage3_60[27], stage3_60[28], stage3_60[29], stage3_60[30], stage3_60[31], stage3_60[32]},
      {stage3_62[18], stage3_62[19], stage3_62[20], stage3_62[21], stage3_62[22], stage3_62[23]},
      {stage4_64[3],stage4_63[6],stage4_62[10],stage4_61[11],stage4_60[11]}
   );
   gpc606_5 gpc5329 (
      {stage3_62[24], stage3_62[25], stage3_62[26], stage3_62[27], 1'b0, 1'b0},
      {stage3_64[0], stage3_64[1], stage3_64[2], stage3_64[3], stage3_64[4], stage3_64[5]},
      {stage4_66[0],stage4_65[0],stage4_64[4],stage4_63[7],stage4_62[11]}
   );
   gpc606_5 gpc5330 (
      {stage3_63[0], stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[1],stage4_65[1],stage4_64[5],stage4_63[8]}
   );
   gpc606_5 gpc5331 (
      {stage3_63[6], stage3_63[7], stage3_63[8], stage3_63[9], stage3_63[10], stage3_63[11]},
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage4_67[1],stage4_66[2],stage4_65[2],stage4_64[6],stage4_63[9]}
   );
   gpc606_5 gpc5332 (
      {stage3_63[12], stage3_63[13], stage3_63[14], stage3_63[15], stage3_63[16], stage3_63[17]},
      {stage3_65[12], stage3_65[13], stage3_65[14], stage3_65[15], stage3_65[16], stage3_65[17]},
      {stage4_67[2],stage4_66[3],stage4_65[3],stage4_64[7],stage4_63[10]}
   );
   gpc606_5 gpc5333 (
      {stage3_63[18], stage3_63[19], stage3_63[20], stage3_63[21], stage3_63[22], stage3_63[23]},
      {stage3_65[18], stage3_65[19], stage3_65[20], stage3_65[21], stage3_65[22], stage3_65[23]},
      {stage4_67[3],stage4_66[4],stage4_65[4],stage4_64[8],stage4_63[11]}
   );
   gpc606_5 gpc5334 (
      {stage3_63[24], stage3_63[25], stage3_63[26], stage3_63[27], 1'b0, 1'b0},
      {stage3_65[24], stage3_65[25], stage3_65[26], stage3_65[27], 1'b0, 1'b0},
      {stage4_67[4],stage4_66[5],stage4_65[5],stage4_64[9],stage4_63[12]}
   );
   gpc606_5 gpc5335 (
      {stage3_64[6], stage3_64[7], stage3_64[8], stage3_64[9], stage3_64[10], stage3_64[11]},
      {stage3_66[0], stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5]},
      {stage4_68[0],stage4_67[5],stage4_66[6],stage4_65[6],stage4_64[10]}
   );
   gpc606_5 gpc5336 (
      {stage3_64[12], stage3_64[13], stage3_64[14], stage3_64[15], stage3_64[16], stage3_64[17]},
      {stage3_66[6], stage3_66[7], stage3_66[8], stage3_66[9], stage3_66[10], stage3_66[11]},
      {stage4_68[1],stage4_67[6],stage4_66[7],stage4_65[7],stage4_64[11]}
   );
   gpc1_1 gpc5337 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc5338 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc5339 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc5340 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc5341 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc5342 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc5343 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc5344 (
      {stage3_0[7]},
      {stage4_0[7]}
   );
   gpc1_1 gpc5345 (
      {stage3_0[8]},
      {stage4_0[8]}
   );
   gpc1_1 gpc5346 (
      {stage3_0[9]},
      {stage4_0[9]}
   );
   gpc1_1 gpc5347 (
      {stage3_0[10]},
      {stage4_0[10]}
   );
   gpc1_1 gpc5348 (
      {stage3_0[11]},
      {stage4_0[11]}
   );
   gpc1_1 gpc5349 (
      {stage3_0[12]},
      {stage4_0[12]}
   );
   gpc1_1 gpc5350 (
      {stage3_0[13]},
      {stage4_0[13]}
   );
   gpc1_1 gpc5351 (
      {stage3_1[8]},
      {stage4_1[2]}
   );
   gpc1_1 gpc5352 (
      {stage3_1[9]},
      {stage4_1[3]}
   );
   gpc1_1 gpc5353 (
      {stage3_1[10]},
      {stage4_1[4]}
   );
   gpc1_1 gpc5354 (
      {stage3_2[14]},
      {stage4_2[3]}
   );
   gpc1_1 gpc5355 (
      {stage3_2[15]},
      {stage4_2[4]}
   );
   gpc1_1 gpc5356 (
      {stage3_2[16]},
      {stage4_2[5]}
   );
   gpc1_1 gpc5357 (
      {stage3_2[17]},
      {stage4_2[6]}
   );
   gpc1_1 gpc5358 (
      {stage3_3[3]},
      {stage4_3[3]}
   );
   gpc1_1 gpc5359 (
      {stage3_3[4]},
      {stage4_3[4]}
   );
   gpc1_1 gpc5360 (
      {stage3_3[5]},
      {stage4_3[5]}
   );
   gpc1_1 gpc5361 (
      {stage3_3[6]},
      {stage4_3[6]}
   );
   gpc1_1 gpc5362 (
      {stage3_3[7]},
      {stage4_3[7]}
   );
   gpc1_1 gpc5363 (
      {stage3_3[8]},
      {stage4_3[8]}
   );
   gpc1_1 gpc5364 (
      {stage3_3[9]},
      {stage4_3[9]}
   );
   gpc1_1 gpc5365 (
      {stage3_3[10]},
      {stage4_3[10]}
   );
   gpc1_1 gpc5366 (
      {stage3_3[11]},
      {stage4_3[11]}
   );
   gpc1_1 gpc5367 (
      {stage3_3[12]},
      {stage4_3[12]}
   );
   gpc1_1 gpc5368 (
      {stage3_3[13]},
      {stage4_3[13]}
   );
   gpc1_1 gpc5369 (
      {stage3_3[14]},
      {stage4_3[14]}
   );
   gpc1_1 gpc5370 (
      {stage3_3[15]},
      {stage4_3[15]}
   );
   gpc1_1 gpc5371 (
      {stage3_3[16]},
      {stage4_3[16]}
   );
   gpc1_1 gpc5372 (
      {stage3_3[17]},
      {stage4_3[17]}
   );
   gpc1_1 gpc5373 (
      {stage3_3[18]},
      {stage4_3[18]}
   );
   gpc1_1 gpc5374 (
      {stage3_4[15]},
      {stage4_4[4]}
   );
   gpc1_1 gpc5375 (
      {stage3_4[16]},
      {stage4_4[5]}
   );
   gpc1_1 gpc5376 (
      {stage3_4[17]},
      {stage4_4[6]}
   );
   gpc1_1 gpc5377 (
      {stage3_4[18]},
      {stage4_4[7]}
   );
   gpc1_1 gpc5378 (
      {stage3_4[19]},
      {stage4_4[8]}
   );
   gpc1_1 gpc5379 (
      {stage3_4[20]},
      {stage4_4[9]}
   );
   gpc1_1 gpc5380 (
      {stage3_5[24]},
      {stage4_5[9]}
   );
   gpc1_1 gpc5381 (
      {stage3_5[25]},
      {stage4_5[10]}
   );
   gpc1_1 gpc5382 (
      {stage3_5[26]},
      {stage4_5[11]}
   );
   gpc1_1 gpc5383 (
      {stage3_5[27]},
      {stage4_5[12]}
   );
   gpc1_1 gpc5384 (
      {stage3_5[28]},
      {stage4_5[13]}
   );
   gpc1_1 gpc5385 (
      {stage3_5[29]},
      {stage4_5[14]}
   );
   gpc1_1 gpc5386 (
      {stage3_5[30]},
      {stage4_5[15]}
   );
   gpc1_1 gpc5387 (
      {stage3_5[31]},
      {stage4_5[16]}
   );
   gpc1_1 gpc5388 (
      {stage3_5[32]},
      {stage4_5[17]}
   );
   gpc1_1 gpc5389 (
      {stage3_5[33]},
      {stage4_5[18]}
   );
   gpc1_1 gpc5390 (
      {stage3_5[34]},
      {stage4_5[19]}
   );
   gpc1_1 gpc5391 (
      {stage3_6[14]},
      {stage4_6[7]}
   );
   gpc1_1 gpc5392 (
      {stage3_6[15]},
      {stage4_6[8]}
   );
   gpc1_1 gpc5393 (
      {stage3_6[16]},
      {stage4_6[9]}
   );
   gpc1_1 gpc5394 (
      {stage3_7[24]},
      {stage4_7[6]}
   );
   gpc1_1 gpc5395 (
      {stage3_7[25]},
      {stage4_7[7]}
   );
   gpc1_1 gpc5396 (
      {stage3_7[26]},
      {stage4_7[8]}
   );
   gpc1_1 gpc5397 (
      {stage3_7[27]},
      {stage4_7[9]}
   );
   gpc1_1 gpc5398 (
      {stage3_8[2]},
      {stage4_8[6]}
   );
   gpc1_1 gpc5399 (
      {stage3_8[3]},
      {stage4_8[7]}
   );
   gpc1_1 gpc5400 (
      {stage3_8[4]},
      {stage4_8[8]}
   );
   gpc1_1 gpc5401 (
      {stage3_8[5]},
      {stage4_8[9]}
   );
   gpc1_1 gpc5402 (
      {stage3_8[6]},
      {stage4_8[10]}
   );
   gpc1_1 gpc5403 (
      {stage3_8[7]},
      {stage4_8[11]}
   );
   gpc1_1 gpc5404 (
      {stage3_8[8]},
      {stage4_8[12]}
   );
   gpc1_1 gpc5405 (
      {stage3_8[9]},
      {stage4_8[13]}
   );
   gpc1_1 gpc5406 (
      {stage3_8[10]},
      {stage4_8[14]}
   );
   gpc1_1 gpc5407 (
      {stage3_8[11]},
      {stage4_8[15]}
   );
   gpc1_1 gpc5408 (
      {stage3_8[12]},
      {stage4_8[16]}
   );
   gpc1_1 gpc5409 (
      {stage3_8[13]},
      {stage4_8[17]}
   );
   gpc1_1 gpc5410 (
      {stage3_8[14]},
      {stage4_8[18]}
   );
   gpc1_1 gpc5411 (
      {stage3_8[15]},
      {stage4_8[19]}
   );
   gpc1_1 gpc5412 (
      {stage3_8[16]},
      {stage4_8[20]}
   );
   gpc1_1 gpc5413 (
      {stage3_8[17]},
      {stage4_8[21]}
   );
   gpc1_1 gpc5414 (
      {stage3_10[26]},
      {stage4_10[7]}
   );
   gpc1_1 gpc5415 (
      {stage3_10[27]},
      {stage4_10[8]}
   );
   gpc1_1 gpc5416 (
      {stage3_10[28]},
      {stage4_10[9]}
   );
   gpc1_1 gpc5417 (
      {stage3_10[29]},
      {stage4_10[10]}
   );
   gpc1_1 gpc5418 (
      {stage3_10[30]},
      {stage4_10[11]}
   );
   gpc1_1 gpc5419 (
      {stage3_10[31]},
      {stage4_10[12]}
   );
   gpc1_1 gpc5420 (
      {stage3_10[32]},
      {stage4_10[13]}
   );
   gpc1_1 gpc5421 (
      {stage3_11[26]},
      {stage4_11[7]}
   );
   gpc1_1 gpc5422 (
      {stage3_11[27]},
      {stage4_11[8]}
   );
   gpc1_1 gpc5423 (
      {stage3_11[28]},
      {stage4_11[9]}
   );
   gpc1_1 gpc5424 (
      {stage3_11[29]},
      {stage4_11[10]}
   );
   gpc1_1 gpc5425 (
      {stage3_11[30]},
      {stage4_11[11]}
   );
   gpc1_1 gpc5426 (
      {stage3_12[16]},
      {stage4_12[9]}
   );
   gpc1_1 gpc5427 (
      {stage3_12[17]},
      {stage4_12[10]}
   );
   gpc1_1 gpc5428 (
      {stage3_12[18]},
      {stage4_12[11]}
   );
   gpc1_1 gpc5429 (
      {stage3_12[19]},
      {stage4_12[12]}
   );
   gpc1_1 gpc5430 (
      {stage3_12[20]},
      {stage4_12[13]}
   );
   gpc1_1 gpc5431 (
      {stage3_12[21]},
      {stage4_12[14]}
   );
   gpc1_1 gpc5432 (
      {stage3_12[22]},
      {stage4_12[15]}
   );
   gpc1_1 gpc5433 (
      {stage3_12[23]},
      {stage4_12[16]}
   );
   gpc1_1 gpc5434 (
      {stage3_12[24]},
      {stage4_12[17]}
   );
   gpc1_1 gpc5435 (
      {stage3_13[22]},
      {stage4_13[12]}
   );
   gpc1_1 gpc5436 (
      {stage3_13[23]},
      {stage4_13[13]}
   );
   gpc1_1 gpc5437 (
      {stage3_14[24]},
      {stage4_14[9]}
   );
   gpc1_1 gpc5438 (
      {stage3_14[25]},
      {stage4_14[10]}
   );
   gpc1_1 gpc5439 (
      {stage3_14[26]},
      {stage4_14[11]}
   );
   gpc1_1 gpc5440 (
      {stage3_15[40]},
      {stage4_15[11]}
   );
   gpc1_1 gpc5441 (
      {stage3_17[26]},
      {stage4_17[11]}
   );
   gpc1_1 gpc5442 (
      {stage3_17[27]},
      {stage4_17[12]}
   );
   gpc1_1 gpc5443 (
      {stage3_17[28]},
      {stage4_17[13]}
   );
   gpc1_1 gpc5444 (
      {stage3_17[29]},
      {stage4_17[14]}
   );
   gpc1_1 gpc5445 (
      {stage3_18[27]},
      {stage4_18[10]}
   );
   gpc1_1 gpc5446 (
      {stage3_20[23]},
      {stage4_20[10]}
   );
   gpc1_1 gpc5447 (
      {stage3_24[26]},
      {stage4_24[7]}
   );
   gpc1_1 gpc5448 (
      {stage3_24[27]},
      {stage4_24[8]}
   );
   gpc1_1 gpc5449 (
      {stage3_24[28]},
      {stage4_24[9]}
   );
   gpc1_1 gpc5450 (
      {stage3_24[29]},
      {stage4_24[10]}
   );
   gpc1_1 gpc5451 (
      {stage3_24[30]},
      {stage4_24[11]}
   );
   gpc1_1 gpc5452 (
      {stage3_28[28]},
      {stage4_28[11]}
   );
   gpc1_1 gpc5453 (
      {stage3_30[24]},
      {stage4_30[10]}
   );
   gpc1_1 gpc5454 (
      {stage3_30[25]},
      {stage4_30[11]}
   );
   gpc1_1 gpc5455 (
      {stage3_32[24]},
      {stage4_32[14]}
   );
   gpc1_1 gpc5456 (
      {stage3_32[25]},
      {stage4_32[15]}
   );
   gpc1_1 gpc5457 (
      {stage3_32[26]},
      {stage4_32[16]}
   );
   gpc1_1 gpc5458 (
      {stage3_32[27]},
      {stage4_32[17]}
   );
   gpc1_1 gpc5459 (
      {stage3_33[24]},
      {stage4_33[14]}
   );
   gpc1_1 gpc5460 (
      {stage3_33[25]},
      {stage4_33[15]}
   );
   gpc1_1 gpc5461 (
      {stage3_33[26]},
      {stage4_33[16]}
   );
   gpc1_1 gpc5462 (
      {stage3_34[24]},
      {stage4_34[8]}
   );
   gpc1_1 gpc5463 (
      {stage3_34[25]},
      {stage4_34[9]}
   );
   gpc1_1 gpc5464 (
      {stage3_34[26]},
      {stage4_34[10]}
   );
   gpc1_1 gpc5465 (
      {stage3_35[24]},
      {stage4_35[8]}
   );
   gpc1_1 gpc5466 (
      {stage3_35[25]},
      {stage4_35[9]}
   );
   gpc1_1 gpc5467 (
      {stage3_35[26]},
      {stage4_35[10]}
   );
   gpc1_1 gpc5468 (
      {stage3_35[27]},
      {stage4_35[11]}
   );
   gpc1_1 gpc5469 (
      {stage3_35[28]},
      {stage4_35[12]}
   );
   gpc1_1 gpc5470 (
      {stage3_35[29]},
      {stage4_35[13]}
   );
   gpc1_1 gpc5471 (
      {stage3_35[30]},
      {stage4_35[14]}
   );
   gpc1_1 gpc5472 (
      {stage3_35[31]},
      {stage4_35[15]}
   );
   gpc1_1 gpc5473 (
      {stage3_35[32]},
      {stage4_35[16]}
   );
   gpc1_1 gpc5474 (
      {stage3_36[18]},
      {stage4_36[11]}
   );
   gpc1_1 gpc5475 (
      {stage3_36[19]},
      {stage4_36[12]}
   );
   gpc1_1 gpc5476 (
      {stage3_37[17]},
      {stage4_37[10]}
   );
   gpc1_1 gpc5477 (
      {stage3_37[18]},
      {stage4_37[11]}
   );
   gpc1_1 gpc5478 (
      {stage3_42[24]},
      {stage4_42[9]}
   );
   gpc1_1 gpc5479 (
      {stage3_42[25]},
      {stage4_42[10]}
   );
   gpc1_1 gpc5480 (
      {stage3_42[26]},
      {stage4_42[11]}
   );
   gpc1_1 gpc5481 (
      {stage3_42[27]},
      {stage4_42[12]}
   );
   gpc1_1 gpc5482 (
      {stage3_42[28]},
      {stage4_42[13]}
   );
   gpc1_1 gpc5483 (
      {stage3_42[29]},
      {stage4_42[14]}
   );
   gpc1_1 gpc5484 (
      {stage3_43[30]},
      {stage4_43[11]}
   );
   gpc1_1 gpc5485 (
      {stage3_43[31]},
      {stage4_43[12]}
   );
   gpc1_1 gpc5486 (
      {stage3_43[32]},
      {stage4_43[13]}
   );
   gpc1_1 gpc5487 (
      {stage3_43[33]},
      {stage4_43[14]}
   );
   gpc1_1 gpc5488 (
      {stage3_43[34]},
      {stage4_43[15]}
   );
   gpc1_1 gpc5489 (
      {stage3_43[35]},
      {stage4_43[16]}
   );
   gpc1_1 gpc5490 (
      {stage3_43[36]},
      {stage4_43[17]}
   );
   gpc1_1 gpc5491 (
      {stage3_43[37]},
      {stage4_43[18]}
   );
   gpc1_1 gpc5492 (
      {stage3_43[38]},
      {stage4_43[19]}
   );
   gpc1_1 gpc5493 (
      {stage3_44[21]},
      {stage4_44[13]}
   );
   gpc1_1 gpc5494 (
      {stage3_46[37]},
      {stage4_46[12]}
   );
   gpc1_1 gpc5495 (
      {stage3_46[38]},
      {stage4_46[13]}
   );
   gpc1_1 gpc5496 (
      {stage3_46[39]},
      {stage4_46[14]}
   );
   gpc1_1 gpc5497 (
      {stage3_49[46]},
      {stage4_49[14]}
   );
   gpc1_1 gpc5498 (
      {stage3_49[47]},
      {stage4_49[15]}
   );
   gpc1_1 gpc5499 (
      {stage3_49[48]},
      {stage4_49[16]}
   );
   gpc1_1 gpc5500 (
      {stage3_49[49]},
      {stage4_49[17]}
   );
   gpc1_1 gpc5501 (
      {stage3_49[50]},
      {stage4_49[18]}
   );
   gpc1_1 gpc5502 (
      {stage3_49[51]},
      {stage4_49[19]}
   );
   gpc1_1 gpc5503 (
      {stage3_49[52]},
      {stage4_49[20]}
   );
   gpc1_1 gpc5504 (
      {stage3_49[53]},
      {stage4_49[21]}
   );
   gpc1_1 gpc5505 (
      {stage3_49[54]},
      {stage4_49[22]}
   );
   gpc1_1 gpc5506 (
      {stage3_49[55]},
      {stage4_49[23]}
   );
   gpc1_1 gpc5507 (
      {stage3_49[56]},
      {stage4_49[24]}
   );
   gpc1_1 gpc5508 (
      {stage3_49[57]},
      {stage4_49[25]}
   );
   gpc1_1 gpc5509 (
      {stage3_49[58]},
      {stage4_49[26]}
   );
   gpc1_1 gpc5510 (
      {stage3_49[59]},
      {stage4_49[27]}
   );
   gpc1_1 gpc5511 (
      {stage3_49[60]},
      {stage4_49[28]}
   );
   gpc1_1 gpc5512 (
      {stage3_49[61]},
      {stage4_49[29]}
   );
   gpc1_1 gpc5513 (
      {stage3_49[62]},
      {stage4_49[30]}
   );
   gpc1_1 gpc5514 (
      {stage3_49[63]},
      {stage4_49[31]}
   );
   gpc1_1 gpc5515 (
      {stage3_49[64]},
      {stage4_49[32]}
   );
   gpc1_1 gpc5516 (
      {stage3_49[65]},
      {stage4_49[33]}
   );
   gpc1_1 gpc5517 (
      {stage3_49[66]},
      {stage4_49[34]}
   );
   gpc1_1 gpc5518 (
      {stage3_49[67]},
      {stage4_49[35]}
   );
   gpc1_1 gpc5519 (
      {stage3_50[28]},
      {stage4_50[15]}
   );
   gpc1_1 gpc5520 (
      {stage3_50[29]},
      {stage4_50[16]}
   );
   gpc1_1 gpc5521 (
      {stage3_51[47]},
      {stage4_51[19]}
   );
   gpc1_1 gpc5522 (
      {stage3_54[26]},
      {stage4_54[16]}
   );
   gpc1_1 gpc5523 (
      {stage3_54[27]},
      {stage4_54[17]}
   );
   gpc1_1 gpc5524 (
      {stage3_56[24]},
      {stage4_56[10]}
   );
   gpc1_1 gpc5525 (
      {stage3_56[25]},
      {stage4_56[11]}
   );
   gpc1_1 gpc5526 (
      {stage3_57[31]},
      {stage4_57[10]}
   );
   gpc1_1 gpc5527 (
      {stage3_57[32]},
      {stage4_57[11]}
   );
   gpc1_1 gpc5528 (
      {stage3_58[22]},
      {stage4_58[13]}
   );
   gpc1_1 gpc5529 (
      {stage3_58[23]},
      {stage4_58[14]}
   );
   gpc1_1 gpc5530 (
      {stage3_58[24]},
      {stage4_58[15]}
   );
   gpc1_1 gpc5531 (
      {stage3_58[25]},
      {stage4_58[16]}
   );
   gpc1_1 gpc5532 (
      {stage3_58[26]},
      {stage4_58[17]}
   );
   gpc1_1 gpc5533 (
      {stage3_58[27]},
      {stage4_58[18]}
   );
   gpc1_1 gpc5534 (
      {stage3_58[28]},
      {stage4_58[19]}
   );
   gpc1_1 gpc5535 (
      {stage3_60[33]},
      {stage4_60[12]}
   );
   gpc1_1 gpc5536 (
      {stage3_60[34]},
      {stage4_60[13]}
   );
   gpc1_1 gpc5537 (
      {stage3_66[12]},
      {stage4_66[8]}
   );
   gpc1_1 gpc5538 (
      {stage3_66[13]},
      {stage4_66[9]}
   );
   gpc1_1 gpc5539 (
      {stage3_66[14]},
      {stage4_66[10]}
   );
   gpc1_1 gpc5540 (
      {stage3_66[15]},
      {stage4_66[11]}
   );
   gpc1_1 gpc5541 (
      {stage3_66[16]},
      {stage4_66[12]}
   );
   gpc1_1 gpc5542 (
      {stage3_66[17]},
      {stage4_66[13]}
   );
   gpc1_1 gpc5543 (
      {stage3_66[18]},
      {stage4_66[14]}
   );
   gpc1_1 gpc5544 (
      {stage3_66[19]},
      {stage4_66[15]}
   );
   gpc1_1 gpc5545 (
      {stage3_66[20]},
      {stage4_66[16]}
   );
   gpc1_1 gpc5546 (
      {stage3_66[21]},
      {stage4_66[17]}
   );
   gpc1_1 gpc5547 (
      {stage3_66[22]},
      {stage4_66[18]}
   );
   gpc1_1 gpc5548 (
      {stage3_66[23]},
      {stage4_66[19]}
   );
   gpc1_1 gpc5549 (
      {stage3_66[24]},
      {stage4_66[20]}
   );
   gpc1_1 gpc5550 (
      {stage3_66[25]},
      {stage4_66[21]}
   );
   gpc1_1 gpc5551 (
      {stage3_66[26]},
      {stage4_66[22]}
   );
   gpc1_1 gpc5552 (
      {stage3_66[27]},
      {stage4_66[23]}
   );
   gpc1_1 gpc5553 (
      {stage3_67[0]},
      {stage4_67[7]}
   );
   gpc1_1 gpc5554 (
      {stage3_67[1]},
      {stage4_67[8]}
   );
   gpc1_1 gpc5555 (
      {stage3_68[0]},
      {stage4_68[2]}
   );
   gpc1_1 gpc5556 (
      {stage3_69[0]},
      {stage4_69[0]}
   );
   gpc2135_5 gpc5557 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0]},
      {stage4_3[0], stage4_3[1]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc606_5 gpc5558 (
      {stage4_0[5], stage4_0[6], stage4_0[7], stage4_0[8], stage4_0[9], stage4_0[10]},
      {stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5], stage4_2[6]},
      {stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1],stage5_0[1]}
   );
   gpc2135_5 gpc5559 (
      {stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5], stage4_3[6]},
      {stage4_4[0], stage4_4[1], stage4_4[2]},
      {stage4_5[0]},
      {stage4_6[0], stage4_6[1]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[2],stage5_3[2]}
   );
   gpc615_5 gpc5560 (
      {stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage4_4[3]},
      {stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6]},
      {stage5_7[1],stage5_6[1],stage5_5[1],stage5_4[3],stage5_3[3]}
   );
   gpc615_5 gpc5561 (
      {stage4_3[12], stage4_3[13], stage4_3[14], stage4_3[15], stage4_3[16]},
      {stage4_4[4]},
      {stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11], stage4_5[12]},
      {stage5_7[2],stage5_6[2],stage5_5[2],stage5_4[4],stage5_3[4]}
   );
   gpc1163_5 gpc5562 (
      {stage4_5[13], stage4_5[14], stage4_5[15]},
      {stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5], stage4_6[6], stage4_6[7]},
      {stage4_7[0]},
      {stage4_8[0]},
      {stage5_9[0],stage5_8[0],stage5_7[3],stage5_6[3],stage5_5[3]}
   );
   gpc117_4 gpc5563 (
      {stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5], stage4_7[6], stage4_7[7]},
      {stage4_8[1]},
      {stage4_9[0]},
      {stage5_10[0],stage5_9[1],stage5_8[1],stage5_7[4]}
   );
   gpc117_4 gpc5564 (
      {stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5], stage4_8[6], stage4_8[7], stage4_8[8]},
      {stage4_9[1]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[1],stage5_9[2],stage5_8[2]}
   );
   gpc117_4 gpc5565 (
      {stage4_8[9], stage4_8[10], stage4_8[11], stage4_8[12], stage4_8[13], stage4_8[14], stage4_8[15]},
      {stage4_9[2]},
      {stage4_10[1]},
      {stage5_11[1],stage5_10[2],stage5_9[3],stage5_8[3]}
   );
   gpc606_5 gpc5566 (
      {stage4_8[16], stage4_8[17], stage4_8[18], stage4_8[19], stage4_8[20], stage4_8[21]},
      {stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage5_12[0],stage5_11[2],stage5_10[3],stage5_9[4],stage5_8[4]}
   );
   gpc615_5 gpc5567 (
      {stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11], stage4_10[12]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[0],stage5_12[1],stage5_11[3],stage5_10[4]}
   );
   gpc606_5 gpc5568 (
      {stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage5_15[0],stage5_14[1],stage5_13[1],stage5_12[2],stage5_11[4]}
   );
   gpc606_5 gpc5569 (
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[1],stage5_14[2],stage5_13[2],stage5_12[3]}
   );
   gpc615_5 gpc5570 (
      {stage4_12[12], stage4_12[13], stage4_12[14], stage4_12[15], stage4_12[16]},
      {stage4_13[6]},
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10], stage4_14[11]},
      {stage5_16[1],stage5_15[2],stage5_14[3],stage5_13[3],stage5_12[4]}
   );
   gpc606_5 gpc5571 (
      {stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[2],stage5_15[3],stage5_14[4],stage5_13[4]}
   );
   gpc615_5 gpc5572 (
      {stage4_15[6], stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10]},
      {stage4_16[0]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[0],stage5_17[1],stage5_16[3],stage5_15[4]}
   );
   gpc207_4 gpc5573 (
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5], stage4_16[6], stage4_16[7]},
      {stage4_18[0], stage4_18[1]},
      {stage5_19[1],stage5_18[1],stage5_17[2],stage5_16[4]}
   );
   gpc207_4 gpc5574 (
      {stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11], stage4_16[12], 1'b0, 1'b0},
      {stage4_18[2], stage4_18[3]},
      {stage5_19[2],stage5_18[2],stage5_17[3],stage5_16[5]}
   );
   gpc606_5 gpc5575 (
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[0],stage5_19[3],stage5_18[3],stage5_17[4]}
   );
   gpc615_5 gpc5576 (
      {stage4_18[4], stage4_18[5], stage4_18[6], stage4_18[7], stage4_18[8]},
      {stage4_19[6]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[1],stage5_20[1],stage5_19[4],stage5_18[4]}
   );
   gpc623_5 gpc5577 (
      {stage4_18[9], stage4_18[10], 1'b0},
      {stage4_19[7], stage4_19[8]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], 1'b0},
      {stage5_22[1],stage5_21[2],stage5_20[2],stage5_19[5],stage5_18[5]}
   );
   gpc135_4 gpc5578 (
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4]},
      {stage4_23[0], stage4_23[1], stage4_23[2]},
      {stage4_24[0]},
      {stage5_25[0],stage5_24[0],stage5_23[0],stage5_22[2]}
   );
   gpc2135_5 gpc5579 (
      {stage4_22[5], stage4_22[6], stage4_22[7], stage4_22[8], stage4_22[9]},
      {stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[1]},
      {stage4_25[0], stage4_25[1]},
      {stage5_26[0],stage5_25[1],stage5_24[1],stage5_23[1],stage5_22[3]}
   );
   gpc2135_5 gpc5580 (
      {stage4_22[10], stage4_22[11], stage4_22[12], stage4_22[13], stage4_22[14]},
      {stage4_23[6], stage4_23[7], stage4_23[8]},
      {stage4_24[2]},
      {stage4_25[2], stage4_25[3]},
      {stage5_26[1],stage5_25[2],stage5_24[2],stage5_23[2],stage5_22[4]}
   );
   gpc606_5 gpc5581 (
      {stage4_24[3], stage4_24[4], stage4_24[5], stage4_24[6], stage4_24[7], stage4_24[8]},
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5]},
      {stage5_28[0],stage5_27[0],stage5_26[2],stage5_25[3],stage5_24[3]}
   );
   gpc23_3 gpc5582 (
      {stage4_25[4], stage4_25[5], stage4_25[6]},
      {stage4_26[6], stage4_26[7]},
      {stage5_27[1],stage5_26[3],stage5_25[4]}
   );
   gpc7_3 gpc5583 (
      {stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11], stage4_25[12], stage4_25[13]},
      {stage5_27[2],stage5_26[4],stage5_25[5]}
   );
   gpc615_5 gpc5584 (
      {stage4_26[8], stage4_26[9], stage4_26[10], stage4_26[11], stage4_26[12]},
      {stage4_27[0]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[3],stage5_26[5]}
   );
   gpc1343_5 gpc5585 (
      {stage4_27[1], stage4_27[2], stage4_27[3]},
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9]},
      {stage4_29[0], stage4_29[1], stage4_29[2]},
      {stage4_30[0]},
      {stage5_31[0],stage5_30[1],stage5_29[1],stage5_28[2],stage5_27[4]}
   );
   gpc1423_5 gpc5586 (
      {stage4_27[4], stage4_27[5], stage4_27[6]},
      {stage4_28[10], stage4_28[11]},
      {stage4_29[3], stage4_29[4], stage4_29[5], stage4_29[6]},
      {stage4_30[1]},
      {stage5_31[1],stage5_30[2],stage5_29[2],stage5_28[3],stage5_27[5]}
   );
   gpc606_5 gpc5587 (
      {stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10], stage4_29[11], stage4_29[12]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[2],stage5_30[3],stage5_29[3]}
   );
   gpc615_5 gpc5588 (
      {stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5], stage4_30[6]},
      {stage4_31[6]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[1],stage5_32[1],stage5_31[3],stage5_30[4]}
   );
   gpc615_5 gpc5589 (
      {stage4_30[7], stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11]},
      {stage4_31[7]},
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11]},
      {stage5_34[1],stage5_33[2],stage5_32[2],stage5_31[4],stage5_30[5]}
   );
   gpc606_5 gpc5590 (
      {stage4_32[12], stage4_32[13], stage4_32[14], stage4_32[15], stage4_32[16], stage4_32[17]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[0],stage5_34[2],stage5_33[3],stage5_32[3]}
   );
   gpc606_5 gpc5591 (
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[1],stage5_35[1],stage5_34[3],stage5_33[4]}
   );
   gpc606_5 gpc5592 (
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10], stage4_35[11]},
      {stage5_37[1],stage5_36[2],stage5_35[2],stage5_34[4],stage5_33[5]}
   );
   gpc606_5 gpc5593 (
      {stage4_33[12], stage4_33[13], stage4_33[14], stage4_33[15], stage4_33[16], 1'b0},
      {stage4_35[12], stage4_35[13], stage4_35[14], stage4_35[15], stage4_35[16], 1'b0},
      {stage5_37[2],stage5_36[3],stage5_35[3],stage5_34[5],stage5_33[6]}
   );
   gpc615_5 gpc5594 (
      {stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9], stage4_34[10]},
      {1'b0},
      {stage4_36[0], stage4_36[1], stage4_36[2], stage4_36[3], stage4_36[4], stage4_36[5]},
      {stage5_38[0],stage5_37[3],stage5_36[4],stage5_35[4],stage5_34[6]}
   );
   gpc606_5 gpc5595 (
      {stage4_36[6], stage4_36[7], stage4_36[8], stage4_36[9], stage4_36[10], stage4_36[11]},
      {stage4_38[0], stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4], stage4_38[5]},
      {stage5_40[0],stage5_39[0],stage5_38[1],stage5_37[4],stage5_36[5]}
   );
   gpc606_5 gpc5596 (
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage4_39[0], stage4_39[1], stage4_39[2], stage4_39[3], stage4_39[4], stage4_39[5]},
      {stage5_41[0],stage5_40[1],stage5_39[1],stage5_38[2],stage5_37[5]}
   );
   gpc606_5 gpc5597 (
      {stage4_39[6], stage4_39[7], stage4_39[8], 1'b0, 1'b0, 1'b0},
      {stage4_41[0], stage4_41[1], stage4_41[2], stage4_41[3], stage4_41[4], stage4_41[5]},
      {stage5_43[0],stage5_42[0],stage5_41[1],stage5_40[2],stage5_39[2]}
   );
   gpc606_5 gpc5598 (
      {stage4_40[0], stage4_40[1], stage4_40[2], stage4_40[3], stage4_40[4], stage4_40[5]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[1],stage5_42[1],stage5_41[2],stage5_40[3]}
   );
   gpc606_5 gpc5599 (
      {stage4_40[6], stage4_40[7], stage4_40[8], stage4_40[9], stage4_40[10], stage4_40[11]},
      {stage4_42[6], stage4_42[7], stage4_42[8], stage4_42[9], stage4_42[10], stage4_42[11]},
      {stage5_44[1],stage5_43[2],stage5_42[2],stage5_41[3],stage5_40[4]}
   );
   gpc606_5 gpc5600 (
      {stage4_41[6], stage4_41[7], stage4_41[8], stage4_41[9], stage4_41[10], stage4_41[11]},
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], stage4_43[5]},
      {stage5_45[0],stage5_44[2],stage5_43[3],stage5_42[3],stage5_41[4]}
   );
   gpc615_5 gpc5601 (
      {stage4_43[6], stage4_43[7], stage4_43[8], stage4_43[9], stage4_43[10]},
      {stage4_44[0]},
      {stage4_45[0], stage4_45[1], stage4_45[2], stage4_45[3], stage4_45[4], stage4_45[5]},
      {stage5_47[0],stage5_46[0],stage5_45[1],stage5_44[3],stage5_43[4]}
   );
   gpc615_5 gpc5602 (
      {stage4_43[11], stage4_43[12], stage4_43[13], stage4_43[14], stage4_43[15]},
      {stage4_44[1]},
      {stage4_45[6], stage4_45[7], stage4_45[8], stage4_45[9], stage4_45[10], stage4_45[11]},
      {stage5_47[1],stage5_46[1],stage5_45[2],stage5_44[4],stage5_43[5]}
   );
   gpc606_5 gpc5603 (
      {stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5], stage4_44[6], stage4_44[7]},
      {stage4_46[0], stage4_46[1], stage4_46[2], stage4_46[3], stage4_46[4], stage4_46[5]},
      {stage5_48[0],stage5_47[2],stage5_46[2],stage5_45[3],stage5_44[5]}
   );
   gpc606_5 gpc5604 (
      {stage4_44[8], stage4_44[9], stage4_44[10], stage4_44[11], stage4_44[12], stage4_44[13]},
      {stage4_46[6], stage4_46[7], stage4_46[8], stage4_46[9], stage4_46[10], stage4_46[11]},
      {stage5_48[1],stage5_47[3],stage5_46[3],stage5_45[4],stage5_44[6]}
   );
   gpc615_5 gpc5605 (
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4]},
      {stage4_48[0]},
      {stage4_49[0], stage4_49[1], stage4_49[2], stage4_49[3], stage4_49[4], stage4_49[5]},
      {stage5_51[0],stage5_50[0],stage5_49[0],stage5_48[2],stage5_47[4]}
   );
   gpc615_5 gpc5606 (
      {stage4_47[5], stage4_47[6], stage4_47[7], stage4_47[8], stage4_47[9]},
      {stage4_48[1]},
      {stage4_49[6], stage4_49[7], stage4_49[8], stage4_49[9], stage4_49[10], stage4_49[11]},
      {stage5_51[1],stage5_50[1],stage5_49[1],stage5_48[3],stage5_47[5]}
   );
   gpc615_5 gpc5607 (
      {stage4_47[10], stage4_47[11], stage4_47[12], stage4_47[13], stage4_47[14]},
      {stage4_48[2]},
      {stage4_49[12], stage4_49[13], stage4_49[14], stage4_49[15], stage4_49[16], stage4_49[17]},
      {stage5_51[2],stage5_50[2],stage5_49[2],stage5_48[4],stage5_47[6]}
   );
   gpc606_5 gpc5608 (
      {stage4_48[3], stage4_48[4], stage4_48[5], stage4_48[6], stage4_48[7], stage4_48[8]},
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], stage4_50[4], stage4_50[5]},
      {stage5_52[0],stage5_51[3],stage5_50[3],stage5_49[3],stage5_48[5]}
   );
   gpc606_5 gpc5609 (
      {stage4_48[9], stage4_48[10], stage4_48[11], stage4_48[12], stage4_48[13], stage4_48[14]},
      {stage4_50[6], stage4_50[7], stage4_50[8], stage4_50[9], stage4_50[10], stage4_50[11]},
      {stage5_52[1],stage5_51[4],stage5_50[4],stage5_49[4],stage5_48[6]}
   );
   gpc606_5 gpc5610 (
      {stage4_49[18], stage4_49[19], stage4_49[20], stage4_49[21], stage4_49[22], stage4_49[23]},
      {stage4_51[0], stage4_51[1], stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5]},
      {stage5_53[0],stage5_52[2],stage5_51[5],stage5_50[5],stage5_49[5]}
   );
   gpc606_5 gpc5611 (
      {stage4_49[24], stage4_49[25], stage4_49[26], stage4_49[27], stage4_49[28], stage4_49[29]},
      {stage4_51[6], stage4_51[7], stage4_51[8], stage4_51[9], stage4_51[10], stage4_51[11]},
      {stage5_53[1],stage5_52[3],stage5_51[6],stage5_50[6],stage5_49[6]}
   );
   gpc606_5 gpc5612 (
      {stage4_49[30], stage4_49[31], stage4_49[32], stage4_49[33], stage4_49[34], stage4_49[35]},
      {stage4_51[12], stage4_51[13], stage4_51[14], stage4_51[15], stage4_51[16], stage4_51[17]},
      {stage5_53[2],stage5_52[4],stage5_51[7],stage5_50[7],stage5_49[7]}
   );
   gpc615_5 gpc5613 (
      {stage4_50[12], stage4_50[13], stage4_50[14], stage4_50[15], stage4_50[16]},
      {stage4_51[18]},
      {stage4_52[0], stage4_52[1], stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5]},
      {stage5_54[0],stage5_53[3],stage5_52[5],stage5_51[8],stage5_50[8]}
   );
   gpc7_3 gpc5614 (
      {stage4_52[6], stage4_52[7], stage4_52[8], stage4_52[9], stage4_52[10], stage4_52[11], stage4_52[12]},
      {stage5_54[1],stage5_53[4],stage5_52[6]}
   );
   gpc606_5 gpc5615 (
      {stage4_53[0], stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5]},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5]},
      {stage5_57[0],stage5_56[0],stage5_55[0],stage5_54[2],stage5_53[5]}
   );
   gpc207_4 gpc5616 (
      {stage4_54[0], stage4_54[1], stage4_54[2], stage4_54[3], stage4_54[4], stage4_54[5], stage4_54[6]},
      {stage4_56[0], stage4_56[1]},
      {stage5_57[1],stage5_56[1],stage5_55[1],stage5_54[3]}
   );
   gpc207_4 gpc5617 (
      {stage4_54[7], stage4_54[8], stage4_54[9], stage4_54[10], stage4_54[11], stage4_54[12], stage4_54[13]},
      {stage4_56[2], stage4_56[3]},
      {stage5_57[2],stage5_56[2],stage5_55[2],stage5_54[4]}
   );
   gpc207_4 gpc5618 (
      {stage4_54[14], stage4_54[15], stage4_54[16], stage4_54[17], 1'b0, 1'b0, 1'b0},
      {stage4_56[4], stage4_56[5]},
      {stage5_57[3],stage5_56[3],stage5_55[3],stage5_54[5]}
   );
   gpc606_5 gpc5619 (
      {stage4_55[6], stage4_55[7], stage4_55[8], stage4_55[9], stage4_55[10], stage4_55[11]},
      {stage4_57[0], stage4_57[1], stage4_57[2], stage4_57[3], stage4_57[4], stage4_57[5]},
      {stage5_59[0],stage5_58[0],stage5_57[4],stage5_56[4],stage5_55[4]}
   );
   gpc606_5 gpc5620 (
      {stage4_56[6], stage4_56[7], stage4_56[8], stage4_56[9], stage4_56[10], stage4_56[11]},
      {stage4_58[0], stage4_58[1], stage4_58[2], stage4_58[3], stage4_58[4], stage4_58[5]},
      {stage5_60[0],stage5_59[1],stage5_58[1],stage5_57[5],stage5_56[5]}
   );
   gpc7_3 gpc5621 (
      {stage4_57[6], stage4_57[7], stage4_57[8], stage4_57[9], stage4_57[10], stage4_57[11], 1'b0},
      {stage5_59[2],stage5_58[2],stage5_57[6]}
   );
   gpc7_3 gpc5622 (
      {stage4_58[6], stage4_58[7], stage4_58[8], stage4_58[9], stage4_58[10], stage4_58[11], stage4_58[12]},
      {stage5_60[1],stage5_59[3],stage5_58[3]}
   );
   gpc7_3 gpc5623 (
      {stage4_58[13], stage4_58[14], stage4_58[15], stage4_58[16], stage4_58[17], stage4_58[18], stage4_58[19]},
      {stage5_60[2],stage5_59[4],stage5_58[4]}
   );
   gpc606_5 gpc5624 (
      {stage4_59[0], stage4_59[1], stage4_59[2], stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[0],stage5_61[0],stage5_60[3],stage5_59[5]}
   );
   gpc606_5 gpc5625 (
      {stage4_59[6], stage4_59[7], stage4_59[8], stage4_59[9], stage4_59[10], stage4_59[11]},
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], stage4_61[10], stage4_61[11]},
      {stage5_63[1],stage5_62[1],stage5_61[1],stage5_60[4],stage5_59[6]}
   );
   gpc606_5 gpc5626 (
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[2],stage5_62[2],stage5_61[2],stage5_60[5]}
   );
   gpc606_5 gpc5627 (
      {stage4_60[6], stage4_60[7], stage4_60[8], stage4_60[9], stage4_60[10], stage4_60[11]},
      {stage4_62[6], stage4_62[7], stage4_62[8], stage4_62[9], stage4_62[10], stage4_62[11]},
      {stage5_64[1],stage5_63[3],stage5_62[3],stage5_61[3],stage5_60[6]}
   );
   gpc117_4 gpc5628 (
      {stage4_63[0], stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4], stage4_63[5], stage4_63[6]},
      {stage4_64[0]},
      {stage4_65[0]},
      {stage5_66[0],stage5_65[0],stage5_64[2],stage5_63[4]}
   );
   gpc117_4 gpc5629 (
      {stage4_63[7], stage4_63[8], stage4_63[9], stage4_63[10], stage4_63[11], stage4_63[12], 1'b0},
      {stage4_64[1]},
      {stage4_65[1]},
      {stage5_66[1],stage5_65[1],stage5_64[3],stage5_63[5]}
   );
   gpc606_5 gpc5630 (
      {stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5], stage4_64[6], stage4_64[7]},
      {stage4_66[0], stage4_66[1], stage4_66[2], stage4_66[3], stage4_66[4], stage4_66[5]},
      {stage5_68[0],stage5_67[0],stage5_66[2],stage5_65[2],stage5_64[4]}
   );
   gpc606_5 gpc5631 (
      {stage4_64[8], stage4_64[9], stage4_64[10], stage4_64[11], 1'b0, 1'b0},
      {stage4_66[6], stage4_66[7], stage4_66[8], stage4_66[9], stage4_66[10], stage4_66[11]},
      {stage5_68[1],stage5_67[1],stage5_66[3],stage5_65[3],stage5_64[5]}
   );
   gpc606_5 gpc5632 (
      {stage4_65[2], stage4_65[3], stage4_65[4], stage4_65[5], stage4_65[6], stage4_65[7]},
      {stage4_67[0], stage4_67[1], stage4_67[2], stage4_67[3], stage4_67[4], stage4_67[5]},
      {stage5_69[0],stage5_68[2],stage5_67[2],stage5_66[4],stage5_65[4]}
   );
   gpc207_4 gpc5633 (
      {stage4_66[12], stage4_66[13], stage4_66[14], stage4_66[15], stage4_66[16], stage4_66[17], stage4_66[18]},
      {stage4_68[0], stage4_68[1]},
      {stage5_69[1],stage5_68[3],stage5_67[3],stage5_66[5]}
   );
   gpc1_1 gpc5634 (
      {stage4_0[11]},
      {stage5_0[2]}
   );
   gpc1_1 gpc5635 (
      {stage4_0[12]},
      {stage5_0[3]}
   );
   gpc1_1 gpc5636 (
      {stage4_0[13]},
      {stage5_0[4]}
   );
   gpc1_1 gpc5637 (
      {stage4_1[3]},
      {stage5_1[2]}
   );
   gpc1_1 gpc5638 (
      {stage4_1[4]},
      {stage5_1[3]}
   );
   gpc1_1 gpc5639 (
      {stage4_3[17]},
      {stage5_3[5]}
   );
   gpc1_1 gpc5640 (
      {stage4_3[18]},
      {stage5_3[6]}
   );
   gpc1_1 gpc5641 (
      {stage4_4[5]},
      {stage5_4[5]}
   );
   gpc1_1 gpc5642 (
      {stage4_4[6]},
      {stage5_4[6]}
   );
   gpc1_1 gpc5643 (
      {stage4_4[7]},
      {stage5_4[7]}
   );
   gpc1_1 gpc5644 (
      {stage4_4[8]},
      {stage5_4[8]}
   );
   gpc1_1 gpc5645 (
      {stage4_4[9]},
      {stage5_4[9]}
   );
   gpc1_1 gpc5646 (
      {stage4_5[16]},
      {stage5_5[4]}
   );
   gpc1_1 gpc5647 (
      {stage4_5[17]},
      {stage5_5[5]}
   );
   gpc1_1 gpc5648 (
      {stage4_5[18]},
      {stage5_5[6]}
   );
   gpc1_1 gpc5649 (
      {stage4_5[19]},
      {stage5_5[7]}
   );
   gpc1_1 gpc5650 (
      {stage4_6[8]},
      {stage5_6[4]}
   );
   gpc1_1 gpc5651 (
      {stage4_6[9]},
      {stage5_6[5]}
   );
   gpc1_1 gpc5652 (
      {stage4_7[8]},
      {stage5_7[5]}
   );
   gpc1_1 gpc5653 (
      {stage4_7[9]},
      {stage5_7[6]}
   );
   gpc1_1 gpc5654 (
      {stage4_9[3]},
      {stage5_9[5]}
   );
   gpc1_1 gpc5655 (
      {stage4_9[4]},
      {stage5_9[6]}
   );
   gpc1_1 gpc5656 (
      {stage4_9[5]},
      {stage5_9[7]}
   );
   gpc1_1 gpc5657 (
      {stage4_9[6]},
      {stage5_9[8]}
   );
   gpc1_1 gpc5658 (
      {stage4_9[7]},
      {stage5_9[9]}
   );
   gpc1_1 gpc5659 (
      {stage4_10[13]},
      {stage5_10[5]}
   );
   gpc1_1 gpc5660 (
      {stage4_11[7]},
      {stage5_11[5]}
   );
   gpc1_1 gpc5661 (
      {stage4_11[8]},
      {stage5_11[6]}
   );
   gpc1_1 gpc5662 (
      {stage4_11[9]},
      {stage5_11[7]}
   );
   gpc1_1 gpc5663 (
      {stage4_11[10]},
      {stage5_11[8]}
   );
   gpc1_1 gpc5664 (
      {stage4_11[11]},
      {stage5_11[9]}
   );
   gpc1_1 gpc5665 (
      {stage4_12[17]},
      {stage5_12[5]}
   );
   gpc1_1 gpc5666 (
      {stage4_13[13]},
      {stage5_13[5]}
   );
   gpc1_1 gpc5667 (
      {stage4_15[11]},
      {stage5_15[5]}
   );
   gpc1_1 gpc5668 (
      {stage4_17[12]},
      {stage5_17[5]}
   );
   gpc1_1 gpc5669 (
      {stage4_17[13]},
      {stage5_17[6]}
   );
   gpc1_1 gpc5670 (
      {stage4_17[14]},
      {stage5_17[7]}
   );
   gpc1_1 gpc5671 (
      {stage4_19[9]},
      {stage5_19[6]}
   );
   gpc1_1 gpc5672 (
      {stage4_19[10]},
      {stage5_19[7]}
   );
   gpc1_1 gpc5673 (
      {stage4_19[11]},
      {stage5_19[8]}
   );
   gpc1_1 gpc5674 (
      {stage4_19[12]},
      {stage5_19[9]}
   );
   gpc1_1 gpc5675 (
      {stage4_19[13]},
      {stage5_19[10]}
   );
   gpc1_1 gpc5676 (
      {stage4_21[0]},
      {stage5_21[3]}
   );
   gpc1_1 gpc5677 (
      {stage4_21[1]},
      {stage5_21[4]}
   );
   gpc1_1 gpc5678 (
      {stage4_21[2]},
      {stage5_21[5]}
   );
   gpc1_1 gpc5679 (
      {stage4_21[3]},
      {stage5_21[6]}
   );
   gpc1_1 gpc5680 (
      {stage4_21[4]},
      {stage5_21[7]}
   );
   gpc1_1 gpc5681 (
      {stage4_21[5]},
      {stage5_21[8]}
   );
   gpc1_1 gpc5682 (
      {stage4_21[6]},
      {stage5_21[9]}
   );
   gpc1_1 gpc5683 (
      {stage4_21[7]},
      {stage5_21[10]}
   );
   gpc1_1 gpc5684 (
      {stage4_21[8]},
      {stage5_21[11]}
   );
   gpc1_1 gpc5685 (
      {stage4_24[9]},
      {stage5_24[4]}
   );
   gpc1_1 gpc5686 (
      {stage4_24[10]},
      {stage5_24[5]}
   );
   gpc1_1 gpc5687 (
      {stage4_24[11]},
      {stage5_24[6]}
   );
   gpc1_1 gpc5688 (
      {stage4_29[13]},
      {stage5_29[4]}
   );
   gpc1_1 gpc5689 (
      {stage4_29[14]},
      {stage5_29[5]}
   );
   gpc1_1 gpc5690 (
      {stage4_29[15]},
      {stage5_29[6]}
   );
   gpc1_1 gpc5691 (
      {stage4_29[16]},
      {stage5_29[7]}
   );
   gpc1_1 gpc5692 (
      {stage4_31[8]},
      {stage5_31[5]}
   );
   gpc1_1 gpc5693 (
      {stage4_31[9]},
      {stage5_31[6]}
   );
   gpc1_1 gpc5694 (
      {stage4_36[12]},
      {stage5_36[6]}
   );
   gpc1_1 gpc5695 (
      {stage4_37[6]},
      {stage5_37[6]}
   );
   gpc1_1 gpc5696 (
      {stage4_37[7]},
      {stage5_37[7]}
   );
   gpc1_1 gpc5697 (
      {stage4_37[8]},
      {stage5_37[8]}
   );
   gpc1_1 gpc5698 (
      {stage4_37[9]},
      {stage5_37[9]}
   );
   gpc1_1 gpc5699 (
      {stage4_37[10]},
      {stage5_37[10]}
   );
   gpc1_1 gpc5700 (
      {stage4_37[11]},
      {stage5_37[11]}
   );
   gpc1_1 gpc5701 (
      {stage4_38[6]},
      {stage5_38[3]}
   );
   gpc1_1 gpc5702 (
      {stage4_40[12]},
      {stage5_40[5]}
   );
   gpc1_1 gpc5703 (
      {stage4_42[12]},
      {stage5_42[4]}
   );
   gpc1_1 gpc5704 (
      {stage4_42[13]},
      {stage5_42[5]}
   );
   gpc1_1 gpc5705 (
      {stage4_42[14]},
      {stage5_42[6]}
   );
   gpc1_1 gpc5706 (
      {stage4_43[16]},
      {stage5_43[6]}
   );
   gpc1_1 gpc5707 (
      {stage4_43[17]},
      {stage5_43[7]}
   );
   gpc1_1 gpc5708 (
      {stage4_43[18]},
      {stage5_43[8]}
   );
   gpc1_1 gpc5709 (
      {stage4_43[19]},
      {stage5_43[9]}
   );
   gpc1_1 gpc5710 (
      {stage4_46[12]},
      {stage5_46[4]}
   );
   gpc1_1 gpc5711 (
      {stage4_46[13]},
      {stage5_46[5]}
   );
   gpc1_1 gpc5712 (
      {stage4_46[14]},
      {stage5_46[6]}
   );
   gpc1_1 gpc5713 (
      {stage4_51[19]},
      {stage5_51[9]}
   );
   gpc1_1 gpc5714 (
      {stage4_52[13]},
      {stage5_52[7]}
   );
   gpc1_1 gpc5715 (
      {stage4_53[6]},
      {stage5_53[6]}
   );
   gpc1_1 gpc5716 (
      {stage4_53[7]},
      {stage5_53[7]}
   );
   gpc1_1 gpc5717 (
      {stage4_53[8]},
      {stage5_53[8]}
   );
   gpc1_1 gpc5718 (
      {stage4_53[9]},
      {stage5_53[9]}
   );
   gpc1_1 gpc5719 (
      {stage4_53[10]},
      {stage5_53[10]}
   );
   gpc1_1 gpc5720 (
      {stage4_53[11]},
      {stage5_53[11]}
   );
   gpc1_1 gpc5721 (
      {stage4_53[12]},
      {stage5_53[12]}
   );
   gpc1_1 gpc5722 (
      {stage4_53[13]},
      {stage5_53[13]}
   );
   gpc1_1 gpc5723 (
      {stage4_53[14]},
      {stage5_53[14]}
   );
   gpc1_1 gpc5724 (
      {stage4_55[12]},
      {stage5_55[5]}
   );
   gpc1_1 gpc5725 (
      {stage4_60[12]},
      {stage5_60[7]}
   );
   gpc1_1 gpc5726 (
      {stage4_60[13]},
      {stage5_60[8]}
   );
   gpc1_1 gpc5727 (
      {stage4_66[19]},
      {stage5_66[6]}
   );
   gpc1_1 gpc5728 (
      {stage4_66[20]},
      {stage5_66[7]}
   );
   gpc1_1 gpc5729 (
      {stage4_66[21]},
      {stage5_66[8]}
   );
   gpc1_1 gpc5730 (
      {stage4_66[22]},
      {stage5_66[9]}
   );
   gpc1_1 gpc5731 (
      {stage4_66[23]},
      {stage5_66[10]}
   );
   gpc1_1 gpc5732 (
      {stage4_67[6]},
      {stage5_67[4]}
   );
   gpc1_1 gpc5733 (
      {stage4_67[7]},
      {stage5_67[5]}
   );
   gpc1_1 gpc5734 (
      {stage4_67[8]},
      {stage5_67[6]}
   );
   gpc1_1 gpc5735 (
      {stage4_68[2]},
      {stage5_68[4]}
   );
   gpc1_1 gpc5736 (
      {stage4_69[0]},
      {stage5_69[2]}
   );
   gpc223_4 gpc5737 (
      {stage5_2[0], stage5_2[1], 1'b0},
      {stage5_3[0], stage5_3[1]},
      {stage5_4[0], stage5_4[1]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc615_5 gpc5738 (
      {stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5], stage5_3[6]},
      {stage5_4[2]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc615_5 gpc5739 (
      {stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6], stage5_4[7]},
      {stage5_5[6]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5]},
      {stage6_8[0],stage6_7[1],stage6_6[1],stage6_5[2],stage6_4[2]}
   );
   gpc207_4 gpc5740 (
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5], stage5_7[6]},
      {stage5_9[0], stage5_9[1]},
      {stage6_10[0],stage6_9[0],stage6_8[1],stage6_7[2]}
   );
   gpc615_5 gpc5741 (
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4]},
      {stage5_9[2]},
      {stage5_10[0], stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage6_12[0],stage6_11[0],stage6_10[1],stage6_9[1],stage6_8[2]}
   );
   gpc606_5 gpc5742 (
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc7_3 gpc5743 (
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], 1'b0},
      {stage6_14[1],stage6_13[1],stage6_12[2]}
   );
   gpc615_5 gpc5744 (
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4]},
      {stage5_16[0]},
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage6_19[0],stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[1]}
   );
   gpc1415_5 gpc5745 (
      {stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage5_17[6]},
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3]},
      {stage5_19[0]},
      {stage6_20[0],stage6_19[1],stage6_18[1],stage6_17[1],stage6_16[1]}
   );
   gpc615_5 gpc5746 (
      {stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage5_20[0]},
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage6_23[0],stage6_22[0],stage6_21[0],stage6_20[1],stage6_19[2]}
   );
   gpc615_5 gpc5747 (
      {stage5_19[6], stage5_19[7], stage5_19[8], stage5_19[9], stage5_19[10]},
      {stage5_20[1]},
      {stage5_21[6], stage5_21[7], stage5_21[8], stage5_21[9], stage5_21[10], stage5_21[11]},
      {stage6_23[1],stage6_22[1],stage6_21[1],stage6_20[2],stage6_19[3]}
   );
   gpc615_5 gpc5748 (
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4]},
      {stage5_23[0]},
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5]},
      {stage6_26[0],stage6_25[0],stage6_24[0],stage6_23[2],stage6_22[2]}
   );
   gpc207_4 gpc5749 (
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5], 1'b0},
      {stage5_28[0], stage5_28[1]},
      {stage6_29[0],stage6_28[0],stage6_27[0],stage6_26[1]}
   );
   gpc1325_5 gpc5750 (
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3], stage5_27[4]},
      {stage5_28[2], stage5_28[3]},
      {stage5_29[0], stage5_29[1], stage5_29[2]},
      {stage5_30[0]},
      {stage6_31[0],stage6_30[0],stage6_29[1],stage6_28[1],stage6_27[1]}
   );
   gpc615_5 gpc5751 (
      {stage5_29[3], stage5_29[4], stage5_29[5], stage5_29[6], stage5_29[7]},
      {stage5_30[1]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[0],stage6_31[1],stage6_30[1],stage6_29[2]}
   );
   gpc2135_5 gpc5752 (
      {stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5], 1'b0},
      {stage5_31[6], 1'b0, 1'b0},
      {stage5_32[0]},
      {stage5_33[0], stage5_33[1]},
      {stage6_34[0],stage6_33[1],stage6_32[1],stage6_31[2],stage6_30[2]}
   );
   gpc615_5 gpc5753 (
      {stage5_32[1], stage5_32[2], stage5_32[3], 1'b0, 1'b0},
      {stage5_33[2]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5]},
      {stage6_36[0],stage6_35[0],stage6_34[1],stage6_33[2],stage6_32[2]}
   );
   gpc117_4 gpc5754 (
      {stage5_33[3], stage5_33[4], stage5_33[5], stage5_33[6], 1'b0, 1'b0, 1'b0},
      {stage5_34[6]},
      {stage5_35[0]},
      {stage6_36[1],stage6_35[1],stage6_34[2],stage6_33[3]}
   );
   gpc623_5 gpc5755 (
      {stage5_35[1], stage5_35[2], stage5_35[3]},
      {stage5_36[0], stage5_36[1]},
      {stage5_37[0], stage5_37[1], stage5_37[2], stage5_37[3], stage5_37[4], stage5_37[5]},
      {stage6_39[0],stage6_38[0],stage6_37[0],stage6_36[2],stage6_35[2]}
   );
   gpc606_5 gpc5756 (
      {stage5_36[2], stage5_36[3], stage5_36[4], stage5_36[5], stage5_36[6], 1'b0},
      {stage5_38[0], stage5_38[1], stage5_38[2], stage5_38[3], 1'b0, 1'b0},
      {stage6_40[0],stage6_39[1],stage6_38[1],stage6_37[1],stage6_36[3]}
   );
   gpc1163_5 gpc5757 (
      {stage5_39[0], stage5_39[1], stage5_39[2]},
      {stage5_40[0], stage5_40[1], stage5_40[2], stage5_40[3], stage5_40[4], stage5_40[5]},
      {stage5_41[0]},
      {stage5_42[0]},
      {stage6_43[0],stage6_42[0],stage6_41[0],stage6_40[1],stage6_39[2]}
   );
   gpc1415_5 gpc5758 (
      {stage5_41[1], stage5_41[2], stage5_41[3], stage5_41[4], 1'b0},
      {stage5_42[1]},
      {stage5_43[0], stage5_43[1], stage5_43[2], stage5_43[3]},
      {stage5_44[0]},
      {stage6_45[0],stage6_44[0],stage6_43[1],stage6_42[1],stage6_41[1]}
   );
   gpc135_4 gpc5759 (
      {stage5_42[2], stage5_42[3], stage5_42[4], stage5_42[5], stage5_42[6]},
      {stage5_43[4], stage5_43[5], stage5_43[6]},
      {stage5_44[1]},
      {stage6_45[1],stage6_44[1],stage6_43[2],stage6_42[2]}
   );
   gpc606_5 gpc5760 (
      {stage5_44[2], stage5_44[3], stage5_44[4], stage5_44[5], stage5_44[6], 1'b0},
      {stage5_46[0], stage5_46[1], stage5_46[2], stage5_46[3], stage5_46[4], stage5_46[5]},
      {stage6_48[0],stage6_47[0],stage6_46[0],stage6_45[2],stage6_44[2]}
   );
   gpc2135_5 gpc5761 (
      {stage5_45[0], stage5_45[1], stage5_45[2], stage5_45[3], stage5_45[4]},
      {stage5_46[6], 1'b0, 1'b0},
      {stage5_47[0]},
      {stage5_48[0], stage5_48[1]},
      {stage6_49[0],stage6_48[1],stage6_47[1],stage6_46[1],stage6_45[3]}
   );
   gpc623_5 gpc5762 (
      {stage5_47[1], stage5_47[2], stage5_47[3]},
      {stage5_48[2], stage5_48[3]},
      {stage5_49[0], stage5_49[1], stage5_49[2], stage5_49[3], stage5_49[4], stage5_49[5]},
      {stage6_51[0],stage6_50[0],stage6_49[1],stage6_48[2],stage6_47[2]}
   );
   gpc223_4 gpc5763 (
      {stage5_48[4], stage5_48[5], stage5_48[6]},
      {stage5_49[6], stage5_49[7]},
      {stage5_50[0], stage5_50[1]},
      {stage6_51[1],stage6_50[1],stage6_49[2],stage6_48[3]}
   );
   gpc606_5 gpc5764 (
      {stage5_50[2], stage5_50[3], stage5_50[4], stage5_50[5], stage5_50[6], stage5_50[7]},
      {stage5_52[0], stage5_52[1], stage5_52[2], stage5_52[3], stage5_52[4], stage5_52[5]},
      {stage6_54[0],stage6_53[0],stage6_52[0],stage6_51[2],stage6_50[2]}
   );
   gpc615_5 gpc5765 (
      {stage5_51[0], stage5_51[1], stage5_51[2], stage5_51[3], stage5_51[4]},
      {stage5_52[6]},
      {stage5_53[0], stage5_53[1], stage5_53[2], stage5_53[3], stage5_53[4], stage5_53[5]},
      {stage6_55[0],stage6_54[1],stage6_53[1],stage6_52[1],stage6_51[3]}
   );
   gpc615_5 gpc5766 (
      {stage5_51[5], stage5_51[6], stage5_51[7], stage5_51[8], stage5_51[9]},
      {stage5_52[7]},
      {stage5_53[6], stage5_53[7], stage5_53[8], stage5_53[9], stage5_53[10], stage5_53[11]},
      {stage6_55[1],stage6_54[2],stage6_53[2],stage6_52[2],stage6_51[4]}
   );
   gpc1163_5 gpc5767 (
      {stage5_53[12], stage5_53[13], stage5_53[14]},
      {stage5_54[0], stage5_54[1], stage5_54[2], stage5_54[3], stage5_54[4], stage5_54[5]},
      {stage5_55[0]},
      {stage5_56[0]},
      {stage6_57[0],stage6_56[0],stage6_55[2],stage6_54[3],stage6_53[3]}
   );
   gpc615_5 gpc5768 (
      {stage5_55[1], stage5_55[2], stage5_55[3], stage5_55[4], stage5_55[5]},
      {stage5_56[1]},
      {stage5_57[0], stage5_57[1], stage5_57[2], stage5_57[3], stage5_57[4], stage5_57[5]},
      {stage6_59[0],stage6_58[0],stage6_57[1],stage6_56[1],stage6_55[3]}
   );
   gpc615_5 gpc5769 (
      {stage5_58[0], stage5_58[1], stage5_58[2], stage5_58[3], stage5_58[4]},
      {stage5_59[0]},
      {stage5_60[0], stage5_60[1], stage5_60[2], stage5_60[3], stage5_60[4], stage5_60[5]},
      {stage6_62[0],stage6_61[0],stage6_60[0],stage6_59[1],stage6_58[1]}
   );
   gpc3_2 gpc5770 (
      {stage5_59[1], stage5_59[2], stage5_59[3]},
      {stage6_60[1],stage6_59[2]}
   );
   gpc606_5 gpc5771 (
      {stage5_63[0], stage5_63[1], stage5_63[2], stage5_63[3], stage5_63[4], stage5_63[5]},
      {stage5_65[0], stage5_65[1], stage5_65[2], stage5_65[3], stage5_65[4], 1'b0},
      {stage6_67[0],stage6_66[0],stage6_65[0],stage6_64[0],stage6_63[0]}
   );
   gpc606_5 gpc5772 (
      {stage5_64[0], stage5_64[1], stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5]},
      {stage5_66[0], stage5_66[1], stage5_66[2], stage5_66[3], stage5_66[4], stage5_66[5]},
      {stage6_68[0],stage6_67[1],stage6_66[1],stage6_65[1],stage6_64[1]}
   );
   gpc606_5 gpc5773 (
      {stage5_66[6], stage5_66[7], stage5_66[8], stage5_66[9], stage5_66[10], 1'b0},
      {stage5_68[0], stage5_68[1], stage5_68[2], stage5_68[3], stage5_68[4], 1'b0},
      {stage6_70[0],stage6_69[0],stage6_68[1],stage6_67[2],stage6_66[2]}
   );
   gpc606_5 gpc5774 (
      {stage5_67[0], stage5_67[1], stage5_67[2], stage5_67[3], stage5_67[4], stage5_67[5]},
      {stage5_69[0], stage5_69[1], stage5_69[2], 1'b0, 1'b0, 1'b0},
      {stage6_71[0],stage6_70[1],stage6_69[1],stage6_68[2],stage6_67[3]}
   );
   gpc1_1 gpc5775 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc5776 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc5777 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc5778 (
      {stage5_0[3]},
      {stage6_0[3]}
   );
   gpc1_1 gpc5779 (
      {stage5_0[4]},
      {stage6_0[4]}
   );
   gpc1_1 gpc5780 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc5781 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc5782 (
      {stage5_1[2]},
      {stage6_1[2]}
   );
   gpc1_1 gpc5783 (
      {stage5_1[3]},
      {stage6_1[3]}
   );
   gpc1_1 gpc5784 (
      {stage5_4[8]},
      {stage6_4[3]}
   );
   gpc1_1 gpc5785 (
      {stage5_4[9]},
      {stage6_4[4]}
   );
   gpc1_1 gpc5786 (
      {stage5_5[7]},
      {stage6_5[3]}
   );
   gpc1_1 gpc5787 (
      {stage5_9[3]},
      {stage6_9[2]}
   );
   gpc1_1 gpc5788 (
      {stage5_9[4]},
      {stage6_9[3]}
   );
   gpc1_1 gpc5789 (
      {stage5_9[5]},
      {stage6_9[4]}
   );
   gpc1_1 gpc5790 (
      {stage5_9[6]},
      {stage6_9[5]}
   );
   gpc1_1 gpc5791 (
      {stage5_9[7]},
      {stage6_9[6]}
   );
   gpc1_1 gpc5792 (
      {stage5_9[8]},
      {stage6_9[7]}
   );
   gpc1_1 gpc5793 (
      {stage5_9[9]},
      {stage6_9[8]}
   );
   gpc1_1 gpc5794 (
      {stage5_11[6]},
      {stage6_11[2]}
   );
   gpc1_1 gpc5795 (
      {stage5_11[7]},
      {stage6_11[3]}
   );
   gpc1_1 gpc5796 (
      {stage5_11[8]},
      {stage6_11[4]}
   );
   gpc1_1 gpc5797 (
      {stage5_11[9]},
      {stage6_11[5]}
   );
   gpc1_1 gpc5798 (
      {stage5_14[0]},
      {stage6_14[2]}
   );
   gpc1_1 gpc5799 (
      {stage5_14[1]},
      {stage6_14[3]}
   );
   gpc1_1 gpc5800 (
      {stage5_14[2]},
      {stage6_14[4]}
   );
   gpc1_1 gpc5801 (
      {stage5_14[3]},
      {stage6_14[5]}
   );
   gpc1_1 gpc5802 (
      {stage5_14[4]},
      {stage6_14[6]}
   );
   gpc1_1 gpc5803 (
      {stage5_15[5]},
      {stage6_15[2]}
   );
   gpc1_1 gpc5804 (
      {stage5_17[7]},
      {stage6_17[2]}
   );
   gpc1_1 gpc5805 (
      {stage5_18[4]},
      {stage6_18[2]}
   );
   gpc1_1 gpc5806 (
      {stage5_18[5]},
      {stage6_18[3]}
   );
   gpc1_1 gpc5807 (
      {stage5_20[2]},
      {stage6_20[3]}
   );
   gpc1_1 gpc5808 (
      {stage5_23[1]},
      {stage6_23[3]}
   );
   gpc1_1 gpc5809 (
      {stage5_23[2]},
      {stage6_23[4]}
   );
   gpc1_1 gpc5810 (
      {stage5_24[6]},
      {stage6_24[1]}
   );
   gpc1_1 gpc5811 (
      {stage5_25[0]},
      {stage6_25[1]}
   );
   gpc1_1 gpc5812 (
      {stage5_25[1]},
      {stage6_25[2]}
   );
   gpc1_1 gpc5813 (
      {stage5_25[2]},
      {stage6_25[3]}
   );
   gpc1_1 gpc5814 (
      {stage5_25[3]},
      {stage6_25[4]}
   );
   gpc1_1 gpc5815 (
      {stage5_25[4]},
      {stage6_25[5]}
   );
   gpc1_1 gpc5816 (
      {stage5_25[5]},
      {stage6_25[6]}
   );
   gpc1_1 gpc5817 (
      {stage5_27[5]},
      {stage6_27[2]}
   );
   gpc1_1 gpc5818 (
      {stage5_35[4]},
      {stage6_35[3]}
   );
   gpc1_1 gpc5819 (
      {stage5_37[6]},
      {stage6_37[2]}
   );
   gpc1_1 gpc5820 (
      {stage5_37[7]},
      {stage6_37[3]}
   );
   gpc1_1 gpc5821 (
      {stage5_37[8]},
      {stage6_37[4]}
   );
   gpc1_1 gpc5822 (
      {stage5_37[9]},
      {stage6_37[5]}
   );
   gpc1_1 gpc5823 (
      {stage5_37[10]},
      {stage6_37[6]}
   );
   gpc1_1 gpc5824 (
      {stage5_37[11]},
      {stage6_37[7]}
   );
   gpc1_1 gpc5825 (
      {stage5_43[7]},
      {stage6_43[3]}
   );
   gpc1_1 gpc5826 (
      {stage5_43[8]},
      {stage6_43[4]}
   );
   gpc1_1 gpc5827 (
      {stage5_43[9]},
      {stage6_43[5]}
   );
   gpc1_1 gpc5828 (
      {stage5_47[4]},
      {stage6_47[3]}
   );
   gpc1_1 gpc5829 (
      {stage5_47[5]},
      {stage6_47[4]}
   );
   gpc1_1 gpc5830 (
      {stage5_47[6]},
      {stage6_47[5]}
   );
   gpc1_1 gpc5831 (
      {stage5_50[8]},
      {stage6_50[3]}
   );
   gpc1_1 gpc5832 (
      {stage5_56[2]},
      {stage6_56[2]}
   );
   gpc1_1 gpc5833 (
      {stage5_56[3]},
      {stage6_56[3]}
   );
   gpc1_1 gpc5834 (
      {stage5_56[4]},
      {stage6_56[4]}
   );
   gpc1_1 gpc5835 (
      {stage5_56[5]},
      {stage6_56[5]}
   );
   gpc1_1 gpc5836 (
      {stage5_57[6]},
      {stage6_57[2]}
   );
   gpc1_1 gpc5837 (
      {stage5_59[4]},
      {stage6_59[3]}
   );
   gpc1_1 gpc5838 (
      {stage5_59[5]},
      {stage6_59[4]}
   );
   gpc1_1 gpc5839 (
      {stage5_59[6]},
      {stage6_59[5]}
   );
   gpc1_1 gpc5840 (
      {stage5_60[6]},
      {stage6_60[2]}
   );
   gpc1_1 gpc5841 (
      {stage5_60[7]},
      {stage6_60[3]}
   );
   gpc1_1 gpc5842 (
      {stage5_60[8]},
      {stage6_60[4]}
   );
   gpc1_1 gpc5843 (
      {stage5_61[0]},
      {stage6_61[1]}
   );
   gpc1_1 gpc5844 (
      {stage5_61[1]},
      {stage6_61[2]}
   );
   gpc1_1 gpc5845 (
      {stage5_61[2]},
      {stage6_61[3]}
   );
   gpc1_1 gpc5846 (
      {stage5_61[3]},
      {stage6_61[4]}
   );
   gpc1_1 gpc5847 (
      {stage5_62[0]},
      {stage6_62[1]}
   );
   gpc1_1 gpc5848 (
      {stage5_62[1]},
      {stage6_62[2]}
   );
   gpc1_1 gpc5849 (
      {stage5_62[2]},
      {stage6_62[3]}
   );
   gpc1_1 gpc5850 (
      {stage5_62[3]},
      {stage6_62[4]}
   );
   gpc1_1 gpc5851 (
      {stage5_67[6]},
      {stage6_67[4]}
   );
   gpc135_4 gpc5852 (
      {stage6_0[0], stage6_0[1], stage6_0[2], stage6_0[3], stage6_0[4]},
      {stage6_1[0], stage6_1[1], stage6_1[2]},
      {stage6_2[0]},
      {stage7_3[0],stage7_2[0],stage7_1[0],stage7_0[0]}
   );
   gpc1343_5 gpc5853 (
      {stage6_3[0], stage6_3[1], 1'b0},
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3]},
      {stage6_5[0], stage6_5[1], stage6_5[2]},
      {stage6_6[0]},
      {stage7_7[0],stage7_6[0],stage7_5[0],stage7_4[0],stage7_3[1]}
   );
   gpc1423_5 gpc5854 (
      {stage6_7[0], stage6_7[1], stage6_7[2]},
      {stage6_8[0], stage6_8[1]},
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3]},
      {stage6_10[0]},
      {stage7_11[0],stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[1]}
   );
   gpc615_5 gpc5855 (
      {stage6_9[4], stage6_9[5], stage6_9[6], stage6_9[7], stage6_9[8]},
      {stage6_10[1]},
      {stage6_11[0], stage6_11[1], stage6_11[2], stage6_11[3], stage6_11[4], stage6_11[5]},
      {stage7_13[0],stage7_12[0],stage7_11[1],stage7_10[1],stage7_9[1]}
   );
   gpc623_5 gpc5856 (
      {stage6_12[0], stage6_12[1], stage6_12[2]},
      {stage6_13[0], stage6_13[1]},
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], stage6_14[5]},
      {stage7_16[0],stage7_15[0],stage7_14[0],stage7_13[1],stage7_12[1]}
   );
   gpc2223_5 gpc5857 (
      {stage6_15[0], stage6_15[1], stage6_15[2]},
      {stage6_16[0], stage6_16[1]},
      {stage6_17[0], stage6_17[1]},
      {stage6_18[0], stage6_18[1]},
      {stage7_19[0],stage7_18[0],stage7_17[0],stage7_16[1],stage7_15[1]}
   );
   gpc1343_5 gpc5858 (
      {stage6_18[2], stage6_18[3], 1'b0},
      {stage6_19[0], stage6_19[1], stage6_19[2], stage6_19[3]},
      {stage6_20[0], stage6_20[1], stage6_20[2]},
      {stage6_21[0]},
      {stage7_22[0],stage7_21[0],stage7_20[0],stage7_19[1],stage7_18[1]}
   );
   gpc3_2 gpc5859 (
      {stage6_22[0], stage6_22[1], stage6_22[2]},
      {stage7_23[0],stage7_22[1]}
   );
   gpc1415_5 gpc5860 (
      {stage6_23[0], stage6_23[1], stage6_23[2], stage6_23[3], stage6_23[4]},
      {stage6_24[0]},
      {stage6_25[0], stage6_25[1], stage6_25[2], stage6_25[3]},
      {stage6_26[0]},
      {stage7_27[0],stage7_26[0],stage7_25[0],stage7_24[0],stage7_23[1]}
   );
   gpc1343_5 gpc5861 (
      {stage6_25[4], stage6_25[5], stage6_25[6]},
      {stage6_26[1], 1'b0, 1'b0, 1'b0},
      {stage6_27[0], stage6_27[1], stage6_27[2]},
      {stage6_28[0]},
      {stage7_29[0],stage7_28[0],stage7_27[1],stage7_26[1],stage7_25[1]}
   );
   gpc1423_5 gpc5862 (
      {stage6_29[0], stage6_29[1], stage6_29[2]},
      {stage6_30[0], stage6_30[1]},
      {stage6_31[0], stage6_31[1], stage6_31[2], 1'b0},
      {stage6_32[0]},
      {stage7_33[0],stage7_32[0],stage7_31[0],stage7_30[0],stage7_29[1]}
   );
   gpc1343_5 gpc5863 (
      {stage6_32[1], stage6_32[2], 1'b0},
      {stage6_33[0], stage6_33[1], stage6_33[2], stage6_33[3]},
      {stage6_34[0], stage6_34[1], stage6_34[2]},
      {stage6_35[0]},
      {stage7_36[0],stage7_35[0],stage7_34[0],stage7_33[1],stage7_32[1]}
   );
   gpc1343_5 gpc5864 (
      {stage6_35[1], stage6_35[2], stage6_35[3]},
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3]},
      {stage6_37[0], stage6_37[1], stage6_37[2]},
      {stage6_38[0]},
      {stage7_39[0],stage7_38[0],stage7_37[0],stage7_36[1],stage7_35[1]}
   );
   gpc1325_5 gpc5865 (
      {stage6_37[3], stage6_37[4], stage6_37[5], stage6_37[6], stage6_37[7]},
      {stage6_38[1], 1'b0},
      {stage6_39[0], stage6_39[1], stage6_39[2]},
      {stage6_40[0]},
      {stage7_41[0],stage7_40[0],stage7_39[1],stage7_38[1],stage7_37[1]}
   );
   gpc223_4 gpc5866 (
      {stage6_41[0], stage6_41[1], 1'b0},
      {stage6_42[0], stage6_42[1]},
      {stage6_43[0], stage6_43[1]},
      {stage7_44[0],stage7_43[0],stage7_42[0],stage7_41[1]}
   );
   gpc1343_5 gpc5867 (
      {stage6_42[2], 1'b0, 1'b0},
      {stage6_43[2], stage6_43[3], stage6_43[4], stage6_43[5]},
      {stage6_44[0], stage6_44[1], stage6_44[2]},
      {stage6_45[0]},
      {stage7_46[0],stage7_45[0],stage7_44[1],stage7_43[1],stage7_42[1]}
   );
   gpc623_5 gpc5868 (
      {stage6_45[1], stage6_45[2], stage6_45[3]},
      {stage6_46[0], stage6_46[1]},
      {stage6_47[0], stage6_47[1], stage6_47[2], stage6_47[3], stage6_47[4], stage6_47[5]},
      {stage7_49[0],stage7_48[0],stage7_47[0],stage7_46[1],stage7_45[1]}
   );
   gpc2135_5 gpc5869 (
      {stage6_48[0], stage6_48[1], stage6_48[2], stage6_48[3], 1'b0},
      {stage6_49[0], stage6_49[1], stage6_49[2]},
      {stage6_50[0]},
      {stage6_51[0], stage6_51[1]},
      {stage7_52[0],stage7_51[0],stage7_50[0],stage7_49[1],stage7_48[1]}
   );
   gpc1343_5 gpc5870 (
      {stage6_50[1], stage6_50[2], stage6_50[3]},
      {stage6_51[2], stage6_51[3], stage6_51[4], 1'b0},
      {stage6_52[0], stage6_52[1], stage6_52[2]},
      {stage6_53[0]},
      {stage7_54[0],stage7_53[0],stage7_52[1],stage7_51[1],stage7_50[1]}
   );
   gpc1343_5 gpc5871 (
      {stage6_53[1], stage6_53[2], stage6_53[3]},
      {stage6_54[0], stage6_54[1], stage6_54[2], stage6_54[3]},
      {stage6_55[0], stage6_55[1], stage6_55[2]},
      {stage6_56[0]},
      {stage7_57[0],stage7_56[0],stage7_55[0],stage7_54[1],stage7_53[1]}
   );
   gpc135_4 gpc5872 (
      {stage6_56[1], stage6_56[2], stage6_56[3], stage6_56[4], stage6_56[5]},
      {stage6_57[0], stage6_57[1], stage6_57[2]},
      {stage6_58[0]},
      {stage7_59[0],stage7_58[0],stage7_57[1],stage7_56[1]}
   );
   gpc1406_5 gpc5873 (
      {stage6_59[0], stage6_59[1], stage6_59[2], stage6_59[3], stage6_59[4], stage6_59[5]},
      {stage6_61[0], stage6_61[1], stage6_61[2], stage6_61[3]},
      {stage6_62[0]},
      {stage7_63[0],stage7_62[0],stage7_61[0],stage7_60[0],stage7_59[1]}
   );
   gpc1415_5 gpc5874 (
      {stage6_60[0], stage6_60[1], stage6_60[2], stage6_60[3], stage6_60[4]},
      {stage6_61[4]},
      {stage6_62[1], stage6_62[2], stage6_62[3], stage6_62[4]},
      {stage6_63[0]},
      {stage7_64[0],stage7_63[1],stage7_62[1],stage7_61[1],stage7_60[1]}
   );
   gpc23_3 gpc5875 (
      {stage6_64[0], stage6_64[1], 1'b0},
      {stage6_65[0], stage6_65[1]},
      {stage7_66[0],stage7_65[0],stage7_64[1]}
   );
   gpc1343_5 gpc5876 (
      {stage6_66[0], stage6_66[1], stage6_66[2]},
      {stage6_67[0], stage6_67[1], stage6_67[2], stage6_67[3]},
      {stage6_68[0], stage6_68[1], stage6_68[2]},
      {stage6_69[0]},
      {stage7_70[0],stage7_69[0],stage7_68[0],stage7_67[0],stage7_66[1]}
   );
   gpc2223_5 gpc5877 (
      {1'b0, 1'b0, 1'b0},
      {stage6_69[1], 1'b0},
      {stage6_70[0], stage6_70[1]},
      {stage6_71[0], 1'b0},
      {stage7_71[0],stage7_70[1],stage7_69[1],stage7_68[1]}
   );
   gpc1_1 gpc5878 (
      {stage6_1[3]},
      {stage7_1[1]}
   );
   gpc1_1 gpc5879 (
      {stage6_4[4]},
      {stage7_4[1]}
   );
   gpc1_1 gpc5880 (
      {stage6_5[3]},
      {stage7_5[1]}
   );
   gpc1_1 gpc5881 (
      {stage6_6[1]},
      {stage7_6[1]}
   );
   gpc1_1 gpc5882 (
      {stage6_8[2]},
      {stage7_8[1]}
   );
   gpc1_1 gpc5883 (
      {stage6_14[6]},
      {stage7_14[1]}
   );
   gpc1_1 gpc5884 (
      {stage6_17[2]},
      {stage7_17[1]}
   );
   gpc1_1 gpc5885 (
      {stage6_20[3]},
      {stage7_20[1]}
   );
   gpc1_1 gpc5886 (
      {stage6_21[1]},
      {stage7_21[1]}
   );
   gpc1_1 gpc5887 (
      {stage6_24[1]},
      {stage7_24[1]}
   );
   gpc1_1 gpc5888 (
      {stage6_28[1]},
      {stage7_28[1]}
   );
   gpc1_1 gpc5889 (
      {stage6_30[2]},
      {stage7_30[1]}
   );
   gpc1_1 gpc5890 (
      {stage6_40[1]},
      {stage7_40[1]}
   );
   gpc1_1 gpc5891 (
      {stage6_55[3]},
      {stage7_55[1]}
   );
   gpc1_1 gpc5892 (
      {stage6_58[1]},
      {stage7_58[1]}
   );
   gpc1_1 gpc5893 (
      {stage6_67[4]},
      {stage7_67[1]}
   );
endmodule

module testbench();
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    reg [255:0] src16;
    reg [255:0] src17;
    reg [255:0] src18;
    reg [255:0] src19;
    reg [255:0] src20;
    reg [255:0] src21;
    reg [255:0] src22;
    reg [255:0] src23;
    reg [255:0] src24;
    reg [255:0] src25;
    reg [255:0] src26;
    reg [255:0] src27;
    reg [255:0] src28;
    reg [255:0] src29;
    reg [255:0] src30;
    reg [255:0] src31;
    reg [255:0] src32;
    reg [255:0] src33;
    reg [255:0] src34;
    reg [255:0] src35;
    reg [255:0] src36;
    reg [255:0] src37;
    reg [255:0] src38;
    reg [255:0] src39;
    reg [255:0] src40;
    reg [255:0] src41;
    reg [255:0] src42;
    reg [255:0] src43;
    reg [255:0] src44;
    reg [255:0] src45;
    reg [255:0] src46;
    reg [255:0] src47;
    reg [255:0] src48;
    reg [255:0] src49;
    reg [255:0] src50;
    reg [255:0] src51;
    reg [255:0] src52;
    reg [255:0] src53;
    reg [255:0] src54;
    reg [255:0] src55;
    reg [255:0] src56;
    reg [255:0] src57;
    reg [255:0] src58;
    reg [255:0] src59;
    reg [255:0] src60;
    reg [255:0] src61;
    reg [255:0] src62;
    reg [255:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [0:0] dst71;
    wire [71:0] srcsum;
    wire [71:0] dstsum;
    wire test;
    compressor_CLA256_64 compressor_CLA256_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70),
        .dst71(dst71));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127] + src32[128] + src32[129] + src32[130] + src32[131] + src32[132] + src32[133] + src32[134] + src32[135] + src32[136] + src32[137] + src32[138] + src32[139] + src32[140] + src32[141] + src32[142] + src32[143] + src32[144] + src32[145] + src32[146] + src32[147] + src32[148] + src32[149] + src32[150] + src32[151] + src32[152] + src32[153] + src32[154] + src32[155] + src32[156] + src32[157] + src32[158] + src32[159] + src32[160] + src32[161] + src32[162] + src32[163] + src32[164] + src32[165] + src32[166] + src32[167] + src32[168] + src32[169] + src32[170] + src32[171] + src32[172] + src32[173] + src32[174] + src32[175] + src32[176] + src32[177] + src32[178] + src32[179] + src32[180] + src32[181] + src32[182] + src32[183] + src32[184] + src32[185] + src32[186] + src32[187] + src32[188] + src32[189] + src32[190] + src32[191] + src32[192] + src32[193] + src32[194] + src32[195] + src32[196] + src32[197] + src32[198] + src32[199] + src32[200] + src32[201] + src32[202] + src32[203] + src32[204] + src32[205] + src32[206] + src32[207] + src32[208] + src32[209] + src32[210] + src32[211] + src32[212] + src32[213] + src32[214] + src32[215] + src32[216] + src32[217] + src32[218] + src32[219] + src32[220] + src32[221] + src32[222] + src32[223] + src32[224] + src32[225] + src32[226] + src32[227] + src32[228] + src32[229] + src32[230] + src32[231] + src32[232] + src32[233] + src32[234] + src32[235] + src32[236] + src32[237] + src32[238] + src32[239] + src32[240] + src32[241] + src32[242] + src32[243] + src32[244] + src32[245] + src32[246] + src32[247] + src32[248] + src32[249] + src32[250] + src32[251] + src32[252] + src32[253] + src32[254] + src32[255])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127] + src33[128] + src33[129] + src33[130] + src33[131] + src33[132] + src33[133] + src33[134] + src33[135] + src33[136] + src33[137] + src33[138] + src33[139] + src33[140] + src33[141] + src33[142] + src33[143] + src33[144] + src33[145] + src33[146] + src33[147] + src33[148] + src33[149] + src33[150] + src33[151] + src33[152] + src33[153] + src33[154] + src33[155] + src33[156] + src33[157] + src33[158] + src33[159] + src33[160] + src33[161] + src33[162] + src33[163] + src33[164] + src33[165] + src33[166] + src33[167] + src33[168] + src33[169] + src33[170] + src33[171] + src33[172] + src33[173] + src33[174] + src33[175] + src33[176] + src33[177] + src33[178] + src33[179] + src33[180] + src33[181] + src33[182] + src33[183] + src33[184] + src33[185] + src33[186] + src33[187] + src33[188] + src33[189] + src33[190] + src33[191] + src33[192] + src33[193] + src33[194] + src33[195] + src33[196] + src33[197] + src33[198] + src33[199] + src33[200] + src33[201] + src33[202] + src33[203] + src33[204] + src33[205] + src33[206] + src33[207] + src33[208] + src33[209] + src33[210] + src33[211] + src33[212] + src33[213] + src33[214] + src33[215] + src33[216] + src33[217] + src33[218] + src33[219] + src33[220] + src33[221] + src33[222] + src33[223] + src33[224] + src33[225] + src33[226] + src33[227] + src33[228] + src33[229] + src33[230] + src33[231] + src33[232] + src33[233] + src33[234] + src33[235] + src33[236] + src33[237] + src33[238] + src33[239] + src33[240] + src33[241] + src33[242] + src33[243] + src33[244] + src33[245] + src33[246] + src33[247] + src33[248] + src33[249] + src33[250] + src33[251] + src33[252] + src33[253] + src33[254] + src33[255])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127] + src34[128] + src34[129] + src34[130] + src34[131] + src34[132] + src34[133] + src34[134] + src34[135] + src34[136] + src34[137] + src34[138] + src34[139] + src34[140] + src34[141] + src34[142] + src34[143] + src34[144] + src34[145] + src34[146] + src34[147] + src34[148] + src34[149] + src34[150] + src34[151] + src34[152] + src34[153] + src34[154] + src34[155] + src34[156] + src34[157] + src34[158] + src34[159] + src34[160] + src34[161] + src34[162] + src34[163] + src34[164] + src34[165] + src34[166] + src34[167] + src34[168] + src34[169] + src34[170] + src34[171] + src34[172] + src34[173] + src34[174] + src34[175] + src34[176] + src34[177] + src34[178] + src34[179] + src34[180] + src34[181] + src34[182] + src34[183] + src34[184] + src34[185] + src34[186] + src34[187] + src34[188] + src34[189] + src34[190] + src34[191] + src34[192] + src34[193] + src34[194] + src34[195] + src34[196] + src34[197] + src34[198] + src34[199] + src34[200] + src34[201] + src34[202] + src34[203] + src34[204] + src34[205] + src34[206] + src34[207] + src34[208] + src34[209] + src34[210] + src34[211] + src34[212] + src34[213] + src34[214] + src34[215] + src34[216] + src34[217] + src34[218] + src34[219] + src34[220] + src34[221] + src34[222] + src34[223] + src34[224] + src34[225] + src34[226] + src34[227] + src34[228] + src34[229] + src34[230] + src34[231] + src34[232] + src34[233] + src34[234] + src34[235] + src34[236] + src34[237] + src34[238] + src34[239] + src34[240] + src34[241] + src34[242] + src34[243] + src34[244] + src34[245] + src34[246] + src34[247] + src34[248] + src34[249] + src34[250] + src34[251] + src34[252] + src34[253] + src34[254] + src34[255])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127] + src35[128] + src35[129] + src35[130] + src35[131] + src35[132] + src35[133] + src35[134] + src35[135] + src35[136] + src35[137] + src35[138] + src35[139] + src35[140] + src35[141] + src35[142] + src35[143] + src35[144] + src35[145] + src35[146] + src35[147] + src35[148] + src35[149] + src35[150] + src35[151] + src35[152] + src35[153] + src35[154] + src35[155] + src35[156] + src35[157] + src35[158] + src35[159] + src35[160] + src35[161] + src35[162] + src35[163] + src35[164] + src35[165] + src35[166] + src35[167] + src35[168] + src35[169] + src35[170] + src35[171] + src35[172] + src35[173] + src35[174] + src35[175] + src35[176] + src35[177] + src35[178] + src35[179] + src35[180] + src35[181] + src35[182] + src35[183] + src35[184] + src35[185] + src35[186] + src35[187] + src35[188] + src35[189] + src35[190] + src35[191] + src35[192] + src35[193] + src35[194] + src35[195] + src35[196] + src35[197] + src35[198] + src35[199] + src35[200] + src35[201] + src35[202] + src35[203] + src35[204] + src35[205] + src35[206] + src35[207] + src35[208] + src35[209] + src35[210] + src35[211] + src35[212] + src35[213] + src35[214] + src35[215] + src35[216] + src35[217] + src35[218] + src35[219] + src35[220] + src35[221] + src35[222] + src35[223] + src35[224] + src35[225] + src35[226] + src35[227] + src35[228] + src35[229] + src35[230] + src35[231] + src35[232] + src35[233] + src35[234] + src35[235] + src35[236] + src35[237] + src35[238] + src35[239] + src35[240] + src35[241] + src35[242] + src35[243] + src35[244] + src35[245] + src35[246] + src35[247] + src35[248] + src35[249] + src35[250] + src35[251] + src35[252] + src35[253] + src35[254] + src35[255])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127] + src36[128] + src36[129] + src36[130] + src36[131] + src36[132] + src36[133] + src36[134] + src36[135] + src36[136] + src36[137] + src36[138] + src36[139] + src36[140] + src36[141] + src36[142] + src36[143] + src36[144] + src36[145] + src36[146] + src36[147] + src36[148] + src36[149] + src36[150] + src36[151] + src36[152] + src36[153] + src36[154] + src36[155] + src36[156] + src36[157] + src36[158] + src36[159] + src36[160] + src36[161] + src36[162] + src36[163] + src36[164] + src36[165] + src36[166] + src36[167] + src36[168] + src36[169] + src36[170] + src36[171] + src36[172] + src36[173] + src36[174] + src36[175] + src36[176] + src36[177] + src36[178] + src36[179] + src36[180] + src36[181] + src36[182] + src36[183] + src36[184] + src36[185] + src36[186] + src36[187] + src36[188] + src36[189] + src36[190] + src36[191] + src36[192] + src36[193] + src36[194] + src36[195] + src36[196] + src36[197] + src36[198] + src36[199] + src36[200] + src36[201] + src36[202] + src36[203] + src36[204] + src36[205] + src36[206] + src36[207] + src36[208] + src36[209] + src36[210] + src36[211] + src36[212] + src36[213] + src36[214] + src36[215] + src36[216] + src36[217] + src36[218] + src36[219] + src36[220] + src36[221] + src36[222] + src36[223] + src36[224] + src36[225] + src36[226] + src36[227] + src36[228] + src36[229] + src36[230] + src36[231] + src36[232] + src36[233] + src36[234] + src36[235] + src36[236] + src36[237] + src36[238] + src36[239] + src36[240] + src36[241] + src36[242] + src36[243] + src36[244] + src36[245] + src36[246] + src36[247] + src36[248] + src36[249] + src36[250] + src36[251] + src36[252] + src36[253] + src36[254] + src36[255])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127] + src37[128] + src37[129] + src37[130] + src37[131] + src37[132] + src37[133] + src37[134] + src37[135] + src37[136] + src37[137] + src37[138] + src37[139] + src37[140] + src37[141] + src37[142] + src37[143] + src37[144] + src37[145] + src37[146] + src37[147] + src37[148] + src37[149] + src37[150] + src37[151] + src37[152] + src37[153] + src37[154] + src37[155] + src37[156] + src37[157] + src37[158] + src37[159] + src37[160] + src37[161] + src37[162] + src37[163] + src37[164] + src37[165] + src37[166] + src37[167] + src37[168] + src37[169] + src37[170] + src37[171] + src37[172] + src37[173] + src37[174] + src37[175] + src37[176] + src37[177] + src37[178] + src37[179] + src37[180] + src37[181] + src37[182] + src37[183] + src37[184] + src37[185] + src37[186] + src37[187] + src37[188] + src37[189] + src37[190] + src37[191] + src37[192] + src37[193] + src37[194] + src37[195] + src37[196] + src37[197] + src37[198] + src37[199] + src37[200] + src37[201] + src37[202] + src37[203] + src37[204] + src37[205] + src37[206] + src37[207] + src37[208] + src37[209] + src37[210] + src37[211] + src37[212] + src37[213] + src37[214] + src37[215] + src37[216] + src37[217] + src37[218] + src37[219] + src37[220] + src37[221] + src37[222] + src37[223] + src37[224] + src37[225] + src37[226] + src37[227] + src37[228] + src37[229] + src37[230] + src37[231] + src37[232] + src37[233] + src37[234] + src37[235] + src37[236] + src37[237] + src37[238] + src37[239] + src37[240] + src37[241] + src37[242] + src37[243] + src37[244] + src37[245] + src37[246] + src37[247] + src37[248] + src37[249] + src37[250] + src37[251] + src37[252] + src37[253] + src37[254] + src37[255])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127] + src38[128] + src38[129] + src38[130] + src38[131] + src38[132] + src38[133] + src38[134] + src38[135] + src38[136] + src38[137] + src38[138] + src38[139] + src38[140] + src38[141] + src38[142] + src38[143] + src38[144] + src38[145] + src38[146] + src38[147] + src38[148] + src38[149] + src38[150] + src38[151] + src38[152] + src38[153] + src38[154] + src38[155] + src38[156] + src38[157] + src38[158] + src38[159] + src38[160] + src38[161] + src38[162] + src38[163] + src38[164] + src38[165] + src38[166] + src38[167] + src38[168] + src38[169] + src38[170] + src38[171] + src38[172] + src38[173] + src38[174] + src38[175] + src38[176] + src38[177] + src38[178] + src38[179] + src38[180] + src38[181] + src38[182] + src38[183] + src38[184] + src38[185] + src38[186] + src38[187] + src38[188] + src38[189] + src38[190] + src38[191] + src38[192] + src38[193] + src38[194] + src38[195] + src38[196] + src38[197] + src38[198] + src38[199] + src38[200] + src38[201] + src38[202] + src38[203] + src38[204] + src38[205] + src38[206] + src38[207] + src38[208] + src38[209] + src38[210] + src38[211] + src38[212] + src38[213] + src38[214] + src38[215] + src38[216] + src38[217] + src38[218] + src38[219] + src38[220] + src38[221] + src38[222] + src38[223] + src38[224] + src38[225] + src38[226] + src38[227] + src38[228] + src38[229] + src38[230] + src38[231] + src38[232] + src38[233] + src38[234] + src38[235] + src38[236] + src38[237] + src38[238] + src38[239] + src38[240] + src38[241] + src38[242] + src38[243] + src38[244] + src38[245] + src38[246] + src38[247] + src38[248] + src38[249] + src38[250] + src38[251] + src38[252] + src38[253] + src38[254] + src38[255])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127] + src39[128] + src39[129] + src39[130] + src39[131] + src39[132] + src39[133] + src39[134] + src39[135] + src39[136] + src39[137] + src39[138] + src39[139] + src39[140] + src39[141] + src39[142] + src39[143] + src39[144] + src39[145] + src39[146] + src39[147] + src39[148] + src39[149] + src39[150] + src39[151] + src39[152] + src39[153] + src39[154] + src39[155] + src39[156] + src39[157] + src39[158] + src39[159] + src39[160] + src39[161] + src39[162] + src39[163] + src39[164] + src39[165] + src39[166] + src39[167] + src39[168] + src39[169] + src39[170] + src39[171] + src39[172] + src39[173] + src39[174] + src39[175] + src39[176] + src39[177] + src39[178] + src39[179] + src39[180] + src39[181] + src39[182] + src39[183] + src39[184] + src39[185] + src39[186] + src39[187] + src39[188] + src39[189] + src39[190] + src39[191] + src39[192] + src39[193] + src39[194] + src39[195] + src39[196] + src39[197] + src39[198] + src39[199] + src39[200] + src39[201] + src39[202] + src39[203] + src39[204] + src39[205] + src39[206] + src39[207] + src39[208] + src39[209] + src39[210] + src39[211] + src39[212] + src39[213] + src39[214] + src39[215] + src39[216] + src39[217] + src39[218] + src39[219] + src39[220] + src39[221] + src39[222] + src39[223] + src39[224] + src39[225] + src39[226] + src39[227] + src39[228] + src39[229] + src39[230] + src39[231] + src39[232] + src39[233] + src39[234] + src39[235] + src39[236] + src39[237] + src39[238] + src39[239] + src39[240] + src39[241] + src39[242] + src39[243] + src39[244] + src39[245] + src39[246] + src39[247] + src39[248] + src39[249] + src39[250] + src39[251] + src39[252] + src39[253] + src39[254] + src39[255])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127] + src40[128] + src40[129] + src40[130] + src40[131] + src40[132] + src40[133] + src40[134] + src40[135] + src40[136] + src40[137] + src40[138] + src40[139] + src40[140] + src40[141] + src40[142] + src40[143] + src40[144] + src40[145] + src40[146] + src40[147] + src40[148] + src40[149] + src40[150] + src40[151] + src40[152] + src40[153] + src40[154] + src40[155] + src40[156] + src40[157] + src40[158] + src40[159] + src40[160] + src40[161] + src40[162] + src40[163] + src40[164] + src40[165] + src40[166] + src40[167] + src40[168] + src40[169] + src40[170] + src40[171] + src40[172] + src40[173] + src40[174] + src40[175] + src40[176] + src40[177] + src40[178] + src40[179] + src40[180] + src40[181] + src40[182] + src40[183] + src40[184] + src40[185] + src40[186] + src40[187] + src40[188] + src40[189] + src40[190] + src40[191] + src40[192] + src40[193] + src40[194] + src40[195] + src40[196] + src40[197] + src40[198] + src40[199] + src40[200] + src40[201] + src40[202] + src40[203] + src40[204] + src40[205] + src40[206] + src40[207] + src40[208] + src40[209] + src40[210] + src40[211] + src40[212] + src40[213] + src40[214] + src40[215] + src40[216] + src40[217] + src40[218] + src40[219] + src40[220] + src40[221] + src40[222] + src40[223] + src40[224] + src40[225] + src40[226] + src40[227] + src40[228] + src40[229] + src40[230] + src40[231] + src40[232] + src40[233] + src40[234] + src40[235] + src40[236] + src40[237] + src40[238] + src40[239] + src40[240] + src40[241] + src40[242] + src40[243] + src40[244] + src40[245] + src40[246] + src40[247] + src40[248] + src40[249] + src40[250] + src40[251] + src40[252] + src40[253] + src40[254] + src40[255])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127] + src41[128] + src41[129] + src41[130] + src41[131] + src41[132] + src41[133] + src41[134] + src41[135] + src41[136] + src41[137] + src41[138] + src41[139] + src41[140] + src41[141] + src41[142] + src41[143] + src41[144] + src41[145] + src41[146] + src41[147] + src41[148] + src41[149] + src41[150] + src41[151] + src41[152] + src41[153] + src41[154] + src41[155] + src41[156] + src41[157] + src41[158] + src41[159] + src41[160] + src41[161] + src41[162] + src41[163] + src41[164] + src41[165] + src41[166] + src41[167] + src41[168] + src41[169] + src41[170] + src41[171] + src41[172] + src41[173] + src41[174] + src41[175] + src41[176] + src41[177] + src41[178] + src41[179] + src41[180] + src41[181] + src41[182] + src41[183] + src41[184] + src41[185] + src41[186] + src41[187] + src41[188] + src41[189] + src41[190] + src41[191] + src41[192] + src41[193] + src41[194] + src41[195] + src41[196] + src41[197] + src41[198] + src41[199] + src41[200] + src41[201] + src41[202] + src41[203] + src41[204] + src41[205] + src41[206] + src41[207] + src41[208] + src41[209] + src41[210] + src41[211] + src41[212] + src41[213] + src41[214] + src41[215] + src41[216] + src41[217] + src41[218] + src41[219] + src41[220] + src41[221] + src41[222] + src41[223] + src41[224] + src41[225] + src41[226] + src41[227] + src41[228] + src41[229] + src41[230] + src41[231] + src41[232] + src41[233] + src41[234] + src41[235] + src41[236] + src41[237] + src41[238] + src41[239] + src41[240] + src41[241] + src41[242] + src41[243] + src41[244] + src41[245] + src41[246] + src41[247] + src41[248] + src41[249] + src41[250] + src41[251] + src41[252] + src41[253] + src41[254] + src41[255])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127] + src42[128] + src42[129] + src42[130] + src42[131] + src42[132] + src42[133] + src42[134] + src42[135] + src42[136] + src42[137] + src42[138] + src42[139] + src42[140] + src42[141] + src42[142] + src42[143] + src42[144] + src42[145] + src42[146] + src42[147] + src42[148] + src42[149] + src42[150] + src42[151] + src42[152] + src42[153] + src42[154] + src42[155] + src42[156] + src42[157] + src42[158] + src42[159] + src42[160] + src42[161] + src42[162] + src42[163] + src42[164] + src42[165] + src42[166] + src42[167] + src42[168] + src42[169] + src42[170] + src42[171] + src42[172] + src42[173] + src42[174] + src42[175] + src42[176] + src42[177] + src42[178] + src42[179] + src42[180] + src42[181] + src42[182] + src42[183] + src42[184] + src42[185] + src42[186] + src42[187] + src42[188] + src42[189] + src42[190] + src42[191] + src42[192] + src42[193] + src42[194] + src42[195] + src42[196] + src42[197] + src42[198] + src42[199] + src42[200] + src42[201] + src42[202] + src42[203] + src42[204] + src42[205] + src42[206] + src42[207] + src42[208] + src42[209] + src42[210] + src42[211] + src42[212] + src42[213] + src42[214] + src42[215] + src42[216] + src42[217] + src42[218] + src42[219] + src42[220] + src42[221] + src42[222] + src42[223] + src42[224] + src42[225] + src42[226] + src42[227] + src42[228] + src42[229] + src42[230] + src42[231] + src42[232] + src42[233] + src42[234] + src42[235] + src42[236] + src42[237] + src42[238] + src42[239] + src42[240] + src42[241] + src42[242] + src42[243] + src42[244] + src42[245] + src42[246] + src42[247] + src42[248] + src42[249] + src42[250] + src42[251] + src42[252] + src42[253] + src42[254] + src42[255])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127] + src43[128] + src43[129] + src43[130] + src43[131] + src43[132] + src43[133] + src43[134] + src43[135] + src43[136] + src43[137] + src43[138] + src43[139] + src43[140] + src43[141] + src43[142] + src43[143] + src43[144] + src43[145] + src43[146] + src43[147] + src43[148] + src43[149] + src43[150] + src43[151] + src43[152] + src43[153] + src43[154] + src43[155] + src43[156] + src43[157] + src43[158] + src43[159] + src43[160] + src43[161] + src43[162] + src43[163] + src43[164] + src43[165] + src43[166] + src43[167] + src43[168] + src43[169] + src43[170] + src43[171] + src43[172] + src43[173] + src43[174] + src43[175] + src43[176] + src43[177] + src43[178] + src43[179] + src43[180] + src43[181] + src43[182] + src43[183] + src43[184] + src43[185] + src43[186] + src43[187] + src43[188] + src43[189] + src43[190] + src43[191] + src43[192] + src43[193] + src43[194] + src43[195] + src43[196] + src43[197] + src43[198] + src43[199] + src43[200] + src43[201] + src43[202] + src43[203] + src43[204] + src43[205] + src43[206] + src43[207] + src43[208] + src43[209] + src43[210] + src43[211] + src43[212] + src43[213] + src43[214] + src43[215] + src43[216] + src43[217] + src43[218] + src43[219] + src43[220] + src43[221] + src43[222] + src43[223] + src43[224] + src43[225] + src43[226] + src43[227] + src43[228] + src43[229] + src43[230] + src43[231] + src43[232] + src43[233] + src43[234] + src43[235] + src43[236] + src43[237] + src43[238] + src43[239] + src43[240] + src43[241] + src43[242] + src43[243] + src43[244] + src43[245] + src43[246] + src43[247] + src43[248] + src43[249] + src43[250] + src43[251] + src43[252] + src43[253] + src43[254] + src43[255])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127] + src44[128] + src44[129] + src44[130] + src44[131] + src44[132] + src44[133] + src44[134] + src44[135] + src44[136] + src44[137] + src44[138] + src44[139] + src44[140] + src44[141] + src44[142] + src44[143] + src44[144] + src44[145] + src44[146] + src44[147] + src44[148] + src44[149] + src44[150] + src44[151] + src44[152] + src44[153] + src44[154] + src44[155] + src44[156] + src44[157] + src44[158] + src44[159] + src44[160] + src44[161] + src44[162] + src44[163] + src44[164] + src44[165] + src44[166] + src44[167] + src44[168] + src44[169] + src44[170] + src44[171] + src44[172] + src44[173] + src44[174] + src44[175] + src44[176] + src44[177] + src44[178] + src44[179] + src44[180] + src44[181] + src44[182] + src44[183] + src44[184] + src44[185] + src44[186] + src44[187] + src44[188] + src44[189] + src44[190] + src44[191] + src44[192] + src44[193] + src44[194] + src44[195] + src44[196] + src44[197] + src44[198] + src44[199] + src44[200] + src44[201] + src44[202] + src44[203] + src44[204] + src44[205] + src44[206] + src44[207] + src44[208] + src44[209] + src44[210] + src44[211] + src44[212] + src44[213] + src44[214] + src44[215] + src44[216] + src44[217] + src44[218] + src44[219] + src44[220] + src44[221] + src44[222] + src44[223] + src44[224] + src44[225] + src44[226] + src44[227] + src44[228] + src44[229] + src44[230] + src44[231] + src44[232] + src44[233] + src44[234] + src44[235] + src44[236] + src44[237] + src44[238] + src44[239] + src44[240] + src44[241] + src44[242] + src44[243] + src44[244] + src44[245] + src44[246] + src44[247] + src44[248] + src44[249] + src44[250] + src44[251] + src44[252] + src44[253] + src44[254] + src44[255])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127] + src45[128] + src45[129] + src45[130] + src45[131] + src45[132] + src45[133] + src45[134] + src45[135] + src45[136] + src45[137] + src45[138] + src45[139] + src45[140] + src45[141] + src45[142] + src45[143] + src45[144] + src45[145] + src45[146] + src45[147] + src45[148] + src45[149] + src45[150] + src45[151] + src45[152] + src45[153] + src45[154] + src45[155] + src45[156] + src45[157] + src45[158] + src45[159] + src45[160] + src45[161] + src45[162] + src45[163] + src45[164] + src45[165] + src45[166] + src45[167] + src45[168] + src45[169] + src45[170] + src45[171] + src45[172] + src45[173] + src45[174] + src45[175] + src45[176] + src45[177] + src45[178] + src45[179] + src45[180] + src45[181] + src45[182] + src45[183] + src45[184] + src45[185] + src45[186] + src45[187] + src45[188] + src45[189] + src45[190] + src45[191] + src45[192] + src45[193] + src45[194] + src45[195] + src45[196] + src45[197] + src45[198] + src45[199] + src45[200] + src45[201] + src45[202] + src45[203] + src45[204] + src45[205] + src45[206] + src45[207] + src45[208] + src45[209] + src45[210] + src45[211] + src45[212] + src45[213] + src45[214] + src45[215] + src45[216] + src45[217] + src45[218] + src45[219] + src45[220] + src45[221] + src45[222] + src45[223] + src45[224] + src45[225] + src45[226] + src45[227] + src45[228] + src45[229] + src45[230] + src45[231] + src45[232] + src45[233] + src45[234] + src45[235] + src45[236] + src45[237] + src45[238] + src45[239] + src45[240] + src45[241] + src45[242] + src45[243] + src45[244] + src45[245] + src45[246] + src45[247] + src45[248] + src45[249] + src45[250] + src45[251] + src45[252] + src45[253] + src45[254] + src45[255])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127] + src46[128] + src46[129] + src46[130] + src46[131] + src46[132] + src46[133] + src46[134] + src46[135] + src46[136] + src46[137] + src46[138] + src46[139] + src46[140] + src46[141] + src46[142] + src46[143] + src46[144] + src46[145] + src46[146] + src46[147] + src46[148] + src46[149] + src46[150] + src46[151] + src46[152] + src46[153] + src46[154] + src46[155] + src46[156] + src46[157] + src46[158] + src46[159] + src46[160] + src46[161] + src46[162] + src46[163] + src46[164] + src46[165] + src46[166] + src46[167] + src46[168] + src46[169] + src46[170] + src46[171] + src46[172] + src46[173] + src46[174] + src46[175] + src46[176] + src46[177] + src46[178] + src46[179] + src46[180] + src46[181] + src46[182] + src46[183] + src46[184] + src46[185] + src46[186] + src46[187] + src46[188] + src46[189] + src46[190] + src46[191] + src46[192] + src46[193] + src46[194] + src46[195] + src46[196] + src46[197] + src46[198] + src46[199] + src46[200] + src46[201] + src46[202] + src46[203] + src46[204] + src46[205] + src46[206] + src46[207] + src46[208] + src46[209] + src46[210] + src46[211] + src46[212] + src46[213] + src46[214] + src46[215] + src46[216] + src46[217] + src46[218] + src46[219] + src46[220] + src46[221] + src46[222] + src46[223] + src46[224] + src46[225] + src46[226] + src46[227] + src46[228] + src46[229] + src46[230] + src46[231] + src46[232] + src46[233] + src46[234] + src46[235] + src46[236] + src46[237] + src46[238] + src46[239] + src46[240] + src46[241] + src46[242] + src46[243] + src46[244] + src46[245] + src46[246] + src46[247] + src46[248] + src46[249] + src46[250] + src46[251] + src46[252] + src46[253] + src46[254] + src46[255])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127] + src47[128] + src47[129] + src47[130] + src47[131] + src47[132] + src47[133] + src47[134] + src47[135] + src47[136] + src47[137] + src47[138] + src47[139] + src47[140] + src47[141] + src47[142] + src47[143] + src47[144] + src47[145] + src47[146] + src47[147] + src47[148] + src47[149] + src47[150] + src47[151] + src47[152] + src47[153] + src47[154] + src47[155] + src47[156] + src47[157] + src47[158] + src47[159] + src47[160] + src47[161] + src47[162] + src47[163] + src47[164] + src47[165] + src47[166] + src47[167] + src47[168] + src47[169] + src47[170] + src47[171] + src47[172] + src47[173] + src47[174] + src47[175] + src47[176] + src47[177] + src47[178] + src47[179] + src47[180] + src47[181] + src47[182] + src47[183] + src47[184] + src47[185] + src47[186] + src47[187] + src47[188] + src47[189] + src47[190] + src47[191] + src47[192] + src47[193] + src47[194] + src47[195] + src47[196] + src47[197] + src47[198] + src47[199] + src47[200] + src47[201] + src47[202] + src47[203] + src47[204] + src47[205] + src47[206] + src47[207] + src47[208] + src47[209] + src47[210] + src47[211] + src47[212] + src47[213] + src47[214] + src47[215] + src47[216] + src47[217] + src47[218] + src47[219] + src47[220] + src47[221] + src47[222] + src47[223] + src47[224] + src47[225] + src47[226] + src47[227] + src47[228] + src47[229] + src47[230] + src47[231] + src47[232] + src47[233] + src47[234] + src47[235] + src47[236] + src47[237] + src47[238] + src47[239] + src47[240] + src47[241] + src47[242] + src47[243] + src47[244] + src47[245] + src47[246] + src47[247] + src47[248] + src47[249] + src47[250] + src47[251] + src47[252] + src47[253] + src47[254] + src47[255])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127] + src48[128] + src48[129] + src48[130] + src48[131] + src48[132] + src48[133] + src48[134] + src48[135] + src48[136] + src48[137] + src48[138] + src48[139] + src48[140] + src48[141] + src48[142] + src48[143] + src48[144] + src48[145] + src48[146] + src48[147] + src48[148] + src48[149] + src48[150] + src48[151] + src48[152] + src48[153] + src48[154] + src48[155] + src48[156] + src48[157] + src48[158] + src48[159] + src48[160] + src48[161] + src48[162] + src48[163] + src48[164] + src48[165] + src48[166] + src48[167] + src48[168] + src48[169] + src48[170] + src48[171] + src48[172] + src48[173] + src48[174] + src48[175] + src48[176] + src48[177] + src48[178] + src48[179] + src48[180] + src48[181] + src48[182] + src48[183] + src48[184] + src48[185] + src48[186] + src48[187] + src48[188] + src48[189] + src48[190] + src48[191] + src48[192] + src48[193] + src48[194] + src48[195] + src48[196] + src48[197] + src48[198] + src48[199] + src48[200] + src48[201] + src48[202] + src48[203] + src48[204] + src48[205] + src48[206] + src48[207] + src48[208] + src48[209] + src48[210] + src48[211] + src48[212] + src48[213] + src48[214] + src48[215] + src48[216] + src48[217] + src48[218] + src48[219] + src48[220] + src48[221] + src48[222] + src48[223] + src48[224] + src48[225] + src48[226] + src48[227] + src48[228] + src48[229] + src48[230] + src48[231] + src48[232] + src48[233] + src48[234] + src48[235] + src48[236] + src48[237] + src48[238] + src48[239] + src48[240] + src48[241] + src48[242] + src48[243] + src48[244] + src48[245] + src48[246] + src48[247] + src48[248] + src48[249] + src48[250] + src48[251] + src48[252] + src48[253] + src48[254] + src48[255])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127] + src49[128] + src49[129] + src49[130] + src49[131] + src49[132] + src49[133] + src49[134] + src49[135] + src49[136] + src49[137] + src49[138] + src49[139] + src49[140] + src49[141] + src49[142] + src49[143] + src49[144] + src49[145] + src49[146] + src49[147] + src49[148] + src49[149] + src49[150] + src49[151] + src49[152] + src49[153] + src49[154] + src49[155] + src49[156] + src49[157] + src49[158] + src49[159] + src49[160] + src49[161] + src49[162] + src49[163] + src49[164] + src49[165] + src49[166] + src49[167] + src49[168] + src49[169] + src49[170] + src49[171] + src49[172] + src49[173] + src49[174] + src49[175] + src49[176] + src49[177] + src49[178] + src49[179] + src49[180] + src49[181] + src49[182] + src49[183] + src49[184] + src49[185] + src49[186] + src49[187] + src49[188] + src49[189] + src49[190] + src49[191] + src49[192] + src49[193] + src49[194] + src49[195] + src49[196] + src49[197] + src49[198] + src49[199] + src49[200] + src49[201] + src49[202] + src49[203] + src49[204] + src49[205] + src49[206] + src49[207] + src49[208] + src49[209] + src49[210] + src49[211] + src49[212] + src49[213] + src49[214] + src49[215] + src49[216] + src49[217] + src49[218] + src49[219] + src49[220] + src49[221] + src49[222] + src49[223] + src49[224] + src49[225] + src49[226] + src49[227] + src49[228] + src49[229] + src49[230] + src49[231] + src49[232] + src49[233] + src49[234] + src49[235] + src49[236] + src49[237] + src49[238] + src49[239] + src49[240] + src49[241] + src49[242] + src49[243] + src49[244] + src49[245] + src49[246] + src49[247] + src49[248] + src49[249] + src49[250] + src49[251] + src49[252] + src49[253] + src49[254] + src49[255])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127] + src50[128] + src50[129] + src50[130] + src50[131] + src50[132] + src50[133] + src50[134] + src50[135] + src50[136] + src50[137] + src50[138] + src50[139] + src50[140] + src50[141] + src50[142] + src50[143] + src50[144] + src50[145] + src50[146] + src50[147] + src50[148] + src50[149] + src50[150] + src50[151] + src50[152] + src50[153] + src50[154] + src50[155] + src50[156] + src50[157] + src50[158] + src50[159] + src50[160] + src50[161] + src50[162] + src50[163] + src50[164] + src50[165] + src50[166] + src50[167] + src50[168] + src50[169] + src50[170] + src50[171] + src50[172] + src50[173] + src50[174] + src50[175] + src50[176] + src50[177] + src50[178] + src50[179] + src50[180] + src50[181] + src50[182] + src50[183] + src50[184] + src50[185] + src50[186] + src50[187] + src50[188] + src50[189] + src50[190] + src50[191] + src50[192] + src50[193] + src50[194] + src50[195] + src50[196] + src50[197] + src50[198] + src50[199] + src50[200] + src50[201] + src50[202] + src50[203] + src50[204] + src50[205] + src50[206] + src50[207] + src50[208] + src50[209] + src50[210] + src50[211] + src50[212] + src50[213] + src50[214] + src50[215] + src50[216] + src50[217] + src50[218] + src50[219] + src50[220] + src50[221] + src50[222] + src50[223] + src50[224] + src50[225] + src50[226] + src50[227] + src50[228] + src50[229] + src50[230] + src50[231] + src50[232] + src50[233] + src50[234] + src50[235] + src50[236] + src50[237] + src50[238] + src50[239] + src50[240] + src50[241] + src50[242] + src50[243] + src50[244] + src50[245] + src50[246] + src50[247] + src50[248] + src50[249] + src50[250] + src50[251] + src50[252] + src50[253] + src50[254] + src50[255])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127] + src51[128] + src51[129] + src51[130] + src51[131] + src51[132] + src51[133] + src51[134] + src51[135] + src51[136] + src51[137] + src51[138] + src51[139] + src51[140] + src51[141] + src51[142] + src51[143] + src51[144] + src51[145] + src51[146] + src51[147] + src51[148] + src51[149] + src51[150] + src51[151] + src51[152] + src51[153] + src51[154] + src51[155] + src51[156] + src51[157] + src51[158] + src51[159] + src51[160] + src51[161] + src51[162] + src51[163] + src51[164] + src51[165] + src51[166] + src51[167] + src51[168] + src51[169] + src51[170] + src51[171] + src51[172] + src51[173] + src51[174] + src51[175] + src51[176] + src51[177] + src51[178] + src51[179] + src51[180] + src51[181] + src51[182] + src51[183] + src51[184] + src51[185] + src51[186] + src51[187] + src51[188] + src51[189] + src51[190] + src51[191] + src51[192] + src51[193] + src51[194] + src51[195] + src51[196] + src51[197] + src51[198] + src51[199] + src51[200] + src51[201] + src51[202] + src51[203] + src51[204] + src51[205] + src51[206] + src51[207] + src51[208] + src51[209] + src51[210] + src51[211] + src51[212] + src51[213] + src51[214] + src51[215] + src51[216] + src51[217] + src51[218] + src51[219] + src51[220] + src51[221] + src51[222] + src51[223] + src51[224] + src51[225] + src51[226] + src51[227] + src51[228] + src51[229] + src51[230] + src51[231] + src51[232] + src51[233] + src51[234] + src51[235] + src51[236] + src51[237] + src51[238] + src51[239] + src51[240] + src51[241] + src51[242] + src51[243] + src51[244] + src51[245] + src51[246] + src51[247] + src51[248] + src51[249] + src51[250] + src51[251] + src51[252] + src51[253] + src51[254] + src51[255])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127] + src52[128] + src52[129] + src52[130] + src52[131] + src52[132] + src52[133] + src52[134] + src52[135] + src52[136] + src52[137] + src52[138] + src52[139] + src52[140] + src52[141] + src52[142] + src52[143] + src52[144] + src52[145] + src52[146] + src52[147] + src52[148] + src52[149] + src52[150] + src52[151] + src52[152] + src52[153] + src52[154] + src52[155] + src52[156] + src52[157] + src52[158] + src52[159] + src52[160] + src52[161] + src52[162] + src52[163] + src52[164] + src52[165] + src52[166] + src52[167] + src52[168] + src52[169] + src52[170] + src52[171] + src52[172] + src52[173] + src52[174] + src52[175] + src52[176] + src52[177] + src52[178] + src52[179] + src52[180] + src52[181] + src52[182] + src52[183] + src52[184] + src52[185] + src52[186] + src52[187] + src52[188] + src52[189] + src52[190] + src52[191] + src52[192] + src52[193] + src52[194] + src52[195] + src52[196] + src52[197] + src52[198] + src52[199] + src52[200] + src52[201] + src52[202] + src52[203] + src52[204] + src52[205] + src52[206] + src52[207] + src52[208] + src52[209] + src52[210] + src52[211] + src52[212] + src52[213] + src52[214] + src52[215] + src52[216] + src52[217] + src52[218] + src52[219] + src52[220] + src52[221] + src52[222] + src52[223] + src52[224] + src52[225] + src52[226] + src52[227] + src52[228] + src52[229] + src52[230] + src52[231] + src52[232] + src52[233] + src52[234] + src52[235] + src52[236] + src52[237] + src52[238] + src52[239] + src52[240] + src52[241] + src52[242] + src52[243] + src52[244] + src52[245] + src52[246] + src52[247] + src52[248] + src52[249] + src52[250] + src52[251] + src52[252] + src52[253] + src52[254] + src52[255])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127] + src53[128] + src53[129] + src53[130] + src53[131] + src53[132] + src53[133] + src53[134] + src53[135] + src53[136] + src53[137] + src53[138] + src53[139] + src53[140] + src53[141] + src53[142] + src53[143] + src53[144] + src53[145] + src53[146] + src53[147] + src53[148] + src53[149] + src53[150] + src53[151] + src53[152] + src53[153] + src53[154] + src53[155] + src53[156] + src53[157] + src53[158] + src53[159] + src53[160] + src53[161] + src53[162] + src53[163] + src53[164] + src53[165] + src53[166] + src53[167] + src53[168] + src53[169] + src53[170] + src53[171] + src53[172] + src53[173] + src53[174] + src53[175] + src53[176] + src53[177] + src53[178] + src53[179] + src53[180] + src53[181] + src53[182] + src53[183] + src53[184] + src53[185] + src53[186] + src53[187] + src53[188] + src53[189] + src53[190] + src53[191] + src53[192] + src53[193] + src53[194] + src53[195] + src53[196] + src53[197] + src53[198] + src53[199] + src53[200] + src53[201] + src53[202] + src53[203] + src53[204] + src53[205] + src53[206] + src53[207] + src53[208] + src53[209] + src53[210] + src53[211] + src53[212] + src53[213] + src53[214] + src53[215] + src53[216] + src53[217] + src53[218] + src53[219] + src53[220] + src53[221] + src53[222] + src53[223] + src53[224] + src53[225] + src53[226] + src53[227] + src53[228] + src53[229] + src53[230] + src53[231] + src53[232] + src53[233] + src53[234] + src53[235] + src53[236] + src53[237] + src53[238] + src53[239] + src53[240] + src53[241] + src53[242] + src53[243] + src53[244] + src53[245] + src53[246] + src53[247] + src53[248] + src53[249] + src53[250] + src53[251] + src53[252] + src53[253] + src53[254] + src53[255])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127] + src54[128] + src54[129] + src54[130] + src54[131] + src54[132] + src54[133] + src54[134] + src54[135] + src54[136] + src54[137] + src54[138] + src54[139] + src54[140] + src54[141] + src54[142] + src54[143] + src54[144] + src54[145] + src54[146] + src54[147] + src54[148] + src54[149] + src54[150] + src54[151] + src54[152] + src54[153] + src54[154] + src54[155] + src54[156] + src54[157] + src54[158] + src54[159] + src54[160] + src54[161] + src54[162] + src54[163] + src54[164] + src54[165] + src54[166] + src54[167] + src54[168] + src54[169] + src54[170] + src54[171] + src54[172] + src54[173] + src54[174] + src54[175] + src54[176] + src54[177] + src54[178] + src54[179] + src54[180] + src54[181] + src54[182] + src54[183] + src54[184] + src54[185] + src54[186] + src54[187] + src54[188] + src54[189] + src54[190] + src54[191] + src54[192] + src54[193] + src54[194] + src54[195] + src54[196] + src54[197] + src54[198] + src54[199] + src54[200] + src54[201] + src54[202] + src54[203] + src54[204] + src54[205] + src54[206] + src54[207] + src54[208] + src54[209] + src54[210] + src54[211] + src54[212] + src54[213] + src54[214] + src54[215] + src54[216] + src54[217] + src54[218] + src54[219] + src54[220] + src54[221] + src54[222] + src54[223] + src54[224] + src54[225] + src54[226] + src54[227] + src54[228] + src54[229] + src54[230] + src54[231] + src54[232] + src54[233] + src54[234] + src54[235] + src54[236] + src54[237] + src54[238] + src54[239] + src54[240] + src54[241] + src54[242] + src54[243] + src54[244] + src54[245] + src54[246] + src54[247] + src54[248] + src54[249] + src54[250] + src54[251] + src54[252] + src54[253] + src54[254] + src54[255])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127] + src55[128] + src55[129] + src55[130] + src55[131] + src55[132] + src55[133] + src55[134] + src55[135] + src55[136] + src55[137] + src55[138] + src55[139] + src55[140] + src55[141] + src55[142] + src55[143] + src55[144] + src55[145] + src55[146] + src55[147] + src55[148] + src55[149] + src55[150] + src55[151] + src55[152] + src55[153] + src55[154] + src55[155] + src55[156] + src55[157] + src55[158] + src55[159] + src55[160] + src55[161] + src55[162] + src55[163] + src55[164] + src55[165] + src55[166] + src55[167] + src55[168] + src55[169] + src55[170] + src55[171] + src55[172] + src55[173] + src55[174] + src55[175] + src55[176] + src55[177] + src55[178] + src55[179] + src55[180] + src55[181] + src55[182] + src55[183] + src55[184] + src55[185] + src55[186] + src55[187] + src55[188] + src55[189] + src55[190] + src55[191] + src55[192] + src55[193] + src55[194] + src55[195] + src55[196] + src55[197] + src55[198] + src55[199] + src55[200] + src55[201] + src55[202] + src55[203] + src55[204] + src55[205] + src55[206] + src55[207] + src55[208] + src55[209] + src55[210] + src55[211] + src55[212] + src55[213] + src55[214] + src55[215] + src55[216] + src55[217] + src55[218] + src55[219] + src55[220] + src55[221] + src55[222] + src55[223] + src55[224] + src55[225] + src55[226] + src55[227] + src55[228] + src55[229] + src55[230] + src55[231] + src55[232] + src55[233] + src55[234] + src55[235] + src55[236] + src55[237] + src55[238] + src55[239] + src55[240] + src55[241] + src55[242] + src55[243] + src55[244] + src55[245] + src55[246] + src55[247] + src55[248] + src55[249] + src55[250] + src55[251] + src55[252] + src55[253] + src55[254] + src55[255])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127] + src56[128] + src56[129] + src56[130] + src56[131] + src56[132] + src56[133] + src56[134] + src56[135] + src56[136] + src56[137] + src56[138] + src56[139] + src56[140] + src56[141] + src56[142] + src56[143] + src56[144] + src56[145] + src56[146] + src56[147] + src56[148] + src56[149] + src56[150] + src56[151] + src56[152] + src56[153] + src56[154] + src56[155] + src56[156] + src56[157] + src56[158] + src56[159] + src56[160] + src56[161] + src56[162] + src56[163] + src56[164] + src56[165] + src56[166] + src56[167] + src56[168] + src56[169] + src56[170] + src56[171] + src56[172] + src56[173] + src56[174] + src56[175] + src56[176] + src56[177] + src56[178] + src56[179] + src56[180] + src56[181] + src56[182] + src56[183] + src56[184] + src56[185] + src56[186] + src56[187] + src56[188] + src56[189] + src56[190] + src56[191] + src56[192] + src56[193] + src56[194] + src56[195] + src56[196] + src56[197] + src56[198] + src56[199] + src56[200] + src56[201] + src56[202] + src56[203] + src56[204] + src56[205] + src56[206] + src56[207] + src56[208] + src56[209] + src56[210] + src56[211] + src56[212] + src56[213] + src56[214] + src56[215] + src56[216] + src56[217] + src56[218] + src56[219] + src56[220] + src56[221] + src56[222] + src56[223] + src56[224] + src56[225] + src56[226] + src56[227] + src56[228] + src56[229] + src56[230] + src56[231] + src56[232] + src56[233] + src56[234] + src56[235] + src56[236] + src56[237] + src56[238] + src56[239] + src56[240] + src56[241] + src56[242] + src56[243] + src56[244] + src56[245] + src56[246] + src56[247] + src56[248] + src56[249] + src56[250] + src56[251] + src56[252] + src56[253] + src56[254] + src56[255])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127] + src57[128] + src57[129] + src57[130] + src57[131] + src57[132] + src57[133] + src57[134] + src57[135] + src57[136] + src57[137] + src57[138] + src57[139] + src57[140] + src57[141] + src57[142] + src57[143] + src57[144] + src57[145] + src57[146] + src57[147] + src57[148] + src57[149] + src57[150] + src57[151] + src57[152] + src57[153] + src57[154] + src57[155] + src57[156] + src57[157] + src57[158] + src57[159] + src57[160] + src57[161] + src57[162] + src57[163] + src57[164] + src57[165] + src57[166] + src57[167] + src57[168] + src57[169] + src57[170] + src57[171] + src57[172] + src57[173] + src57[174] + src57[175] + src57[176] + src57[177] + src57[178] + src57[179] + src57[180] + src57[181] + src57[182] + src57[183] + src57[184] + src57[185] + src57[186] + src57[187] + src57[188] + src57[189] + src57[190] + src57[191] + src57[192] + src57[193] + src57[194] + src57[195] + src57[196] + src57[197] + src57[198] + src57[199] + src57[200] + src57[201] + src57[202] + src57[203] + src57[204] + src57[205] + src57[206] + src57[207] + src57[208] + src57[209] + src57[210] + src57[211] + src57[212] + src57[213] + src57[214] + src57[215] + src57[216] + src57[217] + src57[218] + src57[219] + src57[220] + src57[221] + src57[222] + src57[223] + src57[224] + src57[225] + src57[226] + src57[227] + src57[228] + src57[229] + src57[230] + src57[231] + src57[232] + src57[233] + src57[234] + src57[235] + src57[236] + src57[237] + src57[238] + src57[239] + src57[240] + src57[241] + src57[242] + src57[243] + src57[244] + src57[245] + src57[246] + src57[247] + src57[248] + src57[249] + src57[250] + src57[251] + src57[252] + src57[253] + src57[254] + src57[255])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127] + src58[128] + src58[129] + src58[130] + src58[131] + src58[132] + src58[133] + src58[134] + src58[135] + src58[136] + src58[137] + src58[138] + src58[139] + src58[140] + src58[141] + src58[142] + src58[143] + src58[144] + src58[145] + src58[146] + src58[147] + src58[148] + src58[149] + src58[150] + src58[151] + src58[152] + src58[153] + src58[154] + src58[155] + src58[156] + src58[157] + src58[158] + src58[159] + src58[160] + src58[161] + src58[162] + src58[163] + src58[164] + src58[165] + src58[166] + src58[167] + src58[168] + src58[169] + src58[170] + src58[171] + src58[172] + src58[173] + src58[174] + src58[175] + src58[176] + src58[177] + src58[178] + src58[179] + src58[180] + src58[181] + src58[182] + src58[183] + src58[184] + src58[185] + src58[186] + src58[187] + src58[188] + src58[189] + src58[190] + src58[191] + src58[192] + src58[193] + src58[194] + src58[195] + src58[196] + src58[197] + src58[198] + src58[199] + src58[200] + src58[201] + src58[202] + src58[203] + src58[204] + src58[205] + src58[206] + src58[207] + src58[208] + src58[209] + src58[210] + src58[211] + src58[212] + src58[213] + src58[214] + src58[215] + src58[216] + src58[217] + src58[218] + src58[219] + src58[220] + src58[221] + src58[222] + src58[223] + src58[224] + src58[225] + src58[226] + src58[227] + src58[228] + src58[229] + src58[230] + src58[231] + src58[232] + src58[233] + src58[234] + src58[235] + src58[236] + src58[237] + src58[238] + src58[239] + src58[240] + src58[241] + src58[242] + src58[243] + src58[244] + src58[245] + src58[246] + src58[247] + src58[248] + src58[249] + src58[250] + src58[251] + src58[252] + src58[253] + src58[254] + src58[255])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127] + src59[128] + src59[129] + src59[130] + src59[131] + src59[132] + src59[133] + src59[134] + src59[135] + src59[136] + src59[137] + src59[138] + src59[139] + src59[140] + src59[141] + src59[142] + src59[143] + src59[144] + src59[145] + src59[146] + src59[147] + src59[148] + src59[149] + src59[150] + src59[151] + src59[152] + src59[153] + src59[154] + src59[155] + src59[156] + src59[157] + src59[158] + src59[159] + src59[160] + src59[161] + src59[162] + src59[163] + src59[164] + src59[165] + src59[166] + src59[167] + src59[168] + src59[169] + src59[170] + src59[171] + src59[172] + src59[173] + src59[174] + src59[175] + src59[176] + src59[177] + src59[178] + src59[179] + src59[180] + src59[181] + src59[182] + src59[183] + src59[184] + src59[185] + src59[186] + src59[187] + src59[188] + src59[189] + src59[190] + src59[191] + src59[192] + src59[193] + src59[194] + src59[195] + src59[196] + src59[197] + src59[198] + src59[199] + src59[200] + src59[201] + src59[202] + src59[203] + src59[204] + src59[205] + src59[206] + src59[207] + src59[208] + src59[209] + src59[210] + src59[211] + src59[212] + src59[213] + src59[214] + src59[215] + src59[216] + src59[217] + src59[218] + src59[219] + src59[220] + src59[221] + src59[222] + src59[223] + src59[224] + src59[225] + src59[226] + src59[227] + src59[228] + src59[229] + src59[230] + src59[231] + src59[232] + src59[233] + src59[234] + src59[235] + src59[236] + src59[237] + src59[238] + src59[239] + src59[240] + src59[241] + src59[242] + src59[243] + src59[244] + src59[245] + src59[246] + src59[247] + src59[248] + src59[249] + src59[250] + src59[251] + src59[252] + src59[253] + src59[254] + src59[255])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127] + src60[128] + src60[129] + src60[130] + src60[131] + src60[132] + src60[133] + src60[134] + src60[135] + src60[136] + src60[137] + src60[138] + src60[139] + src60[140] + src60[141] + src60[142] + src60[143] + src60[144] + src60[145] + src60[146] + src60[147] + src60[148] + src60[149] + src60[150] + src60[151] + src60[152] + src60[153] + src60[154] + src60[155] + src60[156] + src60[157] + src60[158] + src60[159] + src60[160] + src60[161] + src60[162] + src60[163] + src60[164] + src60[165] + src60[166] + src60[167] + src60[168] + src60[169] + src60[170] + src60[171] + src60[172] + src60[173] + src60[174] + src60[175] + src60[176] + src60[177] + src60[178] + src60[179] + src60[180] + src60[181] + src60[182] + src60[183] + src60[184] + src60[185] + src60[186] + src60[187] + src60[188] + src60[189] + src60[190] + src60[191] + src60[192] + src60[193] + src60[194] + src60[195] + src60[196] + src60[197] + src60[198] + src60[199] + src60[200] + src60[201] + src60[202] + src60[203] + src60[204] + src60[205] + src60[206] + src60[207] + src60[208] + src60[209] + src60[210] + src60[211] + src60[212] + src60[213] + src60[214] + src60[215] + src60[216] + src60[217] + src60[218] + src60[219] + src60[220] + src60[221] + src60[222] + src60[223] + src60[224] + src60[225] + src60[226] + src60[227] + src60[228] + src60[229] + src60[230] + src60[231] + src60[232] + src60[233] + src60[234] + src60[235] + src60[236] + src60[237] + src60[238] + src60[239] + src60[240] + src60[241] + src60[242] + src60[243] + src60[244] + src60[245] + src60[246] + src60[247] + src60[248] + src60[249] + src60[250] + src60[251] + src60[252] + src60[253] + src60[254] + src60[255])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127] + src61[128] + src61[129] + src61[130] + src61[131] + src61[132] + src61[133] + src61[134] + src61[135] + src61[136] + src61[137] + src61[138] + src61[139] + src61[140] + src61[141] + src61[142] + src61[143] + src61[144] + src61[145] + src61[146] + src61[147] + src61[148] + src61[149] + src61[150] + src61[151] + src61[152] + src61[153] + src61[154] + src61[155] + src61[156] + src61[157] + src61[158] + src61[159] + src61[160] + src61[161] + src61[162] + src61[163] + src61[164] + src61[165] + src61[166] + src61[167] + src61[168] + src61[169] + src61[170] + src61[171] + src61[172] + src61[173] + src61[174] + src61[175] + src61[176] + src61[177] + src61[178] + src61[179] + src61[180] + src61[181] + src61[182] + src61[183] + src61[184] + src61[185] + src61[186] + src61[187] + src61[188] + src61[189] + src61[190] + src61[191] + src61[192] + src61[193] + src61[194] + src61[195] + src61[196] + src61[197] + src61[198] + src61[199] + src61[200] + src61[201] + src61[202] + src61[203] + src61[204] + src61[205] + src61[206] + src61[207] + src61[208] + src61[209] + src61[210] + src61[211] + src61[212] + src61[213] + src61[214] + src61[215] + src61[216] + src61[217] + src61[218] + src61[219] + src61[220] + src61[221] + src61[222] + src61[223] + src61[224] + src61[225] + src61[226] + src61[227] + src61[228] + src61[229] + src61[230] + src61[231] + src61[232] + src61[233] + src61[234] + src61[235] + src61[236] + src61[237] + src61[238] + src61[239] + src61[240] + src61[241] + src61[242] + src61[243] + src61[244] + src61[245] + src61[246] + src61[247] + src61[248] + src61[249] + src61[250] + src61[251] + src61[252] + src61[253] + src61[254] + src61[255])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127] + src62[128] + src62[129] + src62[130] + src62[131] + src62[132] + src62[133] + src62[134] + src62[135] + src62[136] + src62[137] + src62[138] + src62[139] + src62[140] + src62[141] + src62[142] + src62[143] + src62[144] + src62[145] + src62[146] + src62[147] + src62[148] + src62[149] + src62[150] + src62[151] + src62[152] + src62[153] + src62[154] + src62[155] + src62[156] + src62[157] + src62[158] + src62[159] + src62[160] + src62[161] + src62[162] + src62[163] + src62[164] + src62[165] + src62[166] + src62[167] + src62[168] + src62[169] + src62[170] + src62[171] + src62[172] + src62[173] + src62[174] + src62[175] + src62[176] + src62[177] + src62[178] + src62[179] + src62[180] + src62[181] + src62[182] + src62[183] + src62[184] + src62[185] + src62[186] + src62[187] + src62[188] + src62[189] + src62[190] + src62[191] + src62[192] + src62[193] + src62[194] + src62[195] + src62[196] + src62[197] + src62[198] + src62[199] + src62[200] + src62[201] + src62[202] + src62[203] + src62[204] + src62[205] + src62[206] + src62[207] + src62[208] + src62[209] + src62[210] + src62[211] + src62[212] + src62[213] + src62[214] + src62[215] + src62[216] + src62[217] + src62[218] + src62[219] + src62[220] + src62[221] + src62[222] + src62[223] + src62[224] + src62[225] + src62[226] + src62[227] + src62[228] + src62[229] + src62[230] + src62[231] + src62[232] + src62[233] + src62[234] + src62[235] + src62[236] + src62[237] + src62[238] + src62[239] + src62[240] + src62[241] + src62[242] + src62[243] + src62[244] + src62[245] + src62[246] + src62[247] + src62[248] + src62[249] + src62[250] + src62[251] + src62[252] + src62[253] + src62[254] + src62[255])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127] + src63[128] + src63[129] + src63[130] + src63[131] + src63[132] + src63[133] + src63[134] + src63[135] + src63[136] + src63[137] + src63[138] + src63[139] + src63[140] + src63[141] + src63[142] + src63[143] + src63[144] + src63[145] + src63[146] + src63[147] + src63[148] + src63[149] + src63[150] + src63[151] + src63[152] + src63[153] + src63[154] + src63[155] + src63[156] + src63[157] + src63[158] + src63[159] + src63[160] + src63[161] + src63[162] + src63[163] + src63[164] + src63[165] + src63[166] + src63[167] + src63[168] + src63[169] + src63[170] + src63[171] + src63[172] + src63[173] + src63[174] + src63[175] + src63[176] + src63[177] + src63[178] + src63[179] + src63[180] + src63[181] + src63[182] + src63[183] + src63[184] + src63[185] + src63[186] + src63[187] + src63[188] + src63[189] + src63[190] + src63[191] + src63[192] + src63[193] + src63[194] + src63[195] + src63[196] + src63[197] + src63[198] + src63[199] + src63[200] + src63[201] + src63[202] + src63[203] + src63[204] + src63[205] + src63[206] + src63[207] + src63[208] + src63[209] + src63[210] + src63[211] + src63[212] + src63[213] + src63[214] + src63[215] + src63[216] + src63[217] + src63[218] + src63[219] + src63[220] + src63[221] + src63[222] + src63[223] + src63[224] + src63[225] + src63[226] + src63[227] + src63[228] + src63[229] + src63[230] + src63[231] + src63[232] + src63[233] + src63[234] + src63[235] + src63[236] + src63[237] + src63[238] + src63[239] + src63[240] + src63[241] + src63[242] + src63[243] + src63[244] + src63[245] + src63[246] + src63[247] + src63[248] + src63[249] + src63[250] + src63[251] + src63[252] + src63[253] + src63[254] + src63[255])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70) + ((dst71[0])<<71);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4e05706c61b65b4cf05c2a64935184e7f5a27e012903cea11fe531762b67cc0d8cf683ce2296fb00e0cde1d9b4c9e98176320f7e0949d60cc94154f0eb88a9046c38d2fe476dca2b280836ea79c9d017ae15c42d7172a57a85df7f38f50bb16f9250622004aada0d942b5780fd5cab9f0adc2562236a4ad863a7b620f125cf2b25e4cc9da3e1ef852379eeba3bfff168336f7b0efc468060c546a4b10609dc37b2cab6879ecbd3553f7069279357a7b1bdfa8b51bf2687e85e09096c30f933ba72512e109d86cf7485b5e40686c601ec954877d8dd22f08ba798752a72859f57f1667f6682b4be1d20c52db9822434b8a144898f36abb86fae5c8a6e895ea79e4bed829d0f86f3a72953322fdb9335212afac35fefc4ea0caa965eeb723787eeb1f9bc31729302c1844ac5edefae24ab5fe3e2827d9c4071e92e45e28f6afeb15673f44f7cb0f8f1d40d8be0bcf83375eba78870e56473b7cdf9c90b8d9a2608be493c3572276b5e2ed4bc7a59902e78439d94173b3a47e0307d5280abf9428a34a6c0924bd07a348d627ec9e0503f7a4f6b2e7faa7bf2172d1ab3e75e64a8a49c14ffd97e7b114fd17a020c637447a281f92f305a62dac9b0400505829826d38a032a65c297dadf7ce48bdcfcfa49216c839286c91c7874801863294e05e6f2e3a9a21a6469ea301dd8d5b15d19473e212178090f4139682617d9542bdf2f6746e0890c80b769a5e2ffc03222001509d785aac01013411488e505f498cb689f884e7675aa0e47cd18cc94c667aa135ea6764fd7de020a378054765b9878c8ae3c9b80e3a595107db9af79d9ac29d5a3b4451c3bf15b81c7dca6c8714f6143aa475b56548e505fb42de8f2fd2f5a2ee53dd682b1346ad320989c316f31c46e4e71525fa70e167c682420ebe1f66fa470f0f2f71938a047f163971e8827415377ebd2bed608fc286d4fb96a5a535d36afb5f5c25c316217e94c77158d3b2787630eb764cb67a30c0585b613cd7ac8f729dee716fa15d5f15a0d04b02b8004fbf566901a82bfad7f23e1ce67ea655559b63337caba41d84aedb6f3540aa441842e6d6f7d8bda28205208e48beabceb850189ea62fda384155f007e039545720adff6e111b782d04a8497cec37b6d4d35ebbed38a847d7e04c4d15224bd916cff20ebe5e6da90f8ac9459b68c13d8a9bc400abcc9fa3f583762e95bdd7706ad0225f0bd881dc31f6d1e89b4e9ea40cb5e793dbad860505e3d06e6236c2eca6dfbfaa83fd19892ffdf12782fd603669495796c1819c116fd59764beeb4dbe348eeea913e5094aff219d65a8da3329674caeb42573f58ab6a00bc48c00f547da03327d1ae33cb1d386391534a012364ce9fddd55108cb1aa0604ae7252f816f9f282db03bc5a75f71045b2c9e36c81c2d3f55b9cffe1f2c39a5351563ccc5c0b134930a8e4f8ddc210afdd76fd44564e875190bb9805319689cb70f99639a8e7bb7b535160d8c2fca953fdddd1bb1d74d0204a717bb454029a57882efe38974b8b8e328d232dba8b36ce05bb55ef86f43e2c1e29c0add1046e4f40a18a93f05ba69732c03432ac5e555cb3087e7130f17e27977cfd2d6737864f497e26b2d359ddc254ba853ced989d9efdc49d155a3e2dbcb49e6a6456788ab8755fd56511be9aa8688129cd2d5563df3f8a3d3668b24df6cc3ed8b6961db5c2125e2b75f9217dec716263946ed412eeac140830afe025ae9415d7a16e6bc6e3fe8351e03b94051f269e35bb6c00da412da57c1a54368fa75ea6a0ad4550f4597dcb146ad10cbf278898ed9cc7c27a4b4219ab2bb3b7941d87fdee72497891f20b36e4854f8f2d974d78b16bddd41f60fbd276cf779dd0b05d706568989d53b95c295cbcd0cdf50a53d9a5f849b8430a3efab13ebce76765768e6a96aeb6ee7caa67e1d85e0a6d1dc8695b917e674d77fd99d580f14d106bdc8b23a9ce39e81fe85c2e7899ff56f72e7848e4aac66e87bfa96e3338eddd91f73ed58e6f057c51ba47ba77d6fdc41ac99cbd3859d8bd9aea1df74f8622d447c9c02825f79e5aafb10a76a36b4837f243d32ee633a1fce274ffe37dc1621e85ed8c2bba9b3b756f328f127c5018cb289d8d9f5ff005a268a056889a7c31d274c2566af89fd94e9ec6c59cfade033ae39ab3568db05e2cf12d2b3e81f9228333bf551a64b75ef6e80d9eb0e27db32a07e651e26f610c71e09f00e7d0d8bf3e0258fbdbecdbb5399d31563364fe4bba92f7534c8f643435780d3c2703b8eba815d042e9096160683a1b2b25890ebdf46acfd8762844bfc97768203bab176449de9e334f90101c65616e0d910d9f719998a1fae73d354df6b12395cc20d181e46465bc9fd931ba8bcaba322126d7794cd2c7d2dc53bdd9ec9686a48616e356ab834182fea68c411ac5e48215f2bf0c5ec0c53c405f4eda3a27c87de4d1fdf4069e40704315d1285aae0daac329b8afe72bb1a2c1c1f41510060f6281c9b7d3124c9044e6123feae46de32e0b38272776f805eb27dd76a3eb7c39828aa8d91772e7ab57e72dc9970aa35d6ab792b48ed86be34f4811289b41bff670b2610269fdf9ff15e57e68975853c6d9408ca95a0a07da01e1f8fb06f83aec02331e57a9621244b75c58458e00876ec31ae1b83661cee2eebc34b3bca4bb0f5724228d2661175291c7a16ccced6ea88a05761ebd3718259e3b74101243af40bfc045eabf43e7bc300c780120c6eb2c374556d57398f9f6efef2b954ea5d4dca178f7596ea18dc5cd0aeefd1735d7dabf12241793443dd33527d4115f5dbbf83c25606ec2336c7b507e6aae02b88a450c22ed92c6a3d3ef930f5873f001fb6c22ecee874d822b66bfb7a47bed01a47e59a3fcb199e1c7c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd2664388c5e6d93745cfa1ee5ba2ffc40c5bfc3941537c42262b2d015ecba778ed301489105ec354e683e96ae1ad67b5a3ba40432d859ce8c52ea6ea3d8896ffbaf4babeb59c600fa3b1a56d2b1fbf622bb1afcbeb26460431d56c83245603f7d733b9dd010a8365f8726f8c26ca0688332d20bdfe279379a9d1e276a237434a601ef81e2d0a99122e1bdf325a06c43a3e291a51a7e97660c2189252afca40dabd2b627450cab19bf7cf208b3299ec5bfcc6f0b1a5ecbc20c96315b2a234ad250dd0862737c4d1ecbae3b0f4d6d5ff22ce42ae12896635762409028074c40a44c43c50f92ba5c0a5019a4d5fa70c30ebc504952d50d94742a32aeb8345b2aebbbc24f6d5f8273d6682e1667989c4c0fced75674ba249e490abf120033d6795a9be11d9ce6e33dbb8c514ba8b9aba60d1b4f4027399e85aa14352f2f84b7f934854710824cd054d44ea037aa9a399831005e9ffc54cf833002a7cc5cbfbee81d76c1ce709127543e7d77b79de39e7071d41ceac3f6ddd69be86cc19894c4e40e84046d0752bbc48a4ef7d04033b445657e5f65c432b9510ce8e24b6de42a48e53f50186faaab24577f4a9381f69353eea92fb1b1459359f6bb261b8b303f8b819c8730b7b9ae37eacad3042f49b68517e549635600a941fc6b420f1b0ccb6573328dd1d1d233f81c5253d691504a9c73704bc0fc50a50e50fb61cfebe8130334b71691183374ea28a7079364374aeaac69450adfb4f24e64aa362f43bb43dec7a1ae41f00269f9b33a528b931df6ced1442082d641779e71ae50a21c2891a8e9dbbaa26b2e47b3a78c21b0aa0c5fc41c80e7346eb69a2f7c3c5d387689a62d6b75de78213127fd4e18c2a074f8647086a6eaaaea2739ba85cd7fa6d65d03f9da578e8ebb59e1f6bfa756ed9f722d37467ac086cbcf6ed069cdc424512214daa9ab874dfc898357b765a47e188cbe7760243600df6f9ac43bfc1314170f6a94878e2eb3901db9c664fdf6457554cf9913f1748e49763b7b512a8b1c3f86c3c24cf644ce6563f9a4645b882dd39de10529285eb46b81b4e60ab991316c91fbfdc977c30cd66f60d0197361df0b0e53bc389c6702c987387c24c59f720487c7e66b6c14ffdf87b813085b561799bf4fed9d2c34f8347b8a4a417405f8441e7a40eb27789b9803310f8b1b81a5ce347468340489ebe40bf85fbc8558f13d3f9ad4a16e9dd8d4ee665348fdf5c9e12881eb6969abf002e04373ce71f1c785b1740078279914363aeac329c291902e7af11931556452dda3415ffdc24e047fe1322b758bb2857f009aafc0656b305944a88c917214798b925ba5f7bd16f2a4c1b1087df86c8fa8c8d37895e146d225288b2c737f9edbded44b0a5ffe517be6429d57b6e54585a5b6bccd099fe8bea9c35b2e6d09058c35d9f5131a7c40e3772fd5ed6c4b953a55e92299b60778410258a178bd2927a5409e2e1f3c894887ffd0462cc944ee6b4bfcdb6240b3ee698c08957513e99104578c209de5f856160ae7f48e311e2301141300ab4615dc3cf0440abe68c4bb589635b467080b655da18e63f307b503c811034de16f45424491b46af429736b2aae697bcd979392a5f466a5102dcc947d472aa89c6b7838f24b6e3214139d8be84666a0947fb31734730204723e96fc4979af611953d8c8ccdb135b15f6f5dff5aa93918502e5c34713d7228da4c0a04c1d0d0d33a0881aacbb07b6be1aa39aeccf5eada4dbcffd43227f4404b6d37f2738713e888bc76af5df21e69fe0f758c1ebd8e14245cc6c2346ce37a9795f60b2768502a924ad7bd7596fd1f256ead89a2e214b215483491bf8326700cc507f3509f14afe2ae0e1cdba41e5bdc3ffa154927e92ff99b4d7e2cc4d9d04c429ea983e853645317fe7ee076c4d5d393a97da6fecad5a661cade78edd3c96b545769e54868de7cfc2f6e10088a94916b798ae0abcaf4cdd9510d8286f3ddedea87f1e9135c251340a86e26a36374e76bfd4e5db6b87960cf5090eaa1b54846cd3132c9e5ca23073d85dcd1998a3fb1a51614e3ef2b67df1fac14c4049114cf8045de0d52c4e797395f189e1b507487013ad8dc113275635ba313c9a6216483125c96643c53ef2177262ef26cf2db6d6c5899c4327610910347b4c3326e7cbbc0b861829753873f147e73c14d9ab61c7fbe670390a040c44aee985d31fdc85030e0ad6987fa87ef53db0cb3a8e3870e6c6bf62c35a58d9e3e2cc5d4df57777f32ebfc2977fae0ba71362daaaa974fe42c895c78e18acdfa752a66a5719f676e995e12537e54b8dc10723dad9bfd994d3a1c03a2423fa6a80b8c587877b43f957e9f2ac9f64eb3dd35a49679e20443cb4db61850e7f40bfd0ab9ab48b18a311ef11ea45d79188c6344bef97984fc218ff9bd153757f18f1d5b9eaacd249726d23f258072a09854b81e56b6196fab0275d7099872b71cd8fa5257af9936ba32d1e4126dca6bacffb21969fe238a9198f4e5a0b368c0d67a84bed719900860aa7a5c5ee75d5ef44662939789931cc604bcf4f28f67e93c91680ba99bf7e1e484fa33b172466a9dff75f4496b53d26617e698063f6ae927a4a24028ff2052c85d2f4f0f8a4d8422467ceebd9292e0e14b4553330a09f391f8c75e50d59300600eef3168179c50e343873bdefe1d2323a139295c7fb707102a350afed213b4b768a58835ecad59452eea6401b7b734c11631b6d1b11e5378fa6de86f167a412283ac5a967895be3ac5f7c484f883480cac9e507e419f1766b593f03cca9c2720b7ddad6fa7ccc8638638047bc8478fb70fbe7fbcdbded8393fe4ae9cbcc770002949e5e8b48db77041d00a6e102590aa2d8b4268d2d210f435a00ef500d903381d201;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h67178e5696b779d7a29bf9d3ab8ccc1df32e42dc2ba7d085048695cb79a54fa01cdc7a7313e29ae38eb7045278e60104911d602f721a6ec908c3ee58f1cb4a43da2db041c370ba698580a47d445702e0f1c31f2105870bc67da213d7b3711f83b9e35df7d1a05e47760dc6ba784a556c24eaa7f0363f1d7f16bc298eec0cb9407226be3ea66b6e51f7716933f66344bf5f8059f128360c35358a88bb9eb5b00b6360b80e9f4d817b3062f03e226eef14166c66a517419f712170ef39edc62dd6324c01410bc572f66002540b5af524d3f4d73e94f9955a1e00f19a757c72fc73564880f3751567cd64aa9693b84e444a775914c5f76e13a7bcc9e1a41a42965ea33122eb929b33d05bf5e31f905a60f5686476fb3caa0198c931ae533edaad65365b2db5a1c37c89ad8995445b8e897938b3d8250e3a00d4f05ea07b133901b449a33f72bacfd98b4f7b4b40618f55eb18ad39891c1a5ad4dee916d99e6099e21feace646d332a386788efa5a439861fdb79254e5de308482bd068caea0ebe6515f8c7f2df8d0bfe86a1d04fc955620900f3f23e2d881f9259b35975896d4f466ebbda40774f62185b8b6b485b8e5385d301d667f7f05f371f8797fb2a60870970147422ccc87dc2b110a444825a687e60de9fe7ffa2aaad2c5fc735b966622b698b56dd31d711c2c333f2ee5be772ab43176c15f363cc3aff772e18993e9c18bdd5badfae1b291c5ac0a698c316543ea3c53050b29c9adb03c917e1596764e40cf9d8b7e0677cd90f30397f8faed07c93fa3e6c891ac839c9afc2fb0f0615f86c8d558a24e76598a8dca9489fdf5033cd5f9e54504cc5fc169b344a1231417bc84cca73076bd833f6b9a214d920a84f6c139a10320d139c0e4268414755f8ab7f6cd6132e75a26ae9e653a37753f2a0676e7790a5a7ea3997a2400faf9495e888319578cdd35d651d9ebf46ecf06d3d96bba02163819010601715588b09b30bd7c7262098b7ae2c1a451d37bbe2a3fe5b831dc3e499518fb667a5adc3b3ce7a29e26659a73cc452d56a2a8991dd785d0ee6715a39e4555d4de64d509f868bd984c3aecf5733d721fe263781b931ef92dac466d88569f334cff212b35f12cc7ba05350d621fe49efaf08fbfba3a4296f1d10e4ccbc2bf74c81a1dac9376ffed726a77fe41642a6641ffd60a662e47598fbc921e3d88049b4879a2518ea541f0f018ef9b29bb8413de933c3ab6eccbb650363b8330fbb3c2db001d538614e4b51f5f625b8429143e89489cd9da62c1b9dea82aa776ff84cbcfbb12db550d991c9dfee57391f09327e55e17e75fd076aa1af68ca985607b7f9b4a8df431482d3ecf95070c836dd975a3dd7d0aaf6f2ebb85478526c70e79c13c57db5f8b8e945dc19305df00b4a02d3778cea416a15a459768ad77ae2c37e39daa4da1b9e969ba12e41256ba359290ef932c6113b8187973ee69aa2eed7e183acb101352b9c9c731e433158fb70f4e3e9f47fc34eda9bb757f8eab775241b2d3ff80cf5bafc846eaf7aeda7a300bc5d64889757ed7e8e017eab60f666af330fb2b425b59566355eaca7615b6e574e0c58a477e91f5093c1208ae6ccbdeebe7fc0bed0068be9837606d2f5e28313f636a8101ed1574cc875f0381d1d651f2cdda11b53a47313cefd3d688941b71891d3a0512c4cfe9533768cbcdd19c5f77ccb9bce6b1ae1d5c6afbf5ae817717ee62fc39e5f268983930677d753bfe44f01c7236200a12e8c37fc10a10b6d40783a75048650f64e025c0022999689d130e9c7860e3be3a19a0f0a09e78ff55af05b3015cf5e406aab91446515b7381e4353c6648bf69bb16dbc231f993bc3d6229a03b55d46040ef9b1ee0af6bd4cbdf032f89ee5cb92c3c0d1a6c6d559a3b6539dc074fa6c4eeb3e75704c3a416f58389fdd95445f9aa84f192d14fbe737e1ab562a9f1464ceb3dc28153700d6993b2a00f842a3571a2b6fa3674ca409bc6d8c51ef4f0630fb664af01acb664f8a137b7abb48c78c5debaa010f9c0666f5d040f2a2a269961a4a8ead9cfbc938e25bea3ab1ebf5d47aff7a79232e43d1967ef842cc87451893b070b3ee10bf409ca14dad469b33e9d592bae9b62aa7e9827dd0ae6f86f0a1f13b4b7e3569980f5f0efada2a439fdbedf68c1d5af703067e321d19d39222808776ada92680b16fa636e9dff06c2f8b2ab5bf2188b0b08c741abd062441f11a349e4f19d23012626cf740ade1d85592c2f2ef3d1871379cef5e7c49451299774a2806e6cbefe0104d73ed4580ff51e5a4f36c5bbb3e1ab5c6724d1f73f9e02e6d6f5a5a02553468809ce7e20c4a99dadc423356e857ba4edeb5639335e400be58b3ec3ae30b29844413d889ad49446b594ca9968af287e595bb0e35de3986cbacb7da59770b83f1a749576f8eed81f22560d65a2f30d899a4fd92a3c95653fc38928ca94e87c3061ff7f5e84f407df18a512c6b45fd6e66af5646df942ad3de2304a6f5a3d85315c16e2c79a730f96bdafb8f821f26bba3d4f934c09b4ccf0065c338700bb9d254051d5ec8165b3d04c91d410faeaaf52404a12d9aebe6e753c86c25cf597b49dfc3253c2ceb28e04165e0e3486a794e3f0809025c61d051a6ba8db430acd140d6b69fdd5a50f91ee890569c939a5691dca155991be37b5de88e094aa97ef2b55ebba99321b54bac4da4778457a4f3de6a06fc38f5b729dc6b34d16b8d77bbbb3f2481bc905d294c3d15f870287b6d83c7f30a5a45f2de7a6f0d7ccfc1ed6b2fb30a4701f68be70d5118ff32141c5e2209c4870a182ce64a770164193a4affdf7365b8c99a9a9e0566ae2de760ab4423a35c1cb249b0608147b4a4960340e1dc7a87343651d8895a580c37ba52b0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h242def6ec0926c38f6165fb3ef8d2bb22aa7a7fc21aae2f9558e3b535dff2a5b057b96285c925c3737ac6bc74b46e7605243dec0227a3a56923355a556df29bdb61fc8731d65134f7cd09e16a73fcc56fdd1de04963e01bb09716a1431e74d000725eafd7ee78036cf844698e28ddfd4d14502635f09e8f8ac93f77d71f82a5aa9d95b22ad962d342ee6c1249cece8ed3828a9d794774c7c979787b9943faedc92f53966ff0d594a3df8807e44c21f63518797abacf0d24cb428105e32d2b9af563e19fe8f0f12b5694689e3e6c379be01e772e8cc34faac55615cc829c1562c485e3a68e038524d2e8df2be00eb2bd5ff5e73a5c713f913311074e50a2cb97c3af4e99b68f003cd94b43ae08aeae324aa0b80b71633d448d4c479a4f1cc892f2d9049c18c3038e5db2fde096d05c1a329f5543b4f911d98d7c368cfedf6c86fa8fcc1ba9c74b35becba480b35b9b1599eab7bec74f7faa6b1f308ef66dbe6515e0f0edad12fde9ae8920e869ac29de5cf090f31e2ae4dac635c55b95cc95f80cfb687d31326a4402f2209be524b87c0bc01c81db2313bf03d517d14af8496a6a4f1c820c1059bab430c7409ebf741e58b171aae3a6ced8933de1952535b11eb19e14d3d8c240c6a2787c68e6de9a28cd10ba0b514261eb86d824024c2361cea6c2c39cb8c1dfbd68d734d5b7697b1dd7fc7a793f2a94b56953bed25cbb0f75f9e42ba4f1b1ff520933808ba9cdf9bd1f76a241f9d8c58a57695935872dc52a054225bc3d8547c2f858078527899a7f74526248873f3f06b758515e7182fad95ff9384ba5630fec525b75c3579c00e2e4cb73faecc47e3472bd7b95aa365e412928625262f57fa617da03f4c6f32153f736d39b54086252b3033e715ee6518c670520cd62610243c8071d2dbfba8e78add48c0b7a2929376f25952375e51854b7bcdebb3538a67f14eaadeb962de562d531e21fdecf6f5dacd419a298f4b0b258917abcbeab7ba8823b92a54e82865c03e98a7bc2cbed88633dbbf7bad7e438d8052274083781eb104449417287453b0fe1b1458f51631e4785b110b9056f64a5dbffbf1e1357e19d7fa46570712c40c1ef1ec7f0fd41f27e57ad2f0f78416d43d577f44070c48f4fa97045cd52b7080d718d105bdb51121087772f3f4c1f724c0c12d51c66586ffe8ef3ff3097e3241fb27b32bd1b503a8baea789ffaea013438bfe2a4ef41348b5280854a75e1a1767833a1a48f89d36eff0305518aefa0eaa14a5ded0c43159c6d93dc0b6f023128b2ac723f545f6af2a858f476cd9a0f7ac2b213024c750ac5b608fe0d13ae7d0c48ff63953b091638f1420afa652a3a8b72c25d98771ee6867faee310dc92de3b5305683c826203ef1f5192c9f70659ec7349165b9cb1cb74ec843c6634950958f676c345fde2e7858f1656d2f32cce29f70bfef31c0727d86792673ffc1d4752d61ec1c32305b801942d54cd963bbe2cea31990f715ddd03bcdf409a949e0c435e688e285fe4fcc979e5a49e1a852636c71ba675a08490ffcc8b6c7626a9647389daba3f176d57c4d1befd5a386de9aed22257935b8b8ddec4aed8df65765a117cc90b3708b07d8b9713482a7f2b27e8736bdf4d498ce9c5a2f26b33a1683c92d474b44868640d350603245e39c5955e3a21d84f9ed78671712dc04ae204b33ee426f82b7acb3d692d1b37636cae1e44842589e07fd7b632151792c5351a34dea08e3330421cf99dd5b9716f5ead9aa039b5a9d0509120c35181ce79c82f4a35e2ee273cd1ce59793b99f17bf736902b3892cf29ba4ba771e5b8593638e39a5f1ab7cbebd4676840bdf790d5d7fb150f53de8812c93c7e8eaee3cc3502560b3fda5beb315bca8fd986573da464c251214c5795ec72adcdbb5bfb09abc5401fc0e7ccaad853d7c6b877b05cbcab8792c04c7d1425c40e37ec230d8acc46771bf871ab8ecdf16c52bd7eb1914343aba9075f1d67829a681b99a017208a29a1038a604064d80728fab988b24afc145ea6fd1edbc73b0862269562d84b7dcd4a63438bd471f52b3713216fac827aeb37c91493ee22024646487b4261cd4b9e8fc624a94f4b5132f1d2598550c5e624896ccffcf05611c450acf612f928ee8ec0937b171b4f71b531a60cec72a87933f266cd8ec6a7b2817a11eadffe0e92dcfe46b8bb6042485c60baa37f2589a7e03bb591d85757a141044107f5b513e03b0e6e464ae8486a7ab8bf4d5bd663aaa0f388af3763ac755dc7f0ff5e8ae39ecb77364e845a10f59ab2bef4ddfa6a043abda99f0bc403429d0c35ce5b9a5530733ddeea13c22a8acf8cc128bccf0dd4cba05a532aa541e8dced9ff4f8ddf27ae9e2a852fe066771c858a756bf1b8b36271b50ec6bf4871c174359db798b49748aefbf9fd315561ddbd4faee1bd2bb82fcaea6c37f1e664bdb40a0e9c494007d73d3c1ec7729e01ab7105a836ebab93feb91a31618338dbe89579e0e0389558edaf3b4e215440b7fd257122d1ca5796bfc449499a44ec1fe18fe3f164dbb2bb45bcd68d0b149cabc00ae76cf1e19350d92dacbd3bca8ef99ee5221cd625fe1eb9b6a28d19a083e0c37dd0f3cce7638130daae6cc2f9729ee16ec2afd41eeed6a4de8484273a18b3e73443d692977e704184a27f2355aefac24bb031343af27fdce81ef1fa05855b535bd829bccf9789a10cfd0e2f152d6f61c61204ef69c3ce95aaa2318c690fa0ab340be88aa3f20e323fe309a6afc4c4fdb86e9beb3a010801106240e72292a1b69f339cd970230e94421f9dc2e27944312a20dda50e8e82e2fb9ec1109e6b69b09f5ad7690aa965973ad222cb03aa517358c031314fece66991a70442320d90e9fda8a2efa48fd5b003b812f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5acb3c8e77dd648bc506af184f719a28abd3ccbac13b123a82db4ac6017f6bd06e24de3f958728cfbc380fed2e577611b4b8fba23995dd6392998e167028a11d0164b0bcb5f2ca17dace86cc35b20d86b2637576b1415160fcd07c64df15151d4615e79838c5b1df7809bc13d57bd4804413a345959c65ba191e2af36416b16d826e55f174d39c6295714d3b25dd3d1d27564b02ca382204906638fbde739f0e0a928f73d8a17c071e20f74c63ca2d59a97fbcba90819cb28b69281fb2977be442671ebea37eef2f24e4e49613c8e7f12ee7fd7253cafbdecaaf1b7bc97054baa98958a267cef04ab0d9c40fc5f5882f9d3292aca7891b0a62e29e1e4a159d95e93e18616f23e137abb35ae72d0e9286a9d30d1d375e9bd4103e1af44c76653e492e66569298c5960d0d6e56587321ebcf5fbea7be39d0270ce7ee0b9dcd038a4acabd98d65c4d2f3d615aac052eb3ef38eab2abe03f2225bd898d9ecfcf1813f6f76217d0026b3f72e2cd039ef734ae52d9fd0c06b30a0618337a7f60d512c10e81060eeea31a2be9eb1a2e427c49bb9e72b4887a220e3d7cf91ce0f688544a37b313f2c741c7372f0ad9e41d102c4f62996084278655a73c25bae688cd6021d4975e936d82056d7773e537b7dda4a0b1b82042ca9af9f146c5d49c350d9d1391e145c8ee3fdc409fda349e5dd2262b37bad5211f08a5b28ebe21ff4fbfc7f6aacc6cee8d3a638021978e9f6069ceb8133f42a1e6cf173c56f9a1cacbdf2f6aad0d2d844cec4d5b979a7c86a6f6981176ddaffd5f1aff239c87bbd905902b3a13f83aff3a6b7c130531e37acf7539d47609330764ee21ee85ac014571486fdd6a8c6d1a393a8ec548a57b9257dfd3ea552106b86a31fd893a671a9b1d2211582b15be47d0b550fef3d99e6396d86b106676ab668afc5f7e8f8d5071d9e8740ff53ed8d569e3c170be442cbc9726cc60d07bff0f0c790739e0ee8da91a41e3f374518f2e6639b1e548880ef7f897ea24d8ccb48336393b405feb91e5f9193cac1c6b1fe781f148b952fbbba893097c595494ad1721e301155f365c75bd2d4e8af734b5ebce642a5a13b595a9327c19c7e9f1eaad9579c4b1a7f7c748afa84284dd66acea3b16c1fc66cef7f04a31d0780ce34756430216e0ae8af53e924423a585a44992eac728a5f82d0152d475a54dfe2577af059dcf68c5f19d616a78530c0af358b7f96db02833e598c3733097c658c0bab9b9f1b7bcfb612ca688d7aafe30720598a63a6259fd8c8ff2305b3f2ec0d8217376a3021cda3eebb120ddb002440470115f26acbfc53340d484f5b254886918ae20a1a03410cad2b2602e698df6d2c83a118bb09956b4f902f4a179caa02ba70df2a6127f04358b0c51b92fb4f78dc3a3c08c6a95b4547d1e347491afe4e052c26473457314373f031ff4e43108a1da6fb1ab65013a056ec23d1bc06f17b4cc33a46857cf96c7a276addc9ba5d8fc24a9f2716ae50c333b5705aa9d6ba0d77c0b984eb1a96e5260e18e6468fb7b9be5c72daba6252069ddc1517d5d173af9575441a37720fcbe5bc7a8d71cf830badca799a47a17911d9316051576a02765370bf9e2c60d8da3507c32d8c18c24f4eb2a604cfe948d7bd9784c77c514d060faf5b91732703c3ecdc0e4481394f5dfc677a273d1aba0c93a3a9f704dbb9d0b18ed835524a07a5bf826d96774d826ad52a3a2ac65417513ed1105bdd0576cd1615074a1238d10df49e7b1bdb72033d777e9cd22478bac6c3d0fb800e4cc8142007b62d2646d0e54936cd25e68bea88bb3049a5e88426911da1e24807f4216c79e6d3e6aba0746e7c9b17590a12ee80c98c4328c3ced70cd143230645a17a6d843ffc278a1a7cb5a18e467762ee13d0157a1f51d8a8b6aa4eda9b96f96a0be9c9db2a1a46dc0c2dd0834aadf621684f792cc5ceca543b4ce5f4d973b40bca0423492c8281aad2804e57e647641563db9e31e0832bf704734a3375e2ae7802efe9ce72806bd1677f0d5dae1632d5762d5f99358a5e7fb3540a8f37cd2c4d5501f94758e3271651ea563b88a6bf35b522c44e2bce85779dd46aa0d3d87a7fe6e7b2959b20c1fc069dcb716271f7d4a81563e68bc960b3dd4aaec6ed462bd2caae3218235e4715c1baf694b35456926c207874a5e3818f71a9ef9c63934ca71bae63084f6d5f93291465df8a06ab6173fecff3ca937b678026cc99f610994e3dce9cc41f47a3b137b536c66f1d19ed360b0842d067a11932d68c3b21c9a4abcaa76c8a7a78d8658b64f20063dc4277eb4a5f6e7621d010cdce6a08ecb87a879cbf41c8aafc888f7a925b1f59c57026b9d37e4c761639e05d22448d790b5065630d73af71f4c89095431f2f22b0a8b43ea93e592d5afba09c2a73f2e4e6afd789df980ecce62b9669d13ead2ec9f14dacb249e31ed9eadc05081e806630b841eac3028b9ba97510af5e700ac8efecdb7a242a66e5c593bfcebfa4b547e4d18f9820deea20c6021ac1beaad122d07270f97e8246c319a25fd6ac507c0fe6e89ecc2c2d8cf228f99814632a57301f2634b3815db0edebe6508c0f53c155748a944eb171abcce0717a3504a30ca1c9be5bb0e95fefe0be211f0e6700ef444a298d7712e2d45e949579449035492509856cc5785ee2163863eb42ea60d291bcaa79b46b1067f1df59cc559e63ae44ff2ce36e36399a79086e03de6cc3b8328fc92cbd7b6f2cf17406fa90fbf56949b99b290e056008fb521896ee3f91f54ca0cc2d63bd1c8b9b613bc423d87413244f0bab4f1464bcb6f5e8f000afd37c9f5787a89a92ce5961c44b8a9854c64c86124641375eb3cbcac457e2ea34f9a4786d74e6b094eddf1343f4cb8e51dd0db1a402495;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hda711949e3484190e2936b48d8652cea9b4cd5e446a6896351fbf15a8d83367e5dabee9b986283f660ee90ab681718e792aa213bd779946ae4ac65fc89b8b9b090ece477544905c804e7bdd880ba902a5015e85387eced8c7dbde9207271196bd96ffa6713febae78ac4a769b33e18a71bd58b099fd5576dfee3c919490b17453705f6efc9dd538d7be77ea25f5458c337b5b610b8a0bdb215e3e0db3f681a496a22f6ce6172d758522c42076699f6e5dff043201b16f9279d27ead4fbd54e52c729331f5ff3dfbb77e360227476902dbfd90e9b85b90b82707b7539893b5d57cec5b882427727ab78ef22a44743e3277d337825b9738973ae71eacfbba588aef943c6620eb3e97a02ccf637908a785758a7b91dd32af9c4e638cfa0adf33b4c517acceaace2be3e0792c864ff317bbb1d2c8e5a1fb2eff8b5dafacb80c157a77606ef0abfb49115ced7adeef1aa4d2f6d6e8c4d53a35e4c543b23faaec52f92fca56f534f869fbbc0036a4b4f413bd0587d66fac2efd3fe891a1781c934edc2219bfb703e67011968bb2423edcc1b7ec9eea22fd3b7f3b005046886507688136eea8972d3fa367296d9046a7993f263d6037561b059e395c272ddaff2e71197522fc64575d56df248d29cce4642b3908b7ec02ede31599c63df2e4fdcc276490473fe6a0f15c33ff8f32db42fd57c63c68cec206453a84d830f21bf9dc85ede47c4278ee426dec7b24511c4ae87f7cdacd7f5be36374d697fc682f76eaa305c32d482b478f96aa09dccc7ce6a3042caa210fc5dbb3e2be575199671f98978aceab1a67620e8d142911a9586e3489b80dde6174c8eabc4a6c6f401ad74865c1abeb075cc50d57b29826b98eb7ca8ba299f1dcaf19831fc143485e2a5c4acb1fc282b0f9ba08bb7559e3a7db41f9f2faf9811e46ae69d3f11d3c3e55eb671e3758c454f3d7a74ba43ed0dd329312877cbfc539fa242c93a02466dc49121764ff6127fe4fa69f47998ffc5d48ca6dd0ec3aafaff9ff3f6f2e8617379bb339f000f70c94de9809209a74acf718f48d5c4f6a63192e7dcca9b475cb3067039efbbe348fd6de11188d33be823040031a5081f36b08f23cce8dcfe3760068bdc0d33121e09479d57e8aa8c48d43be4834e1c6e06d60058db23f32d6a8ecedf8f4d33257dc20b76aa2a0dbbfd3f64b3a2aef850f54810f6a83b89a5248092eb7e115ec9dac9c188089d1c9b65f7e303ea924caabb82fdf281b20c73578173555d18b2a15d3d153aec883d77913d0f8ba0e19fc526b219e271201abc1588ee143e2dda1237c98ae19d98365635d653a2b0ac0918173ce93cfcdcc34de03c8c72b9c907e0496dbc9605c9a8c3402bf4e2570d2154556ea5474f20f956a7570be3f7e8a45c9ae3c10b74bb761f4c4eafc2d2229ee3549d2a263349a128c570215281f589cfc36af4dfc0242f512f205bf1e99c2431d24d6271d5a57d9429d502f1910f7fe1aa8bcc1919b8bdcfdf399c93cdb1e1fe2739123b28f4c4e021035378533500c242a3b7cd3fd52d5cb0ba00a3f64709d9635b9f3de6a7cdd37ad1c0584abbd350e62b7c25f2b12e4ecc401d6e60f5b6d16cff87951eb4f3f8eaa960f6a7479e2d2f53e61eba901dafcf94c6f628811455d687fd188f7f3476f7aa6af292d9feabb65a3bb8192335e6e528428bd4b966c88fdd1193c994be3dd969893061e7de0f3d40c5c438087d80097ce6921a3cab8a0f6f5b9272c96e43b4687eeb09d8094e82f8aae244d250c56b3b20442f37a7cf765862dc8e59bc9d34e0d34fa8d9b3b603cc1b87440663be943d41abfa21adab5ba071ba782ed934f48740cf5588a38776bc204665dbd7ed91e0e5b529f591f44cccc26b9eb7e5e98cae9c84c611ace9029023b99124dc34dbe4a7f1758549b19605b8db06f9df1742bd5a74a11ec6c28824b2b08786ee2a969d825efb9f2b15a4762086a838c9e992b7856187e35ae869757fe7fe3366c8f3dac4252be4cf87b8631e9ccd0e372b566c61ad210ef06060ca6616b7444e60a6448e02c3855ba6b84806c3f491570da26b2ce7ff7427af0eaa668c832ab83e1b12bd022bbdf366a1c7fcc7d54820eff2e0234b5dbd1afefafe9487af3f3092bbcf0a40450bf19732a1bb00635b038d8dda516a462c13908b7befa9a4e40b4522f7578cd2b2aac8cb34edd225ac253b666f041f0cdf00e310cc7a2ae5d5f90749365ff46467791881417cb5b0bb6a6d92c58797bd536ff42fb3140f277c67324f4c8ef087e0ad4a388aa073f1a28d1f5612a72805b565f851aeb912e0106ea35d6ee6c4c108b7bcf89e6122a352b6a71f4ffdc2d136d1171b0f1250c74d263d2d2ce13fc405515e182a5c8ac8fe2ea055e60d1772b4f1d79debe102cbd753400ca7b55abcf93bf56a3887456486749b325db9e8df33345a276ae3cea9b645ca5610acecffd0449eaee8c52520a3b53e3d44e170f7bdeea1b4e87461837b35c4b4bdd822047ff1ba4898237e20e09d0e2dcaa1f2150d97539615089c568053c786405ebb61ca5f43b1e142f73e4e92c82a5bc1804b8993f54b1a97969b29c50cc2826f79578fa81dd851bacf77ec4b18b0f879f85c33ebb2dc57b0a843deb269c4a3ab4e863c57cb47af9a8b6a523a129b84705a9475482ab25c37e8e3691173d6372d90f93955f85da24b80e4955eb544eaaa147c1df5f642ab4d8566347e5a946d4eeccb7c27cd72f4419daa92f3cde4431064f199dbfc3a2234225cca9f0e44c774ec7a31001f488b1540caf299afad14318c2f562a6d2be7140e8a3a68de29d9149a6faf6cdc30af63471045472f167d17282f3840904e92987b56ea40a6d91baf0386d6b4e598c1b3454cf06bc555969528ebd3d97c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2f4c16259e8986435ac86b292200ed2b35e4a1d871fb2e6ed6eabd9b5803aa22c148ecb5867d5a9cca278cf57653c9e6e4e708a60aca0bf9bed960004cd576b03c62ac3f20b0a6d7e8f7a63f4c9be5958fe1ce9ced8d26180f780a8d0bd18d9d24d306228939cc0d35b3d451e05f64f7163fb636804f1e2109d700331c913df900fc70193d7c50654abc5198312dacf258a442cba6b0304b5c9fae50ef87a069b34c53acb25d6c4c366fbe6c1833b3b5c45a251cf5588f2252fbaa90ce199109afcb8226db4288def4de140259a42cd22ca66165b7f194e830c4df0b3db823d2d0e45b200c5c7a9c3058b7b476b9bd6c5593f1d1bec25cc1a66d3b76b761fd16bf688f74c18464c861b1cdd4d58b9f341c0a469dec01f57931f113c23a2f98c4c67a15d55e6a22526ae770ccbba76b9dff1f98e3902359c18cb06d057f255ac9a4aa4cd0fe85a4180e9cb4a7bb128a850e9e818a6a8de9d032516e5c2bf22ea59ac0abd0a80fa83ed9de2bf2f614921e50cfcdab2d60f9b0d570b2c8fa744c5135725db49237d73139934a27d268b6ea396caef60aaf3f3a53d968fcf8bc9ee05c298003625cea949d1e9ea8272279b769cc2b00532026a4b07c79f6442543cd5183b5b3c299db08b5a81c2cb01993021e35635691ccc6ad210f3631856fda4854e926e34e684b5864cf47dd68028f99e000c6f3c9fbfe4a5dd52da348b6eb0e38a8a46b92cd4d6c02ba069e697cdd0aa52329e0c8b0bfa9eb95db4cd93052d97651a07b74b7136708d7d49a2511d1f9960c05fca0de0e77d825691b0a2e7247b878857246f0928e7e2cde6907864aa27a745897abe6bf85b345816327a54326ce7e3972451b0406401ca29762cbde42af9ced8011bbf5899270d8fa42cf6edd1811e63dfcda75db8bddb743b9166a11a2bba2e502a30ec992800628beb4bfafce15c1f85b8fa8070b710ff9a03288d434aa8f1f575c5e7c69df961a726e22217c8ea0b0052039753040067f5f4d88109a4dad108ba8e2d39bdf4670b69d1a3ad946a1a3bbc56467a324d7019a497253673395481bde9e08d13576248729fccfdfcd923aec1da57dcb378024b0032e8d12c61557d593a781f37253480c4b86645132e90ae1745851b54b441196f82ca6e9e1b5ae7c13ae51a2ea22b9a685330e22cc61fa85d8396adf50715e7d8cbda685da7cb4c6eb26835e5508607c13969846d731780c7e9f66d9afb64d4f140f4edf26c558b74c7ef9ca43fab7417fdf14d9df0b8a5327a8ccf51aa65ea9c3bdfaba9b58aa4eb88bc697ad825b70565cefd4026dcfdc6183458e982bbc442c1172250fa98e77769687b60ce625af6202b5e320df043dc55ef06e51de3d61369f19743b908528ff546932eb6a14e8d041410b79d0cd2e1bb0b4219a9b3731b934f59d3d3ca29608d24650db8f58ca0624fa0e37681846734042998aa3fda46df7ac4abb786cc6b7017a68050ba9ecbb3e2f50fc838e1a4929c05e4ff27af65c23011899d4a0a77b0e6282d20764eb9e3fccae6d5ca48e595424594d50983f5878da72ed8b6a0458611d04cd06f782c8c35d2ba97c73277f45f7f78fcc9204e86c909732aa6c480d83153094c3c73fd817922891b9c9685ac4f3af6e3659e0d8906b9e74b55c8b92c7e13ba577d8942e9fdfcd8528da57a8e5d741b1ed7be63fae25d98d344d82e5820037a03a3de2c3a4f1c2c2d66d12e590e8e5f51f07dc6cf9dae06c6fdae7444f87cdf8404bef8969d2551091fc10009b7ef23fb4ecd62062c701b9191285c98f965a4444571ea6f38640d34d85880ebbe1d60749090797f88215911977a02dc013b7e58ecd5d90b855f6ec7aefe33a51f794e16865f5ee019bb5ce224e03262bd5a185357bdddc0f8278d3d1c5bf2664360133f883c7f2fdd0cc3db1f97d89899a90728b4290db419b421b084a9278a808ee7a17c6224fa3efb460d3ca93d032a7583e2c7311f9c201ba21e6e1cbb8f8f93c465fccee8002897dc6e818b5aec5d16cd6e61437f755f16ba61e96522a736a117d51674045967de06e00d3bd9ea019e986430ec402d7ef81a1bce9cb11b4ef223dd516df1fdbc8378b938dac16e3228de479183746868af3f366a0c324175e1a083911a22c0f9abdcfc264bbacd3be5e696dc5c9e5c5a1a8dfe23c3e613d7416efc19439d8ae63fa870347e33ac938976978c9888dd55c44415371f947ab00e152bdbbf39da137440a94f40f74e936b91527fdf4a2f92267f78bb744e37bee2c505c2769e8e4bbf498fb639b213056afb65d7def8a1d2123c750c69422731e099af2bafc65764bfd2d7ea208a2ad0e0c46576318ebb7815ee5288cd6274c76c8c258b996268f2dd95efc8fbfb40353f65685085d5134042c8a258f9e4ce380a97b2b606f8f4bef6d7b6da77a3e917327eea62008f50b30e7414987aaa61a6e8aad6620ebcf3361126be69bf1f20936653c5ab12bbd32c81e72f61ec0068741aeed16ab644bc83a2e9c297809a73f09f9cc2f1188ef2eba0b4609bd7c547edc721c094001757b94c680dcbf38f71833f994055578819bc09438074f1fdeaff03d7d63d070afe7aec32fff66a45eeaa07c152db22492cae043569ef54165a4bada23a4e8aa5f1aa550775eefb590399ee37c49e48f3d5bf97eec6ddd151ed76113f83be37649dec159dd327af268a7f60fadc6b676dfa2535d0402edd5253ee39acbb029213c917fe4bf2089ddbd5816668af9179c29da94377d421230cc5fc55c143e3179f5514902659246032376ba69d75fac959818bada9ad7039f7b443a45aeb7b41764205932d7d867900a2ac99d60ff1349bbed782f471301bb543a99548312bb3e2fc022a9ddb24d8da51a0c2ddea1d864636330;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha72eb4c4fed7e2c662536eb75b8596f9e0a84987a736aa60e06cc17181f8507a67b8d40dcbcae009b5442af7982c9112815beaf163a0d8325b32dccbf7e7d66c6ce49628691fef9db40d894db643d0e6b903ab6817f7ab2c56088e48e9ea704e1afda743cf65a6810f63a72b95a0436eb4ec0364172d57d88a00f230184b86ee2d4af12e7ecc3a98ea94c042d2e58d422d1b0a53d36445f5ff5d31b08208003ae26201c22a5f590a1f64fc5b83999139b62784359ab5f65c93e2128f36be4df6f7016a70ff70de84cb384c99dca97a4f7a50e42a05d383d17c43c429281926fea8474c3297a7ec189d30ead876570c234255e65a0e6627fbefde05ca3cb4c275ad3166c128d023d843fb0dbcd33d5e5d9cebce01ad23c01438125cd6e53bc556f88f7d29a26521861bc6a424dfd639e4030d6a86b01c3c9c31bf5cca2033934413f361cc0114b3d06d20bf9e6e9a96617a8f0a0b8abf229aa6fe14cd1006acd5728ce3dbd66765fbde325e3d9b5ec0cb3c047bed07f7016bdbe3c1ec8f628272dc3ad7c2a30f62ef08fa3d1b603abf3f7933c23ef9cc4490c226bbcb2342e34773f67793331dc9afb84ead2e49fe183168b27e4883905765797edfecd1efb6dd1f2913a90169ca6f877823782ae389ac5acdec33ab3abef80eaa76d7b0e1bdd95b14afaf036fb94c875f703c3af63aa2237470e21243ac8655d2bbafef562477cc21e6da4bf564cca25528a51f7552ef9fe68e586c2b3388a8b958c4e70fd1b6c9c1b5fde83c4e126fb5064d56298766f97459f3f3dd8494575bc3d3bb28c5d325eb836b17279f71b2eef8f000b8b572ccdf7df922678a9df4f88c0b06fca32a32ce9fbd47b02d2291746edafaf0a49b605233ecce95ab819c09d31684b846cf126e9610ce4bb62b614d1c03e3cea64ac265669a6f798452ea726f40c5227ddf434b1e33237367461edf90a2c626fed390ac7bc6aa0dcc4ef6b1186cde1ca4f4ddcff3460ead39f0f572532851ba7f8f52a28aa3f600b0951fbe698fa748d5736bc726949f3c34472466592403ba9fd7b23ff0f5a492238ebae2568fa1ebb4134578949d0893bd33384868b080ba747b323cd3bea9f592364dbc7c5ed64536f9c4354673c9fc4f76c48c0afbb6f331162d700141dd0dea6afd971e47b62cb26c8e9e8fa5ed3686f0c1c31ee6d7555386589b8714fbef66531d8d93f2d342e6207a81f9c1d5266ce86cfb1d2fb229bc1b6b59338ec1314411f1a0983e559cdc679f3f79ebfa9576de5ca578edbfb7151fa973ba04bc56dd1f528a08ed5e3d2f016c8ed345a9027587195332bf896eb948d90ca8b8028b1fe1d8ed488ad640bc89622dd6dd56f3694b10a504a638eefe88b1aecde0eb63fbf6ca522ecd7ad294840e64bba26dbefdb8462e8974812f3923edc89920940806c61ca623c3dec92e33392d680f3dc42777a53b7fdb0b91c6d841ede97f0283f6f1bf664e7205d2cd59a8650e5438a8f68113c1e6bf6d014d0a8e6911e9f1f0dbc88994491a33a20d55715c13dee7da803b58baf7447b422ed3ddc4709e60836f62fe774ece9aab7bce82cd953c63e43625e2d2ab3c82a0a2860f9582955688c9014d0be4864a61decc377c989809a18546a26888d7bafa490c628ed7dbb9e5fd7b5fb24c20a0072884aac75eccd37ee30ccd545658d40612c14306c7505cb982822ec45022359d68c61b9f791517bdb208a413e3f39bfe0ff2b7ab11bd9e59d4ad2b6581ea4b9cc77bc717b1f6026c4c9a22467077ce0d4b7890303e1cfbc7ad2ad962340b7ff47a39fc8d7f393ad39e826f41c2d9240219441bb91d1c0009ae8ab0d1820b07fbde4914033fc103b60087b1ab2021f2fb856a3f836b46e51bee14ece096434184bd964de7bf341b79ba659686135b037c0c26f0abb4334a30d39449cb6e247879385b9c0b18714e76dce6e708295e9541f6abe7a09c82193abf4b05fbda0f5ee1ba43c0d6711651d47b88af0b254df76ce45a1448cb9ccc5be489c8385af52541df2cf71503ed1ef1261a39a75cb7c9552f0fc5ccd0dde86dea72925df22bb992a16b0bf0f75b1871d1e6eaba0e1c376d13fd466f6997e5d5c8fdde6c5fa871df55b6200e689c96471145b042032ecc6b9589adea203de691a1f2869a78a801725459c95b55f0aa9bc338bcb0b613f1bbc90da5cb13d7de3ee580d88e7fc38a2412662353389746970e98884e7e416a1ce684a9d9b892003728141403644e20500648ea8457704aba18be5d7709256fcfc0b74a4a3dfb5433fbceba0433521f7822dda8c413036513fb4d64bf2305881bcebb87b45a0f8b5566bc8fdc3cd9ef807cd1dbc24a461265f439d202a0bcae85e0c818df9209b02bf9cfd4f49f002a1d8f421dd1c81f3a2dcf539a2dde014ec430156e24c398818fa0ae2a0bd15e189df0cbf3cb6ef5afdb0e230b4ca60fb8dd9ad6001b3b25961ce98929885840bc3a20780ccfdee8d6130bdc20f5ff88e6c1970212d866cf400fb5f1fd3af703b5b9029143eb979ea64f3252451f5d80d02c756b10544d545d5ac32af74caa5715a6addf991cbb5b115e31aa47720b67d658ffdfe649488ae4e5b0b4ff9212757ebf8378e403aefde90cda5287fc970fb1223769116aa652d397e81e0c55b36d0da70a853039b9f490193babafcbf91fee3a402cf1de77a685b75324f205bb50bbfdbf781094289e17b4d82a957ef3a838252d3adc1475b48c766ec1d3f6ce5d8d72a59d36e72c2faa50bdc8453a90b01c02e374e2622417e2af62cab3f62cbc429cac94736559ecc10b1d3fdc5b3d41e6b86b81772c2bea31a0fc8e614b8827965aa9aee4523b1cb7cfbbd3b564a00f10a0aea7ed5846bc8ef22944c7b70d2b2a624596;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hba6ecf63902aa098c9cb4169c740f38101ae68876d978145ec3bc8a02d5edcde3259a188b83056b3318b96e649f2afdcf4bd627db087a39d501016dbdf6e0135cb88327622fb9fef3527e1a84fa4bf104898c3e55af3f057b61400b1cb780518e99cedf15134b1148aeef2165ac39ee101480b47316acc44c5867695ae16e48f3fe39290461923cc4e18cafc885ae3823260e2c8d3d1355394fc8a041c9ff786bc92dfd2dc420c744504a12db9e2e02c6bf9abcbe76378d0ecb459dc686e454b9eb526f8a545b6406e5fd9b3b4efcce8931292d4c406243d7ee76858fc0ef513e9bc09cdea2fdae2b55783566c1b707f4988d1973bf17f9cc85803dfda5412ffc88d5266edbcb109b7ee2e07cc98ed951f3f38ef594f266c466bbb077340a5a453c42a5f5086e8ea5c0da0face65477476037770a5c3e8f535664d4af5295325ebec80e8cc74ccf433e91c5291562d34bba51bc266f6da7a529fe2db57ee4834c478797061e118f044570f04bd1516fc75f2809d30021d9558054dc24d9b1c64cbb08932252ca33890c390397e3e1553593c909e751640bf047dbbab5f545559166f450775371d9107e031884ddff86234dd3017601eff3ecb2fa0741691eac604eb1994ccc37b2a9e8c00b096f45acac0599d720ea2450757d974febd27ab8d3d65862bb8ecac5cf306d94ece73fcbe087ff98975d57bf60765e35dfdf0bf988a5efbd21d79c7714bc6acdbe9835e9c62dcb7db8e6331e810b1c7ce3c0d6a2c738cf0826b9b26245a177d0860a06a1b2f9760ab7ea42d2a74ad5c4617966b32739d0904054d5353d05016f29b13e1270544799e852927fca735f43ae3f0a37a8ab1448106e9848711f5698b07794f4984533eafa1499cb2de624789e171352e8a5bfbf4a3378bb3664c601e6e819b71ccbe4ac8f327724f3a71e1b0771546cdabbf875e95fad51de8db7710292a7a32e6c83676b461c8caf1e745d247a05b55d2ef59141be1081f0534d1c242f519d5d59ab3873c2049fb8ac04143791519eae8ceb970419337b5249b868def9f27a5e55714e4c25127218df646d599f8df8bafff522765ce0ffd28b7efa01fc7f5d6e9becc32f8de71654e5e8fb0da71aed209280432f9f1f51f0bb651ba085218351fe3d866b6e01f9e508438d603975b28e1ba6b59c1c3a1bac06aaf1045474e913300ae3b5958c58904e2cb1dfa154ffd72633c1c95ee1290a7e147026ee0071a5136f8dd152eeccb7fef194ff25105395f0503da7722c8e13292de8fcf922b4cfd0c530276980905fe44e0d3066341a774d4d6d6e7c0c2573c269f1bfe16002c76df20f143f45b05a28a0c09777567f3b5219d3bf47afb574da0f40de7a77ad04f35368441ecb7ba215a33f77221941a8882f79b9365157d629f9ba0043f8225f41c512435908a068a4760c706a8ec6fbff0cadd835d3d74ff15c17714ef5211e7ab1a6c73ccf188d45f15dfe7ff8d4ab0a0222193efc86e229aed4c3ad3cb986caea10c161d68a50841e3a3b738b87835f7fdefc2bceeebb590626fce84cdfe0321f469dd3769a58ed199b28427d478346f5b3b189dfa07913e95d0e1285406b5de3bdc5950276779db730b715a71691d83906415a2975e0d4bc51e7d7a48b2d5595f005aa4da0f4c986478e0192d1c2eb7836bedc8fe2aaf7fb161321ec8505c389dd587eae4388b54eab526bd660140a8f2734f18742131924fde83cd5e7238acd2ff418ac7a238e8bd107be9300042b9194a3fa7fa4deaf15edf18a0159e4e5c1fe21010fc2ace7681a92082fc2d511e764e623db64b9037addb5ebb74617ae677b0e3f10f3d09bdce644cb5f27e1df0dd6fccd40d98cb962174cbadbc7f42124520f617534c7d694596563c8fe7ab0e01f20e8d51b0dd9b82237e5640902ea0b27b39175a0d32f0eb36ce20580e438ff7b5205b607bd36b1cd21cf3b1a9ce890c02632d55becf9657adbba18282790b84c10832667c55676adc3a1664d83af83b141c309ec4910de304fee71152b15f9ff7e2becb4814d21c4530a40f6d4354650f3cccc12ad7a221706fd0f44c2b2e39b5ecb2eaa1113cdf3391a9ce35cb0bac429fdfa7331dbad50e9164f29c15d4ecdd2ff86b8b8c8aa285156dce2a3c34102f51d6dae5ebe0d5b388d2fd680c990c630902d7a8e5842ac97fd68ee80b4bec32fdc00179b9efa30c51134596d45e4350907d644d758cad4af1405d885da3c5f0bf632cb025708e03b4310b0cb65880d31b09e3d1d129cd2fee7c099bf5e6c0b4a7fbc21221448b2e939fc3609bb93f44faa6b3aff80045e76db4c4c80031a6df77751508c76bc7f8abf4548a677db8c309e9485a7a2a91e00ce313e99238c890c1961691a75859c24cffc890f425d2d4565422597831131f12737ef480ad31cf935e4e10f5f1f45464bc160baa0f6d51e305c877ac2f38a257df73294f10c1ecea70011b745452071815fd7305d0cb89f040074c200b8e3e8ceb2c28a3c4bd0184d517a661fb1c6903315ab9315b997594586d38fa28b80e2794e2ca9d382c153b4deed7ca68f8afde24a97c3800009f02af3fa5904f40a0d7e655b18ded7abe57fd6694ce54c208acf1ee7dc89719a9f23a1210565b527ae0e5ccfbbb4c62a78e038cb4fe7a1619f4c44bb6ca48b9d383a288c7194ef587507f3c5030671ecaea88fbf8213672341ebd222aa87c775010e05f397cbe229e26d32acb3b6f353fb82336e0e793f9b3b09dec31fa3155647ef38272ef1d17b6af4fe84a55ba0d5b3a60defd704d7655c840d228c27b5f7c9bf06665738085b438fe46e3448cc4256dd48e2d330663d1bb0efb3d6d9512b5d39f1af3c54e59acb48a27f24deeeeecd6472cefa5f4a7efbb2f02c9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h632ff697ba4c5fb50f02b8a8b30475c1ba6c93079c18dd727741d27b3eadca609a63d39e18a7850f71ef80760f6b628610aa8dd3c78cc8eae34eb561ebf79d730300ec303b76e3e827b53b643c3c606ffbe8577fca45d93c2dd8dbdbbd1cb670a614ca57e5fb003dbe62d84ab5589eeff26a35e0735d43c15e2768df554b62009639c4a5100caa68adf612e7e6d5f2a42b586db3773b131cb015e7c6daae72b80c9c985fbfcf981ffea506c60e120a01599904fbb39d1bb0b2786657008fc6522676187d7d8d61dc28fcd88b46405b5cab3861de7add211ada9833fc4e5d8ac428cfd5f96d8c78a84728b35c67b9a0e29f3240b0650778097390ee1ebf5233fa67e934cfaaf4a1b6ad7ace8b79a20263211a40c143246a861da953f9d97fb2e15c2bf28c791f67f5bca7db7d4bb9127b8f767ffa236f890a388baff1c00eb2d4674e08fc649fdfd561fc7b7d347e5688e617d469ebcad2cf138ab383b6632243773205ae299b727c28257f0bd31ec52cdfc4a83a3dfe8a88a1312d0589ba0bc4d133eb8b64ac5e6b9d12c018c51b18c196ce4dd13beed73735c4fbea9c6807779409b5bfb40a6551ea5d178c36c3ac612dd5801042e286cf8c6d00fa1d5207d536339b7d3e7e1ae301eeadb8ffd0aaa6b4117dba1ea010ec8b1dc8ad945433b7b8aa6b25a7e0fe3e0b90eed238f3a7c8fbf539676a78737839648d29248c4e70f4002565220ecc7f36094fa7f1e86a8a2ad166173513f72bacf487b72fe35748d5eedcb9a00a843213cf3c2fe0273b286865a4d7160b9d43c76df5e9cce7970d83721a70f021bf4e808a8b42e227874dd48e520685d4099a479de8df4edf9c9673a8c735ed78c8b648754a9eb59244ea7e2f3bb6eef155c9d511e21ebabf991ed3a6f106fb53ba91632442ab42a2d05cafe4a785ec47e74f8b8af9d11f105d78e7c245097157f4e43652a5c7b4202df42a758eb72caf68d75da6fd0a6cdd8973183371531036ac23aca6b6be9abf2f4a5402c19ed3088b2d32cc470f91147c4b84d5c2e1568399dd0ba31dbcb3a4fccc20f011165f1f5fe2dd3493961e8d0a247f28860b46505705ef850d4ccca7164057083b80cabe250ae5a72d55ae2fa676cc44683014b97112721b9453a9d14b8fc3c31fa7b6afe6dfa12e908a2c102e6bd132d397d1741df024eee74aa3802892b8a22afd22652197b47589bd4db3fb2b330236c868c602c71f1f5e3dd79377bf15dc525f11c36b8fca92021531dcc6d80c1c163f06c19f04bed7078e927d0e5c7ce11466f513f6b253bbed6326e916268fba4ea8624658883a05e1dde008e8c9253aac43573311f88a643b3601f0ba82074757c92721c978f2fafdf81db33bdecb9fa6a034aef709b7e18b4f03e13ee8c1b681f7a99df47c1a3edfc93e9ba04c3d2b3817d38e8d41556708018c450ba4e3d6a77306a04f90f579538daef9c62ae7af6062af50c07f1bf4b1a5c5097ed4906a91f965c4ff1574d022b50fc6fefb53f35a1ada6340e8be5b89cddf933b4b61568d8992bfad7bd23b108f45c31cd8f073989a462b770ff73efb3ce1250edfd799de6320a3bd08732503599bcc47af5f8b4ce416e6e8feefa4c2144e8c9bcca0066d7511585507572e8f8ce6e8e09a778c6bbff9f624bfbb31ac74e5d91876995480ae6fec14584f13a8c313a0591e77fcae5a3738c8fb5dd4d048136602a222f5c284668e62e8bd9cbe631f1d4c3cd974d115fb3a4069c26041c85ad548df69c0229e0b6f2e9da6d25546fc7195e45ac8b30fa3b542d37e13a6579d4d31ba16da70586090426b3014e075538915d7304362bf63956eab4a22836a821147e39d78f43bfd008466b506e44a6b4413773b14a22a1fdd9baee44b0ebf94dcf0e68e774672ae785a37f9472a100e713b376f75db3790aff26c8f7661120227c4ab29d339642791e5eeb9783a6de9f240522114525c0ba0d3ef7240817724024213564efea876c851e146c7da5778ad1cdb10e77452d47246898075258984bf923788dbc0cc15e19e5f16828ff92ae9b6e84e445f68305a12d784acd3d80044cbd5b0f43de96521c3ab3c47b014f313678aaaf15b11f5528ce481e359ade1428cac13ec1a48342ed139eec06ba5db3f4d746995ebde943f5ac8a4fab3ba743de60e2abe1a05adbd88e6737c8036154da9ecea0d4cd4e013beaf45587ac9456eda625e628129820a09a17821d3c0ffc99f88ba7f959fd562eb529ccb04975c2f8e2ef4bfacbcfb3602727a21f89578ce77db38c3280844ce0626d28379de6389eb13161ce89e993fcd583e0d185e91c4a98ac1c37200c023dabfd2e307780c0f2fbf0bcd3d7d55f93541a3b0370ab0b8c9dff865a6df606abe920f524c8e10bab278d76a9d7fb3f663ab18fd456b51cf8b0e95ac2fe32e747eba251c2e27b0f3899ab61557e3a6807f5242fc950e97334344e0039fa2287e2063448df733ca6e8725aac9e39b5a1333a9e0f4ce93a0b6d4e0c76f780daa1eeffdf8da6a7b45bb0bcee00ab5b731adaa4135fab5bc50144812586208d185ce7090fce04d7b0c0276f5122454f44f3a372320f2ad84ef8a45e12c3d1f552a3f43f84e319b78560524882b5805a1921acaf98e61429cf01448398604facda522f0c64d3601c75b977c20be22d5c485e5f59b73e31e0c48cee483150c54ede90152d6ec15b4dc724b8e7e26d5e0b504a1521dad9295d4a32c4c48f3d1bc59002b2ae6fb31fadeec91875a37eb26beafe373e04177aea9040fc5d0ccf87a31bbafd8f75a3fe6ff21774fa800643ad8ba941aa65b698c748e5364647a69ade0bb6cfc38d65dff824816021ecd7d78149d8efba9fb48e2498b0ea7741a51ba94d8c32343603918b291eada61;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h926d474f1edd37d070d79eecfad1b0889394ce592a461ce6d529c6de0ad758f6488e8cb5bcc2781f6ff68dda18b4becab652dc940e4049a258786dd3e5e2f7ed2f25f5a2796c7f3b1bf48f241ef171f35a89b4d23221ce7bf1a3944348a61390611a759da76849ec7170484e74a1e29ad30f473bb0a40059ff8b65f5140480c9d7a10651e1608da6de8123115b378561704248e074c1551f5e586ef221c8fe8d56adfdc895b56304ac1649c6090538e2e889abffb7def93409dd269a44c0f76f69c932e8564a47ec806a053d0c4bf77d366596826d12452fc7eaa799ac811062494e39b394528ce15fe4a913ad305ef7145039a0776935d1735dbfc7279cd38dc1d376efec9737ded767e82e0498608078e2df998a3ae1acdd8aa15f6e582941e00eab616a204c905eed83e2ea6502b51f4dca4af7a6bdfae88ffbc4fadd427631a5e11f098728cf4bd745bb07d157ffada87c8a9ba4b32d6aae9f652f51c368ac1a1888f36edc9b702e0f97f3dad6513ea621b8175593571bf46e37c502fa6caeda0b7469ae11dd1114b4e28a439e85b8e092ebd912c5faa600a2f540a4af841396a21d25341d8a3e71f65da570bbbc96c0e788c0287b5744693bf58c19ed88aa9511165ff931ba298a8573df9cf48bf17edde56367900a2f9936fff00ebca385075f03870cbafd319c19c82db2507ae0cb5f1a80745f83bdc50755ae394e80d71a5a6612fc2a3f33a0dedf4113e11ebbcf76c0f957feacce6998c68db3b6e2c8aafad8eef7787b3a873baf474181fd99e5054783138b9f902a22e8b95a6205db7f637d6b2279ae9b43c0f1acbe5d660a1afcc6a91daa04fe52027bc32a9c52628d20fc65035cba179cf507c13ac496dece17b0e626e27dbf61bca454da95273671143ffbe33bce60c493e5bce417027b17e4f1b2a1fd29f9dd1424b831ded3192da883b1d927c893d41f56415bf3ab2f528f1e688cbf1cb357ea259253b9309c8c31caa4cab2233fe5d22573f8cd63d20d114f7c74b138070cdfeaa41ea0a68c888ae71c3c6214363250f963752308912ae5878c90e305d8d2d9d19784a435146a7558be7e5b880c3e2ae1dfbde3a86c2df42f7169316e9c07eb598a47248ce2403689965a81526ca9700b8cdb3def8ad9811c6305d42c946c352476558af0497ff180ad2392a12d07ef77fec388146eb1579dc1371a06b348b686cd10727c1d116ae10bad5a8b7adb20ae9e946170d26861e4a0be9569ead7f26ca6a1353abf52f20f92cf6517ab6892602cfcc15aa41aa763038b52320ee2361627d861676d6f33273525ed5ac001c8bfe84aa1394cb2dc15212c4fd6d0061c70ceb0891f8e990a157a02aebda94be18352e0e777bb6498eca132720e5bb5de8b21aa1843795320d384114f765b035ed985f2a6ecbbb2c6e6fb375af6e044d7da0f81f50f5cb345560c23f03021814dcc8facbac0dcca55348c74b602e6a0727f5d32eb829be9939d034712cd8b6d90916d24d2ba3352bdc5aacd4e3515eda7873b2822741828cb1391436e598a96f4cb89356d79fc097465cd68c28a5929460d3ba5686ab5ad6bbeb2b6e2ae864c58bb301d65cac320bcad6e11b92b2f9689e22583545baad7fba863d6dd036226d2d416714de95259988d8b2011112aa0e5adb806c55b21f8855855d06aa036c309a050e6a545fd291fdd5877f515d4d03a0a6ba3a5f9591c2995ffffd8894a26a72352127b6d14400c597d0958fac1d2a969d1c50d1471ea6047d43e39bdf8b2955d334f30ce06991a5bcbbef9f7b65f1fe66aeedea1d716743a27b79291c8a9395038827ed5cbf7e6de9a890bed5e631b3a324628c90712c2706af989be9fcdb45f7088f591655d81381cd808ccda73446e64ef68d67701593e499d15e96ced06b0b7ec0fe8db63e1720258d76f305d6ff6e10915657e82b52ba943fbec3eb6aad3cc50350e9c405ce64bde0bcf706ca09d38daa66531dcc49494fde2f6d9c3af413be0ca1dd18427e122a1a84f3b42f134b08886491695d7418f81cec94028d18c5891f80aa4ef83b6b7ae2022fc7a3b45704c158b4046e960849eac3c4e3af8c995f1f726402e396645bbb94b4b947ca30fe6153bc2d3c0405e02f6641d4e0a77e7c405a5380f5fe146fdd5a6da71bf736f13899330f17837d35fcc494febc4ca2e70d8933403335f58f12153d46581969cd19b39c173d92ae47cef30c1d8cc700076d202237eb7d209b26667edb159c2311886c11c9597ad6ea4fd6a9669556af3030dcbd29837b848c1df39edb5034d170e63fe683b6c85e639b864808e927376169d2e26549309b150cc20204d48b86b26015824c3289e60cdf039742c85e3f2c8854574809a0f83df74c164d252d3fec7dcc144b04cc9f4c8de6efa85b6b3297678bce58657e5a75b3d3b0aed15972320d6dadb1aedbbceebf9201945a35fce8fe73828bf2f9fdaec8ec603921f4fcca930f0688788aa10ba5eb080196e985fdf832771e2e49fedd5bf15874403dce826effbdfc5ae9408610570159d96bf845c94154dc9133261718930307a086efa8d914315a8025cc89b7e02a865471c06281e77635e6102373f8e7e21b808397244ff30f858cf379dd1dc0e9aa262a154de3928fc38f7377ceec38323ccf14a0680242d7a365c98c83c563e81b6a04721ec423c8c58fedf5f4c3a854ba0ea2fb5f5e8651a237bb7a192136a3bd3b688e869391cb47682c068a325ec6ca932c7e43e2dea4756534da47dfe30ca3e6a6f28fda19facb48fd5b037d29d88e46cdf681e1f5c13f454ea14dfda79fa4d9a35f01a5cf19976cba15f70734c4d08a68cd88355a66a074051bdc834c6d62d19f9dd2cdc8651464fa9edd58e96f68f7e8e2a0462;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h155d80c2fbb774ce2858bbe7a13d9b437529e57bb3f563d877df12b80d5d93e13595ac8e978afac3af486478d5886e6d185ec94cc88f4a3e5ce3444bb3d80c657b46c7608ad766107d46a8f921060ffc5cc68cecebf74a9953d349421087edec79b8b362b8105cf1f167629afe43f4a5e9d64a43ee6bfdb2b06291427c5d9a028c2b50f4a47fafe99d460898b649b2f4c428457a77494483832504e5a258c8ee207a5beb8e86b4cc069c6f0ea8b2c2880d0c9543540093f19a1bff73a9a026ce1ea03bc24f2dee29f264244d9730aee6c7830bc17b700ee2b0502748caeecf1b6079fd65095bec6ecd2893d746519744c3aedbb40fb6834fc4ace2022306b411aff6cc1baa44473455fe70b62e57a5e7f7bb6791260d10a8451807df4687f155a03630c11b064327f73d137c37dae69e0c0fa85cb9f3aaa1bd9ff3fc7a1964fd141a882eda3c66abd683b885675217a05cfdb50151d9a92dcea31ff8925a155407c214e2ee3c90b2bcd1326624a6121f3ed3d95e710f8993e4b5514921dc95a10ca27aa4163a4b67f5a2ac6cf3969b4ac563717011e700a641a4f71de2222065066c7c6f57d1931e216e1cc883cec50b57eb8cf53a0f89f4ff2efcf6dab51e4d9c5f10cee1ead0620d24aeefda1125463ee141a5af975ab525af8dc7c1883d743937b7109787b14007655df89e54a41fe8deeb4f1df877c7f0a2dddf1d64d3aa157aaad46eb0e105dfb04d1c71af54243dda6422082c5d1a66f5306538e935d2f182823f2e93034497f18bba6b6e7206ce1d3df60be1b910fc39a22e45eedd89bc366f5298bc78043474a9545e4a94066899c57b1020334ac6b50c95048e4c26d1093dfae6ccdbe01d441f3cd40c40381e70def8d0ad6291688ab6e41efcc1b07574faf047d482faaa026e001044dce4899e04a3da926740831f44a1208730966dfdef780177543b4d091c3a4d445e60c54900f21128b470739a7f17a185cbc92ee5dcce4f57c88e9d2edcf3a5b57e3282ebdb94cf748e990d64110836eb88fadf74ddf57d2fdc31a006daf938fe95b58bac239a3cd64f54bc3a2dae19f93e915190a5e092a1c14a9ff457ba448daf8572347199500611ee4d64b2784671dd2d904422a25bb9991e56a8aa6b69735989fcc54c37bfe326e25c86b45576918e0aa8e51318242490a36dcf66711b4e87b33893bb2531e4f1342c5c145971028e1fd111ee354172763a2a4299fc53201d681b2a77b447068b81cf12cfde3fcdf25107bd7629a5a0438390112bc195027369659fb5cabf667c3c4a4ea3051dd3d9cb99ea899e89b27e3a9fd1fd6f3b92fad8a0e56af103f5b5085f9dfe053e64b1611e725e25275dbcdefded3b57a007ae0d6c9b60d1d269f28cc351f977122ed9169c43e92c500099da82d30a9901b051bc24f44acba7b4fb433ddcd423d75b8113bf5e48d7d1cc5cd8aad3c31d7a901a39033a271eeab35a660db9bf10f82932808cf236f61bed7ee87099bf17028817895c71d60eb7acb6d73e049d0e57ab46d26ce74d52136915b63e3d12849c16658f660ffda11ed6e204db565addcbdb13924e07e44af23e35a77d263d28616a9b5d0e39cdce3078acfd5f4ce86f449cf0ecd14bfe48fb3f958da39e6dac11d1af380aa5826b8cd503779663d327db83ff5172bf6c45e6c7a9d33fff50755c5f6e7d98db84ddf6d4fe9bf1759ca7181e16ffd713bd2d1262896a94ff47c45b386eb8217f905b7115eef8e70dcbc49fe9a390c0a32ab90c6ba034684456ac0718debbfe20ed966deea36724c6177530afdcf45f8e9b5c390ffa9f22542525a5fc277bd0fe515d0f61bea4c5e45b4aadc6958bd868b57761a561724b1d4fd689746aed0f0098c3567bbf7bd0ef5f4f180e4b3a1d9bae7203c2cca7d9e8100420b7ec7960817d7f4ff42535e6d5993e39357fa5a756cf2973214aaa3a427b86d4302302351e0f1266f3c6e9795bd6850025538423403e04a1479621faa71f19d722eb96e79e6cdaf162c4d515a632dea876f3cc0969119256600832de60091499908656f41dc58f8d2051714242d653c71d559b2a7a42d576f63c69c1bf97a61992d6059056fc05f886e6a18a8f538719ba6ed1bb76475aa4a971a30a60e35e6e2587dd22653154ebaeab5c4c59c284355347c924ac0adcae15151b5d0573159229de9ff8fa50c7e127376fc67bff670b199480083f91ec0fb10ccfd5c22c163f70df7a8b03ac35359d7d35466994c536b653b1f198ddc87fe521478b5731c5090fdedcf1ddbacb7ec8358b2617b1f8e00d05e1b9e7a119486440ae606db56b4e20a237290e426519b532f35cb9525b5d9bf7dcb9e80503c8ceb4a3ddb2f25b3513a7a7286952a7700dc0bb18a15c1d06a3a6cfc54c302b40ececfee40bceb95d9516d33fe0c6bd78af0b54113df4354c7b762d75727031dedc1007fb118ce66845fb80853f570edd2120436fa322c5309a5a0b91d48e00563cce8bbe533e94ee2ddcdcdbc85dc693212725a956c0b5a31e5939e61351594c11f2bbcd35516151938a527b19c75cbc9b8b8130f847dd3f04bd8274c5a64505d449c8c0802c3dec0abf77c17c2a56f82304af9b4812269ceebf28f97a8848f2afa8740a4adeaf97dd0ef08fcb900fd0e267999a810846e7464c2300e2ca25f7cd41399b25cfa4b08cf209479763236f13c3e913fed4b943765e2b22c9baebbd6b1f5238893a61f3014382a3e9cbfca27fdf6a1edb412dc16a80f617a23522cb2e0068afbc2b38e88ec53e42adba53caceb31a1798d6b4e4e1e7a5c947edda5e1b6708d6896558819faf019610e7c16b3fd5573efc3d607c7f4236d89a1337dc2ee03588b5b8bbbe6768a1654d67659dfcf38a0bd27a110d541a6b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4df5625c3ecbd0b61fb059b4021c5ffecc7fecbca1b9c76cda9f1098d30b730aa70fe400e58d95c6c16f555749388a13ed679b89b3736cbec37199d1e9c7ed602bff1f640c95ee5754bf71f57bc502fa6eb6e892076299ec449f520e44524f54f1da9cde59da9920672a50b2b23edafdab6e2a478c4b444dbbacbe203d8350025a67bc5207db0c193d78c6037059e6f57933c72a471834140b149cb0bf5792f011d4f4d98be7bd450233437a23cf4c41018062498abef82f410d23f46ebfbfeecbb79067e2bc7393d260fdf19ef112a2c8349e1f68d76d69c4812c183c616785044020147830626746da64cfc439dd12c430d9738a22bb8719fabae55fcb7740e29e7dac3d3a545d8c8d1b28bbb42d7c6f763935abfc8f0df8723775ef9e64aedef1831b81b1be4e4f0d5b5b41ee8c2d48ffac29d4ba70396ecdbc2b1950394cfe36d4b8f9e73c6a4f150e7b2834592749a3ab2212252cc31ce615f59d0185b48384b13bd995d63a6aa47d7e12ad0c062aab74837537f7da911c48328bba0c2c3cf5250e824ba031c50e9163eaba1327e7e46e99574e435555874553aa00db1cdadf17aac2ce5d29e6e2b74444acaa212b83ea4b5070f821248d77005f14d1eab1c52e9497e8d5a88777d485518681ab006b365a0db808df35ef3d5c5376dac35299805138cd14cb76d0f0ec4354e1dcee9ffe559a1b132b001b8290b71cae89ca13787158be2094f02a9d689357d72aad30842cbda46d2f5eb08fcfe390357efb124da45739ba64812c02f2d8f9d4d11c7bfb737e71b7f20b869f5c33a1d624d8a2fe94799b53f528bfa74cb34c601e1ffa63a476ba7536043cd9ce124b7a78b754bf620060db1283bddd92c3c5ed8105a5faccdc992d17632a242b12743e6700df00e1435a538a8e22e3ea27f8f5debd84c402b69e345e8e132f70a1cdf92c44dc865b44d026391e56be8500ac1cb40f02b5929b3a8e19c94542e5f165ffb9b022d4beccb0ccdd79abe3b00af46a062d192e7789e6c75554f707e691353179495d887e64d39759ca91cb892b4eedbdb07a158a6a92e644305ab9518f4a8a16d7aa24d9bf4a8846ba5ad1671395e178795db93bd27c340a62a03bc3a3b94ce8392dcb16d6ec9dbe97a145f1083a6bf0d12e8947801cfac62f366edb33f7124543df8cee146db7ffa77e5e0fa14a23add4e050f04eb92165992d8f94448aac43fb201effca0bbad322efa573f80f6277db1453ca84670d023c8b1b8417ec50f738c6661bf7f6eaa781acc8843e58a720c5ab421ec9ac76d6be5f00e2b0beccdfc856f13ffd774e65b55c8637dbd6c5291e913d43bc4be3f0977b7f935440e6d91c096625e13570b5449027607773257c23e4467bca4fb4457e10a3d2c248c2d5647614ce3fe52c7ab2423918db01a3cd990b99a9db1c1550becd65b131fdca4068435c6192b40f1e26f626627dcee6618175a202c3393935eb45c7e7b73996cc88a82332057f05c41107f245a317dfbc7f2bc7b45889bd0891c5252a28ae883da263710c23060ec47812e8d16c29de632bab031168543ca38b623f81e70a42d9bee229deed60d14b031eece110168eb2880b1abb3d45a1ebb3cca615b225ca03b6112b1a156649121a3332a3f9e716caf96f29d57092b2540b6e4d6e8867112d7ff4b12957fca8817e074f6ac157b99adafbef75eb850f6dc585100a24ef2718978098fb7e90118dc8bb1546ca0c25af37788a7a2353f9e1fdb3337e0510b1ed2e38d517657cad504febea39da0e9f89abb320ab5d7daa580067b34c8e628758c1a4fb1dbab06f93a285c66e771b3b4f36cdf80e53f1954589f22fa0bdd1861599debd08dde108c36f4e30e0f5b242560d2dc777914c7bd7585352e43d942a318ed2a359dcc52c2dc8a27c6ef42d902a08d3b17edf5fdda5bfb342da8fd7165eec2ee6a7603422750beb691f986b8fa6a0f3d05b25211fab20cd17d875293135d86f74a8084911e0ab74fb60459fd7e3fe05bf0fcdadf295f8c1770b7d58ee69690e9a03f39591f4b04e124b29e0d509c72660a44fb2db4b0ea7d32b7d1e8a35ac120acba499e8e09ea568fb2c7bfb08e82069f0621f132dc2d840ee3409d5cc98d749a30b8a6882d86d1d5d0f78879fee06464eae34ac95faeaae4ae94aa966441abd2bd5f978dfd212dba90d9c4b365913b084b4917eb3efdac32983c825d4c2eafdcf24e4ff5cadad11e5a0ed89532b23213edf8525d4a6aeace94c96594e997eaecb6bfc4822578e4bfbd814092488aefdffd1f82829eb1602167c89bd3f352d6cc1726a2be97c885ffee72e8034d213c7380fb9af7fbf52cd42a0f00ba4a367300c4360b9632cc65fabeb4cc71dd56e73fa75ceebff4ded19d65b49c94a1428f16d22bce6c611269451ed55f3827ee7b84098c11a68c97916feb03bba1c7fb7d7d2415319cd5eaf501d8b3fa0f406ef4ef065e1f07e81d731ad1763cf814e4427582e151d22f515039a2f03e76761a9268fb7e2b8c6b193a85d8c9c8ce06a6ceb9198791ff9bd52b66a362e8d1bc87faf995c51bb38cec11da4448db9a10e42a00703c53da2957ceecbcde3f59e3f5a6b53f27ad980ba1e6eea91f2b4d9911ae2237af6a5d3b401916ab972bfd24316b0bb950d3d6d717ee7c7dd9c507403b629dd87cd0f32e062b759d1486f9ad7402efbdbceda9f6edc3da6c69f6543dbb849e089c1b436d2fe32952f25eb50252f85d6c396de96a100b4b8d72a3431adc7a7b363d88dc809f8f53c367efd15fdc2d73db447ae164bee9ccf4e5aca8b592bb303e3dcf40aecb4bc20b60bf85f6f10bdcfd5219fa6e6544633523cba5e7e67e165a5a91f0fcfcd53b24349ed8864852991b8c15327749478c39f294a40;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'heecb467a15b25b5880109ffc3d9b26ec791ecce1823b65732e4c39a0873d3232eab2a27ac2b0ac81779363db8baaf8e6ecf9106442708474d87f524e5489a32046bbf20b4eaa250f5baeb22ffc9e06bcaa0ac527b5369bd3c3a754a4a3336c6a2265ba9a857b6d274e2051048ac7448013d3822cf1bfeb59687153f1024113235e515ee4a3d94128a1826e64b5fd5c6ae7e4e260bc306c090404f11086fef067491b66e574b5779ca7191f2851ac994db83b99c1ab0e1106f314d10daca20696de4e59bf3fe0e06aa52720abc52f4865faddcdba17aa80b9f57b866adf6b8851edb10479763055e76d995f986ddc766bb5e12b95bbd7eea1ac31063553fbf610473653a4f9f1678931fc50d84d7df2a8fe4c1a6ed6d8398f1696a568dd67ad299ceb3b91c62e3035576b49139afaaa0c8a8f49a53bd5eefc487d7cc3105549540a5fb9d6dec328479378fe96a1c8d27e2f79252d29373e4107b0d5d78094e8ca1f914a374eca0c2d00fbc46bb76372d66eec5e7709affd9f899a768786139408680c0bc180b0f585b97bb7edbef860c29f1867d872e789986d04ff83ae84fb8dabb246dbb75d8a738928b9e5f07986c2d10fedb5c7f51071b717c5bccf82ca2324fb1d6b0f922c3e812c5e618bc498c4272c5d0a4e31063a81b8311d66e49efbfb940e4cde8d5070e62a7c1a320e4da60eaac265ce5419d2a640a76c0fc78d176aaef05528fab54540ed0ea39feb7526651e18b48cef4ad2088cff7c7e11a00237d558cb6c21564d3dd72a24057064f89f7c7d40ac993abaef9ac98c8fbe53be952abb52c547f8583530d297a9aebe9c8396caaee11cb6ce491336550c7b70ecbb90d82b9be35d98fd38fa664e4a74085bead4fe95898f6cc1a7d9efc710388744b08f6ea7e3a588fc158f7c45484ee82e09f80ca24871e6b7a6dc02b5d09026d7f483b5fed243d41c1e132318162a8281d49271d671e95048316284f65021fb63bbe1a203c724515c891f85bfa0f7f515312a2dbb07590dd1a228dd20226418a05dbc7e6249a548ba07d45ceebbe207a01c42c4a0b0c415867f1a3cd5aeffd540068b7bb56faede21d5459db847bf5ae8b399f84a472996749807e25f959ea079303775f4139897c6153103183dcc555352cbc8748184331fc0c2d252f1b2c748ccb5248190f65397f42c1c26a680f86fb6806d36253bf7c88d25a150ec21c74ee56c52cde67140dd2f3da0174d1b0d686d1f7d6e39022ec06a1d5fb24f37a0455051c2aad325cfc92c8a90d9a950263243c41d08b33df5905707cc73262719ad77116cd52547df75707e49d2f71bbb14f97f616a37b99b13961d3c246f1e1045b0230c989a9b233fa9215960afbcaade05ab39fdda6f4930d11022c4fce39b51bb745949928ba170d8769a21e99735fdf3441c74f158ad4280da93d2e1d7fa3bc85a9678f92cbcc73508f3c970ef9779c2d8db90a0c1539d4655bf1cc515f12ebd7486419183f75a5eedbb56fa6ddfff8257666799d9f5af2533ecefad95988211d07283c63c890dcdac042fe1a105bbe28fd0f1ac40c0a3fea3665fd3a2339807ee7ce6e428ac2b25100f5f5c69fbc39303d2913e0871542b7bc05cd6a2d343eb84af92cb043ab0f90125d472c2b5f9f2eb9e4a454515a39e1087a7f9ecd7f419d201854573453371a53631f0a4c1c000379cd91dff3d0c7ece5487c78c9e8ca047b51c611c5fdba1595d1e35f01e3fabea0ba5c652feb66e8588950c2ed09ef421a19e11e931364b0d7048d50528387ca8f2b4b303b32c2b4d2a521df28934d283bcb2a7db08a2fa082f4fbdde6ca460fad2b59fde186b979bed6f5498818972619ba588fe79122e33ac2a342d3fb49cdcfa188414cb350201adec11236c3527cea246bc667fdbf1524767091c47fcc0d0926fc172809dde5e18001182ee57cc3247d9758f7a7a00121b923a2cb359764dcfd7816de30dba9a870d0dbe7a451e4e74244c6c661cbc12917abfa6f61b64d90cda04a9e2c2f8d16ec0891f9b8090d1b330de43c579bd13580f125283fa3d5e83531082d6de53c096c5870bcc89da441bd7735dfb61c3e4856d2c08453078eea037182d9de95ff1ba8412c5d5a3f1522b4915b76aee1ffa526fbc16e39605fa529cb45da000d4355486de99283a0211e7dde6ee15c21a684e5f309270b94433178ba4271e268be030d7ec7b31e3a9bb89e53d9cdc1793eeb8c49662469ab5624979bbeaa7500b6b3edcf93f45dcc81695dfa840756bde357e288732878cff1e82bf005308c77f8dc8f74b3e60a42e0643fa5342421f70ee8960e207bd83c9feabbf39f0181a011b71edcfc20204bfa0681ffb477d60fd7fe87b274c73b2828cc0a98d4d439c634a48659b7820b79ce5fa639b772750bf8f7b220e84461f02e5e945a3751a20485c3d47f5ef3a243611b35e329a386dd99a8a191b57b94228666c3483d817c20e5bde1eb7808628e800799a3dbf85c1e3bc2415b5b201ab3268a8456faf548873ea39af147df566ee5b89c42690009d342bf181cb4697ec67565c6d8ccd8620821dfbc8c16cea2386e467551e282307991f9bd5c257af5d8593d676fdacad5ee3d5233c4bf1b3c4e9879f9cae02df504fb1da1dadbd13d2ebed414ed308989e578e56de0f079ee3b6740e37549890d532d5f3f2f93620a8a779c6746e3e0a1b59d5801f3f0b0a807414aa21fe2cee25d3afc1a32534773906bd28f7fe19b6744fcf9298e55bea9ef27601a80c68edbcea8513dcb93e968eb8e9c7cbc7d19344cb89f006bdbf25e0452075f013738167684f813c95d5cb75b59885834733238e6a26fa0a067b1afcfd8a0a5883595eba18d97611a9fd61089d09de281557ebc6eeb75829423247;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h185cb2c9dea32235b930b6e616fffd4e6b6ac4dec14560515e18de1005c7ef38c76b6095fe7bed389b01d732cf73ba24a9b4d3d72f6eee0a937f04de4a9bbb9f5095091e95636dde8348ef40534c621e8a1645bb2a3be7b31e8de3be8d4fa0fb734d279e2fe58274b8b5a27b9b92fc5a1fdbb0faff7e31995bda01cc8db40879436419b635fe0e899605875212f840ef19aeefd4f6777728fe5cdb15372ef9a98a5ac99f45e9f5cc32b4c1ac1e27a75cfdcea2b2207a91a40c274ae8ece9ba27e67866f50050dc7a371673d88383c78db48641447b06d1a22e16ac62de41bb33044cf953a5703493a328de1828d41ff6e5718e5ec06a6aff927aedeb4a284659d7354332a9e5ad70b074f2dccb31c3d4daaafc39ffb3261f7f71c779a6468f89d5c8296bbf67786a494518a55a0b8426987ab7b77847ccf93ca393eafd45fe827f71099b51230bb857a1c5aeba2d81737dfaa32a815438143280fa113c5de18b3a28d737d3e78515e3dcd1f3f02a6f6e1d30b4a119106773094ab76af93e6c4031b99be9a5f18b6efa9d2c0bbcc31fbb835e44c40a7c447743d9ce0cd0dde5ef964c79120509585ad4517d29f339678c37d98116626466c632515cd8b0c7c33c4eafc1de79b8ba14456dd46096be262582a087153bf1b609a6ffef016281576b9d54651f6ecfed1ca2c25fa921d9cc0657c1518fe27e82ff3a6645d8f6588b3b1f5f3cb880493c774ad09d8128b69979ebe9b102575d1f3fbdeb2993f411b825966975fade4e64821f4e77869320a75507b8a2ced82eee0f91007997a862f5f87edda12310dcaf376f1b968d6d391be115ef3cd6cb31f4f59ac12d4b6b1c34e8311d3efab49868baf225b60da7f6e842faa0a3ef7a337fae16dea0cd2e06cf2d02430328245c19c18057347c4f8a0254530c392c9ff5fb95bad5f4f0df7fba2fd98d3915c337546fee98875ea3635db2391a4a0835b1cba8b321ae64073d7334261d72c890637b57251cc9ab8b077cafa99d6e931503838d98bd3193e8015f230edfa8201b15322871e6fae3dedb5162eebc550555ffe4ce91bf41c5456774461bbbc874023c871dc23ceb686536cef773e0554680de1175f7555dfd6b85b0430ddd7f00439f462fb4211802462de9eb3ccde0b6793a9dc7384d9b5933c8f9db0cf398e443a002aa553d5cdb0834e7e60ca17a931849c3a972f8911c88a5d5a1e5b6c21c7e0a9ebd43a51659893ad3a7f1e78ba742a0c9948d0b51c639b11e5012662fb23577e4fe1735ac5c1271783e642ff5fe31d82bb6e3c8a36e0e393f566007ed1240b6e39b2a3dd6d4517ce4200ef617737eebfe5c85414f81c4925b1f7d7f66157bf30fdac37d684c7135ae4162c47b8d35d88a1b8d58a3af97c13ccbfe6b4ec9d7ee8ddf3e8260bc0464313babb61d23bf9591e59089297e76a44c4dc3ef656f031b3f73925237072759610cdb32ec1b60a124be2f6e1e0755f712a67f6502d7aa758bfa2a356ca25ad89ebeb3300d03e82d9dad724459f47662aacdbeb3e15b19fcfad592d1a467aa68e0b2ce829baf64b3edd94dd42e20322751d9575b4ca1aac4c058a67ad4873f4fd7a64afe0559606570a69227177a6cffaf2faa1db2a8b32668f705845f9d429a2b54f00959b5cb8d94cd01624b109b12b48db0447cac96fb12eb27fbb049d021fe424e77a36fc353c854b7e6c079fa719252d31797f094484938753b86c156acd6fd783b492126d31d863d8cf55028adbdc22787a9c58edba4a41d32c0dadd5fd288d41e3109b35abd0ef0eff95695d4e212b2ef6968445c8ea1e208c2c4e2b65072d9f57b92e7861d0654f9b627628e200073996ae60690f29e4d824407fded5df20d4a3db486598e9e1546534f3e33cb905c2206f1c1b96e5830e907e7279e6939eadeaaddf5a0fd9881960ddb0fe739a0043c1bdc2f4d286bece96a14cd4c61fc27e296bfd47026147cb192de87743168f3ce509008ca14d528ae288d95ad93e1e6a6ce8928088407cd409fc651ccd15b3c82d7c8c5ffd5cacf39b3309b4efd386f39088dd3c10c3776f556cb5d687d650a36b1a70a63baffdeb9db8f8afbd5f3234bd7ba02796bae193dbf21a7ad141011d3fc680f67b6fe68b7ef362f5f399df1cac08ede796aceb77a61683834a7dcac5b9b0da0f498843339d9e251c2b29a11fcff5079851abad5e736f3dd02659d8802365662130f1c96444bbde9f43487708026e8bf3c4a49a10430e132f3f411910cd4917c2549be3af2b2914aeaee101bd17ac81a543913cdd2dd5ef3205f38bc354f1dd88433ec7e02b061a70d532d69c1a44974896dfbe7f3266befc92c64850089ef3c1dd92aa808226988f12f8a8cbbde828b59ce3f2ec2f52049907409a290a6ef4c18d99e4695c700b48bf4d5c7e8f372d3c1d2bd72a5db9a2f105cb0294d67149ae52c8c4de9a1950e763355b4dfcdf2b151d7cdfcff6944ebe78203a3529e275b8882255c18b1b8f0dd47c2cc1273d8c17a9384960d0e6e69be0aab9059573a7150437e9714d1456cdbfa62b1ea84a4a77e397bac94cd26aa3cadaef475d95f9c757699dcc7e351b7b448c0a571f656aaee883a7f2a8faf9b0fe5c9b161e4e0a78bdb333818e8fc3bb7b65ad44396ea95343e87041efcf1a270f9b60f316ccd3cf5b56ed2b91ae42f1b7e7df31b8a37969777b29872980eb13ff0dabc4a1d38f38680bb5f4809bff8a905f6c6ec4f5153360d2839b42e2d784427fcf27e480eec17720635b8fb113659ac2eeee8fcf52ab2c428eab4dcbb6daa8f0fc66f04f2af8700e4099c5c7d4fc9bff5d15c9172a60bdf22a928d5d4e72d8da044a11f4a2b3568bb8e9821cd69d8d34860cf3076c141a171b49d635b0d1f6146;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hcbd66ffa0f36254cd35b2fc2536683c61fda534680bdcd71084e9a643a0bb84ffc1e75f7ca670f8d9581a7b1fe81f3fc11392e2c5fcafc9a2033d14c12fe1bbf95cabeab7e1b1305b915e6845b9e93d8505bd01b5f7fabda80d8b7a78f4e2f5af0cb79f13fc389ca1fee35ece73ffb154faa9833f734d3960bf764c30832c329c5e6a9c7ba1294d51215f1ab82d9bff636a047ed5f7e6d17b09d2f6f6a57f9d429f0a48184097c76456cf0738cdfe0b5a7d9728858450acb74db3d79b03c2543de2dd56b94c248072c51c90bffd4fa4b7a0f74dda1369e05fa3cca1bf89b05c6a4dd73c4e8bc000991b289665b50b8b81cd133a170d5e9e2f7dfe08d7f78b869ba6a0d779f354220a5c0923beee7a0d295c2511036b0ae1e16992c162bad5c5caa0bbf7eef48afbac080ea836f72f03cb3b47090ccd8afb7aa2ca5d6621997b32986fc18aaba00be3a501d2bc83f17fc8f7bf76937a84c0f317b1004f5a890283193a27c8bedcc4fabab289ef2858ed27fd4f664d81e04cef25b891e75a26014fc9dd76d4b97a8348f4607bb51caba3a680c67c4012ee99786fb03e9bfc63095d07fe8138a74fb79517b4cf5a8a630624bab96530c5e8bd95691000dc2a441de0bb604000b7b9353ec554ac2b90139e51ed07cdc1f8e24522f2a1c3ffa99dbd71c70662d7f495c03d9a43e8949591bc957cdd0fed8e09c644ee9f56a11c8fe8e3b7a8b1bf9eb6f6f7b8be00a84062d41f0efc8073c84f8d08ea909ffe2173da4835b5eed06ae2559c65acc66ab14755553ce7927f2fb36692601bb8949aa63732a2e44dcbfd8ed39db21bb94b7bbd9bb1271e1af27d9a4ff35e170562ec5b99e95968f4ca48bb587c1322aabeeca95c2d862e8b76904878b4437660555a24ba75e468183acb3ce4d40647afc53939f55c7df722b0e88d61783b826b6a17c96be4fd171adcf82d4df4be3fb3e530933618cd6c9d0a259b581d1548b60327faf997ce6634926b14a49be28caa8e48abdc0983313f52af09934d725d9ee0ae32a9270996a652cc575ce80125132e5f47bdfc80233c87a7090204119110d82eba8172f0f6c00d7a7a4d0dbdc0fada14188880ced5ca77c535fb5cda8b43d14622a6d1a2976f60df082ba9862e6d022ed5eef5b6ce55c68f0a222b75401c7dec8305ca8af324071748a973ad69193e4eea1376f82ebd6c55f9f83271487603f36fc78a51cab919d09cd13a1f9573d277042979b375d61bae3c240995b279b04c0830c7c6b3ce6a053dadb76b9b8fa11c463aae2fcec81bc51bbfe2e80630e116cba8c81a4a88c106375c10257df39ab8b62c6d0b4ed7577ad006aee9bcdca081231c0c19c3a3236de7161f16f5d9944d916dbffa4541947487b6383a97933c6e31e4ba65f8a8de0865b5f034124dd5c321c18ecb9d3d26b9ef62e365fab19389b31ec960065e43ec0015d0c3440e32259d76b87cae7cad060d1175f4aad488d03b490bc87670000e7221a38fbc67609abbd0f1a7206d2f814c328edd9d201e2938630f354b286cfec629a1a9a373bd98bafc0d8d627f55a545466985d048aadfcd238fb843e474245067cdd819ffa2525e62facbc49188f06dc61458092c4a3bdf56a3f661072f7aeecc6f399f1ae0919921ae235b4b9d86f862093f65e8921ba95b71cb40c57262ce85e0d1101d5298f610f45f535beee1013f03d4b282f85fe3e50430e5feee1d9f08baf9bd60cb77d274de718e36e118426aeb957adcc3e7172278e24dff4d62aed5b4a78b420fd560c52103d250ed34fdee0140e7f124516cc6a1136bb0b6e89b01d369711c2febb5862ef1eba97d7d3bee5e514fc5ada24f8e1d03de8a1e66ad8f9960fc21a088b10e34bee0a13feaabcb76d584ceda8ae7b525f2b74bba363361df9be3f76485fde8ebe1c939098bb372557dcda7eda83675f6156fe50a8c99b2205a0ab6f1546002f5a8e60cf58854929472cf46a64317a5e1072b18ea66744fee38de9be6b92dced80829d9b5e5f117b66263ba3bb4d03228f962e92b5c693add9519d7de0fd81fca8e316223b8c2709955e06fe8968f9e9f6dbbbc438d2628ac090fbf622509dd94933de59914d05e7f144e3cff94669a2a409d9e73f7b4e69cf4e2b0919bf872f947d7e0bd8cc061663872b80d0f1233c5d6c48d76671168d3a272e4e22a6120466f2ef13f7eaac5f0f62f58b0eec0580fe7d1bae2bdd93f501c01c1b3516c97341813b64ce5af648c8757382a5c9e9fa78039513ffa14773e6568c6b322350a5b68e370416b282738bfcac676e1a31e43b31e2c9d8b52f8eba2be50a9960c03a1438ae27f66c325ecec409f7dbbd7d7e1814bb0b7fbd0a9172bc262cd622065c12f19a194f40b94f7ceb8768d7ddb0d2717f7c264ed095de0c444b7055b162d435fea66c455565769234e510199fd89d8518fe5d14a89bac795832c227251d7742f8d7f5f44d1bdde3a3f418df73ff606e739252ef8145b20880cb5f7eecff15ee7833d2cc59dc2bbf99031473370cb930b8259abcc6e207d8e1cd17dc6d8a419ba14866d6940ec9063632759500b9239dc8fa233476c8440646042fd128f615877b4b09bd4d5c5239c3e779242d7defbd64928b68204f2bc9937d863136432c1918ab3007f5348b7a77143ef5b709971d76d60863ed91230b59ccc0aa6008303332cf59df7b039dc47c75f7d2c9c73aaac2a15d2aaa17fa53e7941dd455600e7a892ff6a0c47ff83ac4d55168a8c0560c8939f6e8703e883dd4871c4540bcb1c2966fcd61d838e59b5df3129fc722e9bb0a899dbb96f5553e5507e18605406ba7c59eb87299e3a1681831b5837c3ee568a6094f8b60c893fb7dbff85aa1d167e2cee19e9414b826b3f91d2ec439e17c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3b2b507fc125fec01fa2e685ce7905badcd9518357f4c2e4f99578a4e7690d8eac0bfed1e67df53d9316e6431f790ecb3fce487920a064fd85d594ee414faf0e980ad125b143313686bfb2f39ac7caf93a9158a40355ee652189367fcacde97fddb697ef8f5610d2f69bd37021c67efdce00bc804d8323cb503b3fb9cad8502a7dcea6195eb8dd256b5efeba99501faf1605a3bb5718cc1640714d52dd684be137390d2abc396c3d2895f0aaafb5e60d01c10cefe307303803df3a9133515f53a6af95d90cb82403e44370a17a990d99c0bd301800cc567a69f78a7e71948274aef9f442799998654b2aab42583181de3f7b6e1aea67cada067a3af798e9adc121866f6805f1fb3e0b7c117cf64c5e0b9d9f364dfffca4934d6cc14363e2cc1c0c9c26c44117d050743ae25ef2f1380ed1da1b4ca9a6e7da4fcf07a08e1592d179af507d1e8595ee5a02408bcf40c194cc8cadbbe9c134a2f2264a06e7974319819da3e2fc792faa2b586c5833d14129844959f65deeacb82da0aa9f2a5d1210019506e7fd84a05dceaa1688d106f23c95dedcf79ee751ef6442b31eda033af3fb52c7b53cfa0294e247c9a8acb81d80697f22d72586e1abe9fabe2cea0436308239b932ad6207857c4b42219809d7d8c7131db71e8ba879973e4f8494fc2cfe1d69f9b69af0de325450bb7e6f32a16f62a4f71bd5d5b7e8aebc0b1a24d299bd2c8bddbed19d7f0da1651174cc60a6342a3f4cf44e8b4b6f263ed82368306283fbd2ea35a8688cf56d45ed74d21c8a4b896e11ec774781d9e8004f4938537578661a2545bfa625a42ad75088ff99426289c4ef161967762a9abf8bfeebf6684131f7b57a8d96557138c9f1ae0570f23a1b4f89e66208f4f17c5d6674afcab2c5517fa069ed007a677d78bba67d5b384ebcb335053f997f4c3f8d6ed558f82a440d875a4452547045d2810b6a70718d1195956274cdebd53ff0ed16b59ba3b3ddec802f49a856d480e8933b6f45d33fc285a293ce5991cf448f48a7a643e2fe238b8f10ad037c2a6b563d83d039ebdeff4be021e4f9be3dcd69a128dc11071b5b75b9b6f36a4ef477af7ece76bd09a72b71d29d12f94d90a54e51ce7363495a9892963d2519e2b61e62638b81b2b7c265731e2571e793169d018247f66773ae5a2852ac08639d331bb8174fbdf4319bda5ae3182d6b12bc45784f3691d6b7fe668038ac5ab2cf0374f6ce152cecdab4206191bbe62a3b3ee9357bfd411ccefd8e221c7b11af68d9a2d70bb2f6614b847329ad54d004d8fa6d90da4edda51977917f550a5e12e727ccd30a5d0e873ba2a7538a83f1f52aa31422762169492669b3a46b84c00c123559fb18c1b5ab7a1a91933fac9e0f145672c0bf11adc1dea103f74310096fdc07bd779be192dff53715e75a3548856f89194ff29ec0e23c603e382f7568f7e480ed3e4afda55b6183bf7b7e5dd16286ee27637a84cb6b2dfa16a0ffebcc212dcb5c0e211cbe0192f797f32a8f2eade4aca2d0eceb80822cedee47c45230ff35633cfc8152c2fa24797f520dd840e01beb77e0f774bb76b431a8a214221df6b5794092c59d3ae621f158af2deaf8efce0717b88272e451de2599bb8305b2528243fb802dd5f2c984b2fb5db8a86673912d7fcb25a9e3bafb05856bf62e2976d90912d182c940f965c4691aac5a2b26a1a850f3ec9af6af0e71e28834e66f2ce9bac4c9ad3c28cce45803db736985ae7d9eb57cb09cfd1624d33cfa7dd4217de87672f1993bc335a36dcfb94881557351df649d785be055f03dfc391adee687d86d4b82426198447905153f91eaaf1127959e27e4b461fc56c086fd33041cc976edc882ac1bfb8444432b8cfc1a0f970b7559f312cb02665e3b3760eb70dc4dc243f49d6c34df1faa9ab9c4b084a661cba9bf2166c46d1c62acc15a820b1fdca2efb5038cfbd74442f22bd0098627301e2a166828994cac939709ab14d003454fdc03d5b9be2e0c7f37b51db2f1ad09bc0b283b774553a568af40bf5178e6b9cab62690a265bfeaafc38f6ef7766bf8118865928af65111d78484c44e38d81c5bbb217091d42573e4d2fdd719d0ee3fc66cfe6eda78049b206691f054fed8e0792f1aaea76a52aa1b3f054d140ff0b0085fceded37d0389885973856e6bda1632b801aeeba55b3a63e69cc5d68a18a43b2b56f5ad4a830a534533e48eedd8fc5e26c11239d004731b04a45a56aa6f46a5d2f923e5de8be5038e9c139d99d88361c3c474a29fcd82cec941e304bc9f56ca53ec723ae6a778cbcf79d6383180c4e2ab1ff32926cc00e3124c93b8c1bfcbb628c64be0e7d75f4ca1c7627d22c274a47875999fe50edc81724325fd5485bb7a85a153f265ab80d52726981afc70bbdfb644bbe26c15d22e7dce7cac5d50f25eecf06ca358819d776034a2e17f82dc13551bfaa585bffcd38060f0fd1094a8f890ec03adeb6b4d7baa3889719372266435b3307fb3557a4840c03a708b269d9bc82efb07b9a6c602258ef2d691f2e1a929487cb914145f53d616f92c4d86708583a47f511dd74f79fce07161050f41a30148b20b4f5967a92be5d053e25e6a08210c53ecde539821c5d8fddb2b5e1da00caa2ce94a0daeedbcf1085ed163dff5f6c7201522706243d86651e2d7c200a7e6ffa24003928e9017e8105cd2e5188f812cbe16904a4b5f76d491530037434d07624e88276624b7fe93c20eac8e2554f192257052ad34785f79cc97fe4594447a4e8cb63e2a578d091698e5475ede34c9895245db3061ec463b4e9304df38c539003153f063a9005d389bda64ce198bf00f00957152def77addda7c34b134c8e66a515fec8965495c23e39f53d7f2e73b6a47a555388d0801cd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h71b4768d3f76e2c5889765b157e79150fd70e43f334dee2a4bdd0e4750eae1ca824429cd43d0104717c37e70d3b831f077492e914735ba401dbad7165ad254fbdf256a00f7514d42657409e6fb99f8156b5e78b2e60a97924891a1fdd7237045796a1b3849dd72c1925825d539894c2069b258e61bf27a13d5344027e21d3ef7510afd732e33690001ffd40a46354b784674b681742b9954f7ca31edebc6d063644d9d44f44b5719d6cb5224091fb0395ae9b2d90befc63298e219520d4add8363dc2aa50f8673df649a01f7cb75ffe2e85aada77f0d561d970ca1c0f5c6215d6d6ec399413a7ba6d5bd11aabed6a9c35bc58b2b5f0536e77aa861c3f99ba151b3d2561656ae90948b7415e9673ad3c2e23ec447796c68eda4488dd1c33450f261e9eae71686a964b3b259d2dacd0ca0e17119c985b4646288a8ed9f517b8c56ea47f5d1018a953e38369039fbd5f158807ce56fdfa4495735ddc340bf7a3d81b393110414ae290af19b03a10cb36443523c865842eb176f3afc01c1f42d4b6fe69a973853a46020f875dfacaa1c845c68b8f879f051a31dca7a5c771656c7fb01b6e75ceb6e69073c26e38df87f8286fa59946c05cf92c2088a633c7181dd91e780733945fe7c15a8283736ead2447cadc4a4b1d9ddc20cf3f2f08df93bbedb5aca5a1496ce4fd5fad633bdfb39fa82d441ff4798c31ff378d2d232e74c1e4f1aed2ff8ebfe163e48ca7d8a0064a9c8f3cd96405b0b3e9a1b2d00644e6abf1f911bc5c806d3ab96eb789b0a57ae2a92250c95d33e4c5bb960d96c8cf028054ee1fa977749b07792bf2aaf1e67fa0cd968e000fb54bd3a2b296e1fb25e3fc13b95d31f5c36e8e48d06e8cf9e2250adec98a757c77bf39091d7538c6aee7f9ad437312a5ecf9b1e0fe3b13d88b1ffe3a8c33fc2f286bd8cc4e14189a4534e3ae94f09fdb426aaf00be39e1e3d8f826249b9418e6110b369a67176c981a29564e469f6af60987c1d7da5b199c5bb00cbd6943c601b57ac200b62fabce8f6732d1bf788ee9e027662b0c5c5fd5f0ad36da8b8e13fbcbe6a16eeb707c5af97cf4a94347680068149d3e72d273efd58dfc8a07848ff638961e873f99f5c193b3d7097b2fc2e5e172b4bdad5921f0cccbd7a73a33772cd91c015de1948a6e23706613881fcf2e3324a1aa6255255cff635218c2f94308babee012eb04f24b48610b28e153148cdcf2c205bbd5d9e03a6623f8ccdb81c086230880470467c5872e0207117722793204f8bf372ec8f169e067d935dd5f1d7540ff81d2ec6b70a68275a7110516f35bbdb477743af2529de409e586b3abeccda64ded9d6985588ae16aa4ac871d3d208fd8c26419c2ab5ca846c5722d821e96b47697ceef3609579f57735288e4d194603b70fa4f28e5c588cbf976f4b278400931453cad95e6c8caa3534fa5328b1f6d901a17f9aca2d04b137f0d7a635d4ac81aa84480d94a03e993f36a325cd5ab785f66c777843f10a3defad1e2c1d0b2183def5f7fb5c92508b1d5cceafcaec043628c1232692f60acd09212800d03b8fb11903988dff7d51a120380280b21680ea2b107f6f5611edd9d2910d0f77d357283a8a83442e819d09cdfb7b65e92c16ad468823ea812d94877111fdc2c7e7562a62686058bf11482f90a698152e1a3c412d5e54f6d59f52f96bfc093ff5c5f62027d26eea2a364ced51e9af5fee4d1f2086c49aef0ad18e5592b33b742fafa01b3d4f8976ca69f25b2f20ec0ade6f346a9ab008c97df0828e399b48b3fe9e2414e5af31edc1e84d4507a557ea559d80949682997c3fa9feef4504537a41ed6b0043bf30e57e52a336daee7d953c29dd2af4e6aa94f4771a9a30868ca1c19fb0b11750d1f037213ab9c8f30ea85601498a248fefc07d207bf7d5679580a060e16758bda6e7ab2609c9a30fdcd76862f12d90ddc0c832eb46a54ecafa327df1ead26f12a9ce8612c8ae020038516bf45bc5531afeaf032f0bfb49d41a0789f67b518a2f32ba8e75df5339ac9b5ce800a67ce860f9deb903fd1cc1c7f94b6001f6c1b3ba74f580d8efc9df0501a2fa9a90babe6cf96d970f523103624362383bfe64360448f7c2651e9713dc5a333677c87e0fc0e29ad8d34656ce6069f6ec76b3f310279d668ed05d72525d5947125ea788ccaa4d1cc33e8ee13292b05b1e09193a7aadde1d0a2314d403ac6b46a65d3123f2d044a78032e7c8861f95954162565be2b2b6db6742e042e9f7796900de7879698af7e9b369bd9279375e72191a44b7b07f17bec61beb1f44c4410bc6e1bc7f2d0ee6686c86dd3adcbd7f3316b166caedff707625f9ecf05c790ae0097b230839e69dacae44d17edbd237408fa5519cdba35d5e12378bafbeb83844119acd7e3ff6d09a3801874f10d31f306eb7c165033b6f0180e8984746580a0efb94f4808f4cb119701c914ffe421622daf04a2c12045b1867aa7cf40b47f479630298fe458b78be833d9313bf9372f7571b1d428572ce08d574f67ce162a768e2d032f90458d109cd3e7ed6e2d2ecb8cf3ce830e98330b6b3af90aa0c0be101b40ef3b34f5036633d114ad86384728914ac79bb880cfcb37491f957a9ca2eb679c79c4026f5c95c3258a71cb21092a48eb0414cd1f0895cf0b881aad4844915e5c3e87471a86270469074cf07f7c3c5abab793a554020133a7eeb3e7dc136ac29d0492a218c9f633b919806a6da0008a2ab446901651b70a492bab2d2379aa7996298d2f8773f9a290ba3ad1cf73b80f0499829315960c87a238305e6c8f3713fbca22420db3132e268dd78aa818be3977379f09fc013127e51e9081b59382d08c1e9258acb8aee71695e534b484bc97cfc96f67d07ee3867a8cbf35a29;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h9ee4e73ff9edfef7c4eaffd27e7488139f68b98547b6160a33bac91fafb9e404ca2cdd693b3327ace6ca68d94b0ad68c1392fa1645b4e4221ab26a4b94bb361a5b958e81450aed9d061723f4d54f8797ca4c9805a422b2c3a073b85d4d6d467654b02519ebae681ec65399410c40a2c40658332ba799f5b58f0c8c2d0ba7ad127cfbec12ccca439790c3339a61a84e0a9ba2af71b7066d58e904afd9daf782284d3cf5e762858015b7456858e5c8ba2e985d304017ba793766de2b0122280a10000f7aa301896ded10c24a39f2348e946132acf7437dbb9f1ad375f686dcce741ec8e0ef68f959dabb65086d937ad342f2b3371cde1b44bb290147caae1c6a513a747d0ac5eb196b5f6a832bf57491bb48051b7c8fc55a6ed0fd41961c1bcbac5230424a4da5c01abc586d7875d7f1b91f9b4bc68da58ee4748c7b658d8165a5b33fa64c3a86d2396752c8922d1c9598f3c795fc1282e4c1a467861e51391a07a8e5eb1a35fce0a08d65d373042996ce60c8aad4d1f3f400c88274f9bace80b882eb92db75465eb0fa03ba4606e66e274fa545ef6b519b4f84ae01ed5d2ecd0d2db87bb0b96f8770350fff789cdff8d971b18d0cd9db63c1891acc38cbc553bab2b1af640dabe3cf5a7ce54bf4e010712fff87d0360855504cfbfc52609acc4054bf1c8219d998efff5b45fefd5ec1c6920c9506ee2695a4b895e8abfad4f77160f2512ebefc2cf2e3745c9f4837e492cd7599b020aa91368f9a0e4d32ce0a8a5a1ecf63745a7f7b3d837d468a767932edccacbc2525ed13661aaeb0491ef6e33d21f2da6efda4ec2a7563d427088df95898c57c60dc70d709ce4bd17af4e9479c9fa069cb3d91d98edcc0ebc51bc260591a2d2ecc6c5dbbd92109b7c6be27da3c2cb7bdb3d295c287ba9ef8fd4ec91af7b5d09fd6788631e822ab4eaeb664ba59b9f159345de4fba9161d7023a2f5b4448a2d7b7679aa9ab4158492b51fc9e4b272aa6e54412ae219ca26ad92acc54a2651ac3b6b2ce27df9ff54465c1380695435063faa169ac4e175c999792925f80591dd5326c42d961c090a421291b7d905ecfba23518b80a4bd52e33120fdb18905fb2928389221e141a314d201e51ff660c39da0287cd35fd44aa849d1413187ba4c054b5bdd4663c1f6ce596eee952953650b1a60848124c2e6086bf329a2aedc67fb5e5e7fb8fdf44e611bd50450cbbda06e9fefc7a9425253fbb32e422e024e3a3ae177f86f2079ec46e4b876766280440814884586d1ad9a8f1bf69df76763228612488629ffc0eac6df10f05ebfe3f8f7682b4dafe72f09d954fa4dd65912b0891def9bbac791d7b7dd30f46f226698ae02587ac469d1fb68ab23702e32eaa44e35a27d584b92b8a3d6994d9c56681053b74c38efe3de918253396b570bd8d1700e660eed02a73ded599b386659e23ef07b7faaaa4a05b497e74934271b2862a93457104abe07a3156e33eadba1346a39fe9e60e98bb007fc6acfee99616315a179f5dc2b5356be0ed9977c7175853a0384ed06eca0c87c09a2ce4dea0d63498c1b32e378e5d64c41c98ca6ea6c7ff2f622fb20285336c68817e99d9d643dbfb4e357bb4a076c5fbaeb0bd9c5ac0d4e739f2a484a179385997a67108fad25a4d7bed44920db0c9f739f4eddff77664b4ea2bafe3acf209b52c9b64478be424c581b2f57f16a9aa58046e5a8e14e7d626c5462e353cda7ad7dd21d2196857d7800246b8704a515714d62d7138ffea4c14cebc0268c0dc1937502e9ab905785c013834cc1e0ac5c0104ce5d3421385ab02708e2ffcddeb8f15d92b5ba675f518eb2cfaee0de81f6c54a8c047a310c9b9dcd3f522067c653649dae1512758ecf1ae4cb67bb6e199a8cc6a6568f4a87cb4414106a6de1bd2d8f9bebb36e23c91476b04adfbcc2b87c8d9000f42d723932f2a7092b76e4f3ca6c4430a52fc4182abf49d76a7c28439d4b290e9875e5fb9a48f0ff14da49ff3fd161890d301af9f8905c5bc9465e3e0ae924ec6c675c63f334213a6d1f81542af1f0d0add6454ca3b01d1813f1b0c71b5c1a9da433992eb9ced27b491283f0b982206b221980255c911973c299a14d664f5f07b2f9dda4dea58b6f6ac790baa7424224ae0c11acb464117590131201e62f921a5186f380d6e674cfc7110504f12fe37fdac6796aa5890049ded31aed45cbb6b6d9d6054cb40f015b6cd8d9339999facea913cb29307b61b7a454fdc8e78dc4f8ee4ef32ad2d92f19671532e2660a66a7b87263fdd9380d8d477530ab0491309fc8a25d5e8d794cc0aaa3869ed2c50a0cfee1c82d184b35ae88edb5e4045376b25696c4422fcf3c2ea954acaa3395f0b083f113b4adc55da1c3fe1cbaf32a7b094145b3d2c71e6f12070ff5567c480c92b4a4cd69a2cb2a5f1dffbfa77161b4fa1d71b8285f34947d30e1ab08e96c8eb5e441f4cdb184f178179422f7327fa1e80bfc1ae0dd0bf0a3c167d44bb1558340110edbeda5496f2f9a4ec0a582a3e5f2441203f1181d7faf6993e8faebf4bb36ae963ef4922a5063553f6b1be41c503fe69765c8267e3fe58a0b6136eb12a771b88360b205055ce8c319804462d0a5a82f6f6ddfc2791fbf544ef45a507684a9d445fadab4d05174d99c71638b7ea1518e7a461e9cb70e3b580afb9d4220a9fadd162397be994be87fefeb3f24d19a7bc2fcd0964dfdb64cfb8a0773a6b9aebdd845ba86fc706e3fcb6c98be3a7f1ebb4ca0361ef0fb718ef642434f1d53f6bea5a7757e675d7acc205037716d1124bea83cb248e379e2d364e226856e1a2144b19656fdfceb683fe0381d0d25114fe5af957a2b376685bdded80ed7d1e34a72ccd7a7543bb2acbe76e958a54b6f143bb27a6ee;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4e6ba137f628723fc6b1a3b2fe96d148446cfdd0f610acbb9184981cb39b608b352aeaf79b175f00bcce12b02b19be3aad3e4a42c11aba24981095a12fe3cfa4c8a024a11bc91d72fbef61f68789e804fdd62ade21acf76aa4a2dd65bcd269c783760bfa740116604ceb4b724d3af8a874e88b50e300028a335c1df67f18fec0cc46ee3d18c46e2cf4a1aa6fd0439b15059b1ae5845ab6e1b31098f0dfd34bdceda97861399709448d672262e41d97bd046caf36e017b1023eef48bb17ead4b154c1ef0d8f8bbdeb55a4ba49c696a075b866a89b7fef75216149c6e23d8a2d3a49cb6268535184901798d7bceff9d34b2da0796b0ebc007b9051bb443325341886dfecf09978b22cfedd3faee459eb9a251120f8df4c92181b26ce4ae32daaff421a8c393e457660107248b29414d5f96a76ed230381ffdb40acf01ed166c93090456c90e75ad9bddcbd052e6d18c09640390202bde90829352fd315d46f09f281ab4738844892ab091e7742eb7ea3d152de4f98a35606364c054e0d9c0aa169ab16d862e0844fdc759cf4dd18a935253671481848c499c379f2bf42b450ec60663c4d52e1e55914ca3376ee74c5a18aa2122d5a66a6f90149748cc3da649925a8675bda961051bf19f5c03b62748c74866209fc8bb0abde0194ba63ab886981edcfade0a7864575a41033f8fcb220e9f34b7bbd7cff51444376ab577000b706890441d313470c8eda052290b0b59f9ac10fe6cf2d3cf54bd63882b1bb64b914eea077b0662a6252fdaa6a702cbb63c8b01c58f9c65115452dc529ed9f51fa80b429abd1bf75d3aec391b0089ad1fc206e691dd98da86c60895d2e43d7446349d242b3291dace8b376750a5d92d3dc2ac81760f8f2d3d5b5107e02a9ac9ec0c30aa196fecaf86ffed76ef2f3c55aab5fead2e4bdeb878cf88ddeab27fbe9d8a73ff536d162aacd2fdd4d952bf5924034f0fb93e2f08fcd1b4bcfe7afa7ea0f884ad09425d2f37bef5fd8081143ad5a11a177615a8abe4c7c2bb465bea5109df9e8cb1f9bfffbc690d6a7d4799967bb6398c308da1e456a5c3b8dc5bc3a0db8107b122194e828f493162f3d46a2aecc1e4be3b286beaa573d9a344047690414be0295f0782f0d3029d0ce7236608f6ea0009bc111a9d0d5c21c5eb938059eeb5bcda89e8010f905e423f75f69f3a3f7c518b8054ad334865b514d1424cf7e45e30379f4fcf52dfcb02665c4266c5b77fd4315b1b783a6178f4e8252b2f14e8f5345c2d1eaa9498c75f1791b7a8b2df83a624eaeb0871b4feb04098304f1ec41d9555b3715fb9637c13dac02a96d23a85afc24bb456dd8b667feba7f9bb8edd21a5f26d520f274e188a7f263e6d5a8ac7ac072f95de9f0871e5afe76d4f655b65cea2d2ff08e46d26b79b983fa7a27d5aae55d04a3b9750a94fdc1cc62bfe83e75722ebbb5da29f135b697a5d52b9ce78d5e07a198410c9cbea1257a35b8e67fb86c8858b1f94926ab41f2b11f656a5923c8ca439040cc63db8d63e9ce2f94825caaa35003b3746d93f88a4ea48e6a900d340e38f6c7e8f88acc4bbab85e00ee8c72da37a2af32d99bead03dd1a9bc4aaa2aab6dd0aadc4143c0138e2fd66347cdbf142f6fecda799f0cd9472ceedc55153dbfb9a8f490560586a19f5dda3b9b9bc3679915e6c28d34dad53a95d93acc194dd1ea7701972308da623f26794dc663f205704bdb729a7c94be0a01112f99ae3041d389b5ce6bd52a6541a29cccf178e96f1ffd473c7db616eb10cf5a0ddcd373313ddf84c2444721a37636329b8a39e025f976944033484cfe89d85631c462191e4539c68708b713df5bf16a423146c53d04567b0bfd0ff56076195eee2bf9f035f48a5197610dfc85968168d8dbd16174b4027d787cb13ddfd5aee0299f4676ffca34c975538ff759be9635a1be7f98540f66888bab0e0ce01b4228fe163c08bff6ca6a7b5f42ff80762a4fddd918e367cb648eed10b0802f2bf729b523b0f2f1bb16566b0a630e60dcdae8c2df52ac8823c36c0e40fdf995ec298946568e1587d9889807d91728a4fb658300ddd3340495d0a1c64d24c4e1e28a4ea1e3260b512f0feb5e7aa6a95239d1853bd252b403090618197dd7f2ddf087c0139549cf0fe5d69882268717c70e29ab3121898c030b7daf692d16b662ec98a5587213023bd564817858bb6cde29a09267f88357f72bcfe3e090011c37bd4b171afa47ca3dee72d49a4ea709253d744f1dca6fd1cedd789a34da390a13e6ae286c983635f1e91edf11121cc5709ed1d7886bb0a9d7fe1bd12d91ddd3f567243f7a65e9d14a3787806631d6fc95b3a6c956301add5c7cdbc16f7c64285602b57d65cd09a7b6a031ea7d7dcef2735f88e8734867bebaf9da92666fc85f45d1e4758c6d463e143a41d37ff6dcd1ade3e0371555b8540571a61af02b4efc5dffb50c77c4b809f3d7346872ed48309ff1d00d9fa9a469a70a1cf99195cf184c4c368c453f49bc0389ebcd19f43440f45de4088c66db8db4ba7a716f3f6e70f75d657a11730f0544e560ec6f1038a62971db676da45164c6dc8532751d2347a42bc10ff78181f73f95a3442e0b86f1288f34f579dd114242420ae8cb56ddeff043453e7b379b5de96590595c22960033937a89d1624c267d94f63ccf70fa71b95647fd0567855cc818a0ed8845d95ea6c68ad88a9ff8c2b4fcd765ab86364c329f7390e82c4c86ce9f47d53b975f514a0f44ad6cc11be2cd45b2ef30d6ca48e5230e651ccddba8f98d307a2d53dce7fc36cd4e9431fb6ea61b5fd9c5e944bab9e46c7e01365573c83e647307c9c93db73a1d5aadf7632fe0814fd65a01b401b2fe0f989ec3bf9c1f905a4f3fff9612b4d5952f3f811f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5caa1ff2b056a6e43805211b57d5334f00be7a8032ea4f2f5b8e1650e6527850bd3c0a9ade8e3b510226ca3b44c23470be10d5b533301787ce73d303abb7384db2519846236995245b110c38c13066065ee0dcbcf72528933fa274335e50514fb3e5ae37368cc661bc27a1fa502970c4b43daf286fdefd99ff9773e7c445759a8b9f9944e2492792f8163dedccf977ca580c3d562de3c33ff4d83f075fed427c4b53d6f3cd83c079a8dc6039d8eaea81195d8af373891ea5e3df1738637756125ef2e2dfc3e5e817eb21bd436de86a67455ab0bd0c218f7eee90fd93315cf3b266e0990a04d8abc05577fdcc56a122e0dc51a5f05925c2d393d7ecf1961747f68dab9c5ab42696c08a2bed49f1ddafdd00c48d1779f998bfcc04c2a3ab8b127ec762fa27dfac7d6b6beddf6502a9f270c61ffbfe90f1c6aa74d77c6e3317097f90f7d20e3a91da9ea886ae78c701315e5851dc26bbe62bbe391e5bd853524d77513e490104b9e4551032076fcf73b25103f5082386bacb32c2968e80e30a1edd0fa74c283a42c68a07b91d6dc0857bae015bcbe273f317f17b5de829f6719cd8b5c3bdf640c878bc3aa87e45fc41f70101d83e1fcd304161ff7ee8b4f6193011d6c76617cea2d8e9fd8667343eef1cc1adf978d9e0c96a34c5b63ba3ab01e853c8e41677fd2078a26f3038a3ef9c222de8083482bf28281f55a7ce12cc2c329c8e4d793b9c6daa331942717846449c4a266120ed4d6818abb2a65f0b230b0877fa06d0b3112cd661b5fdec6481c0e77d06af9ec375e6f8f5d9256f56f0aca976376c67b436ab9c665d6033d0b2bdacc55f52b9a9e044ab5700a3657f87c1ada9d4d6faa057fd34e356ce39dd1f4bf34c08220ff2640767feeee5923e64b899b1871e37196a7f693fd0b69dea6def7063c1d3914e92b288a00dd1a465195f5524d914feabfc8a27e7d7114c5fd02d32043c3fb11f7a22724f20c2fd9d69cc1d997a988b57dfeb83b63854f43c165681bef56dc0c8574778bb93cc911a6629877d3be874298603b15fe9a286126d9d0678e583b9509c7640de0e8b4d59a3d4f8e0ed68a63f29369dfa5713ab5be7a4f5791e12f64684993d9b398eec53ab222bcde1333373c2873b1206f22b08586f5c1889f0f9476cb36a71e6af61313940d65426d04d1a56f6a67f18cfec20d382d9481f0d8b54badf110327375c300dafb1e81449d57b2d6f1cd2a2d563cee511159afd130a97da5ee7bb976ee9ee70c38a0c73f8fffcc47379252be06f53157e0ea023efdd3e618d6e3def2734f41034dd4757b638704d4789e14056d63033351c6583e4c9455669cc2c68ebf4301bb2d077578825d1818b0853bdff4dc1a39cd81ae7baeca10fad1ca923e6c2f09b8499e9d73b1130b526f05878bb5a167c4e39dd654cc24100101a42fa9737499a6a3dab064a2782eff65c053be36f5768b9d3c3620e22c0e2b7537663fb993d55c852c11d69b8eba98ba23e8cad5c5cbfdea805209bd55ed0e612f5fd2c8cbf2fc5c2a721234da514727560aa217ba1c9db28ad9b28b8c5ba44152bc34e0082e7c8b27c75e6ba7a07ba3ca8c1ff0e562820f4ec72c184b1ba25256703e8c76297daa58bbc3396bc1764a2cf90ad5ba451d51652c8142b29f01f0853165700bad678d6ddbfcc6d80cf4a622d5702c9f3646288853db28e5509615d0cbae3901feb769cac87b153ddaa930f59da607e80d71b2a8e706640118dfbd618d67d928e91ca46a7d808afe6a6ea35085a23a0ea3160aaf24580ee03291d274d1f8617390327efaa128e63c185f3afea66a303c37cde465556a2160f6912f5bfeccd948b0fe4095dd00eaa2f6304f9b5730383a84c234603b9890297f159d51f2e91d55ea698fefbfb61008cd3ea1787e9549dd876bfbec20c63eda38f4ae6134f0fa71bd126bc26eb2ffcdd75ea40efdd2ed464925ae74848d634b68c5500bad4011b728a28c4b2fad314afc06f08ec809efc6a9369f113e0c6ed0781344f4ada2fe17b9fe5112ce18efc6fcc0861bb146a9afd58eac632588ab1c63126e8a9cf9fa5365d9ba34b71ad866c6717a8099eca228861d2ee98b5350801e21987ba515ad1a3944726e815a75033b2fdfe0bf3a1d912bbeddb5399a28cf1fc74d83615be157b584082b41d6c796ca3ef5a443515638f641fa6dce627d3d9ac9a0a2a8b0f873e04a29a816b428295680cf0ba27a74a5d2720a409149ef8e2be1bb373726d099f2dedfada092e395fd98b218bd1afad5fbabe45b383e16f43d3751bdd73d981814d71a9ec087b624fa8560488b1b988444c59b4a77a18662056148874569bf5fe4caa6c23a9e7218aa805f95adaa093da3e9b01f60a3a7207df94be586f649ec01ece682a2aee5644eb485e0150b653a83697cef7f210f9730a68542b345901910440be035df3f4dd183318a23471a2d60bc7e3159b2834e6de8d865836a016b48fce2e251051be03ddb345a314af3fd8721eb65466e740d182612007ba271cb7122d069eb5243d419ea1d519c2f82fb8fad3703b69d95b9e0608bea6b5fc9ab2ea0868e3505c7c009894a3f27019d58f20d2a20842ea966dc2da0a43277814ea27798acec9dfcd0d9d6b87965fbdb027ee15f863b7ba1b480b2c6be639955aa47c44e4268cc3244c02cdb3358b65cd0ebfad80790994a8385ff0ef87287ba044ec420ac32accc83375b78f38204583e589b87b7e643f252120102b2ee0749427b1d934c9a11a5ac7bc84e13bbfb5fb3e4827fdc84164bdd918d426458cd8d35345f3989e857ebcce7746cfcef5da365f4c6954432dc18cc7cd7f3be75623a9ca336b89cefca552e3f856f4a2c87a43d221611ad0494b12a076115640284610b7169c4a44;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf0854d2c41ed4d2bee4f493acdd121b874fb8416eee5f317b91e44196518bf47507c5ade5c872b249f0169e8b1e2e09a6576f5f6ee2c7690df112a3492434a8c0ab835594137c25db1656c665fb408e9ea95d03a128ede452ab22add4b6e79e78a4266734b2f5b67e4c14e027f9dabc95305306fcaed858fbada4cb7fe9ea64ace352e0b84efaa4fa892355fc9d4dff82dbc9becb33f828fde77bc10018f81e83c3537e36b9395e0a58b7a8cb7836221dd5fddae69a1ab60420ff444000f1ac12c89103885e0a95a2e185ee65bb75f99a745c03cace84b8878b3bd3df80e30a2e0dac381d9430880b44908b2e2f411e9ff949063772e41685e0351b8be267e1946ce4d2641bb76664b1fed1fd8acc16de909d5312114061cecff58888c93c35ab88995fa01adfd8edae08cfe1c1ac39177f7aa53bc6d511f33b6adda2e803ae4b5bcc337cd7fbc0e00c3a2db53646f6a6c46c1206795b89d3ffa1591b07ade96f896d8c1adefa373bcbeeb7bfca4f6c130ec1ef8a94856a714546fb1cfe757327643a490eef8580ff9bad56fe2f56e6aac03580d867a46faf6125860961558a9ac85f775e0a147d0a73e3b284b5e17ea70936cac7582f4c2ccba8d0fbf2f03bcac1b01b16166c3d5561ff3b77669c28c1fabf73263e02d6e48d31a4b7fe94d236c9de5f688cb44a479956f31d62f204e808da9fadf9145535a7e6537278c617b3aec4ec3873ac9b99d81f13d70596d69f525c6ba9c398f825c5f1d8abb6fd8df1081fc16bbaa709d9d93ae299f0d9471602485eb5f85a26e793185449e8ac5de478a4888c45ad8a048da526d27ced7aa3b7da73c98925d07c4d3641f59f5ffcdd424bcf0cb9a3a2dc3a35333ca0418af4f1ad88fd8d4c2733360d45b92f12b72800a9a7dc31ef13fafb5eb5d25c3b1071319a13157150fbc91fdf49e6aa8a8844b965527589a9152239f7f885c4e580928c46d87f3ad62ab7212d1de8665565c0ab48859be06d8ab5b9124c1bc31358676b70e600a853ad17a3a7dad051ba68d1ec1ee3a7af3cfc987636448f145cf724a28203c39df92c6e7d4108b685df5ffe7802800478957bc5eb9f217bf57eea63069857bb8034f579ebf9066bf77db3f864d0ecb7671d6c08702947792aa2dfe02add809c51a96952f374a60c712c669f2dd2ba2bed91a64a6067a73b969c06a72dac446ac897faeef91f69447de2fd735c0ea73b1fad32bc403cd79fe8e5243b62971caf521388c69e2e2eaa7ea5b8c53b6311dc6a9dc5c6796df3bcd6e888dd29b8b6ef29f40f09acad446f573326104ac6aa57781a8c6e3228c60a0d019f19718a0aec0c1136f88874fd123b19292c84ebee045ade9421731133b83d76dfc6fa954be7837cbea6fc9857e0e437bdd94654de8d7324570a725bafccff2a7252444098727c32fae131479750d81a5e5da629fef3e2b2b8b14889ecf6539c173a0be261723219bfa1b88753882efdea0a43bb67840ff0ae39b5b0ad4a3d60f6bf59adc3ff0cb7a0d4b0f956cfcf9eff0e7fba068676ed094634093566fec2789b444801e6e6b7ccbec0e889a36126766e4630cbb5281e37bc3adef9fb570dce8d85b7783bb47a59e9bef78aea6967c23463f4fbf3ec25f9ec1d05b7a20ed612222c97f7cff3ee17feee3676a2d48cb09ee97b71efdfdd970ff00bf1b906b527ce6c85bee01b4a8ff30b74b1b5f873e6c0156d678fb9ad7b07152a52a6e61a0a2e66bfc99a01c28295ee9dc566e957c426efc14fc9c97185e38da03739af59ad9c071d24461ef6e60b9fc337625119b5b2ad83886e1103334c17a9519bad96159cb87871fb68246e0bc71a983c907ed8f1fa88ef7817941c7306f61be53c5335ac33d76855a26857dd124d0d817f835c440e30911688787ee8ae747a61a520b22d6dc54d691aa9659d00df08b89c7aa812515a189891f11ce8bd16a6215a360bbb0ab149406889340c5b7fe584dfedfdce2b1bfd48e159c02ac50c8238f4011d3f3a78d872c63c1851e68ead9a7a16a3521a8a7a216a4b4d584e381c04433bf59e9ba12292417bf77d2a599c05f92f4eb2bc65f1889f02805fa67193acd26625db740f73b3a783078ecc3568422580d63eabe3467039865679948088783e377a5abdf146e56de07a78f56c8465e0197b1832e50af9f3f45b4c24af32f908feb503ed0b609c95ff2874abe54c7bc60d0eb2584244cfc54bcede07217170519ebeadc56edecd4ee59187d6c6d2f8fd9a929a41cc461f5e34695af4347f742ac4f86416ed4f9a9e7d4f45fb0815e4f9aa29d636515b07a051adb78eebe783416b3ebdb0103c5a4e41ae9a22c2f402776b007a792c0b7b1f9988559dfe9e7b0b0d8459fa4b83965d862eea9c8db0f5506387ec1b62205f8871ed0889a2f50c128a7be4e8fb63557a9598265059e7ddc70863b76b8847380a4038d2fabec165a2467d02203eaf34fd6baf26ce29d727e0e85b51b2bc10eb31da9b08bb2cfb6548fbc7840af1dec1e95c078850af5aec00af5514b63fa6cdccecab72d91bdc5495ee28c6407edaa92f3fba10a0e69937830acf3577a8cbefdadd1cc73ce67ffb1f6af1988251fb0496c60cc0976e329cf96043ef144329692a245fca455c254b37a8ac46f99e2f6ef435f4b7a5e4aeb0a8a2b72c7bbcb53a81616ced5059e5f678d0b294cefbdac16c144dafa7741a013bb053f2113163068315a04560e74bf06c103e07715adca1b8b42f544d8ad3d79dc5c3fa63ae0c7b3c69f747e1c0b2d75acbc9caf60f6b30094a81184f9d7609907aa77caca1be81cb5548d4589031ea386221a5af0facf3884f71f681dbaee3fd35a2c1dc66608f796118df392c552fd0b4f4223596449c71b6fb872da41a2fd1003d7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1c1c1f2627de7a410c567a1212d18e18a2c4d493a7ea5def561f5d2ea067d891c4249d783ecb7b337e50b3c63be8bc91e3709bb2a678e396b39f4bf9ea427abb459e54ad583857a2a53c03811128138a9abb571edc2f084831ce48f83753eaa46306b30444a4df93494e0b32103acf5791d055673e70f3cfc2ea8fb6d74220951c2ca9be6b2fa2c675b1cc40d7d6840d1a0230c547fd2d375774b64ae89bf0d4059b09a91b4ae852a1f1a1e0ac521910c1ba0113539ebd573ee2e7a83aa44fa9b77f9e4bfdf3a869807a4989947b2e91c17198d6e7b5ee6d94816cca3d94b0ee595c7923745b58a73bf47bc963ab040924f99bb3f381be0b61887e58a069ad89b611a9f62b98b3c82bc7e52009de8fc155082be008ea55c98974f32ac838af4b684e1e3ca1111349c6d0ee774b95635795ee00358c7a308b2cc41ee34340d1ef7996efd2f5915b316e6ba58c83f84e73dccb9145a691e66dca4d8adf8edc62b6fc5f5d917b2e93bbf158bdb7b2bba0eb0be1a38a8c33ff27e36bac29aebf1e73380a3d5bfabfa1081812b9bb5551502ecbd28954d3e65c7438df524c7e3f4ef9698de383827b6017f0ec694b4d77bb392df2f29b540c228c0734294d3a8b7e4f0feeb06c13b7ea81639a1683f9599ec8aa24b048045990d1e4e687cdf5a740da97351457ae3b2eaef1c4ea498c81c5dda06c3d38d8e83ce463001786b8890ffe528da5ccb57c4c8491a11def6d39905c8e1d36b89c9f2bf5bf9ea8c67478363d3f3fa1014a55986e7fc1f3cba55e5cd26996b7d579039614ee28ce34393922666768f910f65c22db4f36b5a746c59f8c76338997858f2c8b8ac418f9e7bd5237d3ea1dcf5436f90d50de002f74afb2f80782f853c9c634d9285ced59cd5a77f07db889a4498e1f63484cb023763db8d927e6371e60c64593306092f4fa46a01e5dc47add67b54010c427a350bacfa8a7e414966ade5bfada318977a4e7f52963455587c5e7d21588f1ce43426338969b6cfc09c54e68acb668f4bf24af0e1036d4de9f20693ac28e958324202fad8dbb367eb645f439326f506a100d5f41a4851b432d00cb8e532711c85621c10235ecce02a90a1f71f077f555713b9825c849141fac0ebd51bf7c7d737d7b98699789e9e743ed17845c008cfe80a08b761cdcdf4d345d29f0321ab9ba2b88cecc4e1e5d926373ae2d9df28ee298602766ba7e8831c6419ede11284267d2620149b9094f26393b244ecf1c2116e46a308d257992f164af49df98f579ddd2bd599621b3c00e0473d889e21a9de7727e01501f6577703c8051c448c38a3cd236559ecdcdaa844edf68edd91a896a62ed509c545a1118657860cef56aa3cecee6b29d49221d05732f5d9c07000fa49f12dd761805b907d0354c9c9bbd4aa05b39a23e3a5bc2da558d85513159272d0381809453efc092cc434990dabeeed96c4060358375e4a7082444af660c2723f37ea803048997bc0c79093da6224e8fdae131f03e79796380faa1ab2f5cb4591872be5916c0800fe2e42aa7edd22076d7cf9b3ede0a2c968a707cfcd7af438105e31f0c3b8cc097b42d68edd704ec97e7100e53e8b1a0790a295b51b6d92181fd4745cddbd9300e9a9a8ee21eaa827b0741b115ee3c8da4d88e56ff6bc0f561d486dbb1f4b13e89141b9f7561e0db6cbda5b4aaf2ae7136a017375baa2882522a0858a2c4398d802bb410bf34ebc378a6069601e900726b5b7b882904a4c07dfac22a290d38f3745aee78d73608f0abfa934df6b850d1eddbbb74f8afc402fd8bdac36888ccdcc3f993898eac002fbaed914583b730ed98fbbe7cb91b9b476f9a52c47f6607ed734da8df3b3c724b9f095f54c082195559ad03eb8f0a0ffb889e1d581983c823235c4656fe41e24958285aa85b953d824361714ed83db5b627fdda75b83263bb70365e5611ee98f915056ab3b7cf1d87ff288f2e3ab8ae3118883008a282beb94f95e5211593bebd61b448c2aef9f65703fc4a390bd13785ccd28a20512bd567818fe51a44114ff1c3929e59f6cc547ba87ace5bd459d437b1ae5abaf9b193b946368d7ce9258aaa732bf600f25f74e566de15bcb34651adf42ace4ac254058c2db62d87481dcccf7bc152b8bb7aa996fd9a3928a707add2ab66ee1dd80582fe2dd6241030c9d5186c0926cacb4442b1bd9fed859e0e0fc7e6c700196a7d3b581d5c65edc9c9ff0a73c4aa1bc482d140c9fc45d5de7257beebeb0f4d0b961979e7d1751f631bd9c1b4c52e3b805cda4a7a5447343afd23439466f771050ae917f36f8a5ce2ab5e6d3cc18bb7a854dd8e34587a7e6aa85e8bad59138f13946f75bf419736a9feaf5605137796e90b1f3a23d92902b6c51ae1acb1374d21378d7249c7517f02bc94424cd0d2a77885de66e1e4c14d633972bc5ea1e7904cf9c058f00f05a762352bb8cc590e87850420b8d1e1964f53497371b5067f18d9fea03ea2ff5f36cbcc3ee7c7689877fa6c6cbdc92db4607639b16dbe1d6acea16487afaf62cca33d912924d1126e43ba305c216c5a782b58672fabb4081e107adfebe9d4e7e17dab35a1e26699d929d698a7735f8f309676f5892ef98de63517f3fd79f29a3a844c319be5a9e0eaf46e1252adb084a57da6310a81307066089449f56c427b50ee3481a49e4cb91637eb35b84c314b6b53eb4fe8fbb40517a7874158ff46af2c0502102504e4a8e494384d728d0453e37960fead59490524e1dad077efc5f030cbfb9f1899b7a8d8f4fb49ada83bbe5cfc79390b4320759369ad1e4c6ec5e40ac4e9598e8a15126c13e529590d0f795cf502d68a3af54296048a521848534610343ff8d44b7a0851d8e888dc2b347065a45d52fbd8a5551641a9991a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h390a8a1599d24375d7959a12cc9617cdd393eee68121c74760badf0c77a90349a13d14c319f14e37e540121e26235e1258c193db3cc679f2ea4bd79322ddcf8ea3bee954001c3fa796ccabe15b0b943b5d498dcd5e916f66b2c838469288fe4c2e56304ea47386e73830f3d3e2bea60720a07b61ea1c04a3aa0bde402d645e906f0a5ad645eea7e95373c451d633ee607dd3ecd01c10d50ef32fcab12871e842e92c5e1664cc9b332dfaf26db19d7e10dc49818bbfe093ad7095ee70ddfd48fcaa830aaf01faf65d5c121c6aa17f5cda7ac4326b8773599f5ee8be9cae030a12ffc629899fc32e0be10996ad006f6ee801c41faff87a0e194875c1646b1f8b3640dbd8fe805102d462f0884eaa6f488a697414469fa066c4994651885e9786577f46b0bc319e22a13425323bc40ff4048372884b3d379f885686f0fef7c28cb8dc9c66b6ceb31a0efb70640990bb2ebe6728273b1968be6f9b38ed19fa4c51504a19a8436725cca37e43f0377034d5837124de63bad5d64e338865e1337ebea374c7c6716c769b9b11e1e63ff56d39bc4c96a3902ca93ead8abc3626f658148f990a9b84699e889a92f516600b2dbc2dd18ec72a66d0480ccf381645e8a56aacb16c705a4637b71e3e10011a1b24847f4bae92ba4aa41c2723bbb8361540857aec7bdeec939595f33024cb6eea5ca7e0e38700388a11e2206844ee92dbeb399bab4c30057fbfe62a78e6d238563808155440689708d3a329423849a4080a502ffaefc6f1087b953110a0abf7a9f47d899499848591a3efda0ee92a59f5b678311abbcb0cf47850d9a1391d827b7a6506f4a585f9eeaef6312bb40dc5040c3b2a78f594d03a8fbb172891a1cf9585462c275443fc6208e6eb5d3f641b62aa1e9421509c8bef76ac27854172c6bea550b9602d77fd5d0ecb3f7761bcc94a14a94eb7f0a1c7cb8afa06d5ff74884bbe74bff7e9d28c44cb064fb809ba4ab4ec6ae8883cc9e87496424efc84c8b0c356bdf05429bba66f76214b1f56d545b0f063f7e7764f046f3626ce3810d57ee61bd3484776df9e24a5d3ff9e3bb1cab3833d6fea7f161b0e553d9b13b9781ff5804ca7073b82bff31f7a709ddc4e75a6836530a6fd4b4e89234ad33e1ba7affaf6b084e3d13ffacc8fbf1e87467a5c54009eab36d20d9ad74e61987f84e4fba55ec0142ffc0e594f050110185879b67e061f358d8efb4462c0ea809200ac44ad633137e60bf243186d269615073065514b91b1b6f946ebffde3a62bcd1c308b2ab7e88bd1f71ecb0dc96cc3f3cfe6d2ca31a4d60a17485dffa67c7f4a679ad813815282c9ce396d62cfd476f958f72db3b5bf8b4b7d3923d9d70709f5ee9cb5d12c4f39eed34ad449b2a5588e1bc0b68672a70142a02adcbeec0ec30c4a6d5d42d0aacd3750becf261fa806f9ec7fc370d9462c2bc2b3c9e9401942e732d2a6e733b8a24e07b0959d302ea98a1c4cf10d1827eb3915a313777751fafcc43e08621a25b075c21c7819ba6be129a5dff4b861a36bac816580d3e31c3b4dcfa20dc94a7ca20c44d8f1385d721e905a1e1be1ed840a3a2bbdd73e1c5c405637e66035fb1a6312aff3b97390c1ffbf4f62c4a5fd2fcafbd5226267fd2ccee557d8d36880102c35546a9e6806672f178402024e7ae22d539d806019c1b28af6c007851f54d3a91d215d8d147a1b592f3332ba5dbcf4626f666f39e48c4f7fe3bed24fc4172e7db4a1f7d05d5a21dd7224b2f2fa6b20f047e0ad749f149619648798bd8ff4c3a68c457faf86a23f9faa5016ad27c3fce8c16c718d839e52b6f1f11e8f0fe156d2942091a4ff78c80e208aa270bbd76dddaaafd02e6e238d642829d3e9149640a907db8d54e42a1387dac60d4442828ecfd3e8f45b6ded7f90a4043759cff98a7e352f30fec4e48aa61ef7b43ff7e70c7a900b5e043e6a863e150092c0006d57be6162e9fdd22d8f9bd20b56ddb7d703c84794ea5c52ba26b965ea0f7c70f9a66c233ed25093071031c5c0505ce86bfe73484160f8502519aec7c6b4ff1d11ce20f9741873ada3fe5e43607e7fe46efaeecd9d9c5b92f1c8f7ff5bd3b59b90cdfe3deda602621403290ee0e849fd408e38d75e688862343e93e722edcc9012e8c058b090e11c47b64d6e208d033360a176401e9f9e5716edc25e035f7064aa3556ba99f2e9273bcf9f3b8e63e28296954738c93b4ebe8b5dceb703e3a4ea39c2c82e40d8f184e96d2ac8c1e9d933ee9df4430fe8e67ae98057d62b9d976437800bae669d3a8c578c8a8379fd8855b4ecd0f967f6dd3c6fa11909c550301a64ac3000e6d2a50055095f07ac7dcef2cf4c1a095e689269523fcfce9a9b01ef220c38ee0c85db0a297e7f651caec305f3a08ef7c3d9b793a994d1ee79688d582b745e540af740743b79f41c676a52b8db9875f4b18aec5224163b987c57d9530ff6976d2dea62b9ea1dc163033f511e4c18d64d47eda3204cfee4ad465b7980b8af14da9a806cb6834ba9809661a7b19cfeee13efccbb8e839396536564392f4de58ff431a6ce8d4d5cde05e42d218bd532fa4d12c6516b7619609713e78114abc12150a76f6a0a52b639bc3362788f5d4b37fed686588b49cbe834aec4b63184aa9e461a3a20ce57eb765d9691cee6bfe4d91ae4c24003b12e0fdd308b7c430285ad584a0752ff39d4295de2d6cdacec49737ffa7891ee1cf5eab720b8349e0ec77fc9024254a54755aecedbcc8942b7f511e625402bbcd73fe91c30a7ca94c59b9726b8810e75a52cfe865e339868a236ee107d7a192cd2fcf437523e4a30f7d5afd66c3cab396a51e034a2232e218e2d6ac976d8712c26a47b1dda078e44ee076dbb331989813eb2e637a7a34dd76c56;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf7c931ad8453d012aa66c9cbf58d4b45e13187d82e0caa01cbaf914d43f43c36538c9649b9c1a2b801b200d2b13ce76946373dc8d6242356a2df558c1e22f1524f71e0b6ad2666fdb82413402852be77317b22973c1139bfcd55e9ec6cd49c765c6268893c2d626bd78316ffe92cef39f7337b7f714d634f405ef11e76cf4930203563a99f17f5045a41750f62378716b7ccaafd7fd9d99d6bfce1f04994dfb8cf41825e5180277bb26d7cb97ba0eb18dccad53a2774ef10a71a6dac699b786e3363e4a3f1a2a20fd0d27d3e06977638b126387a370926eea948843d8e80b1cae79f1aeca010c0123c5c2e03b9e1071a56b10afc7a8f9b4375bcc3b2bdf7bedaffac82ff20fd214ed85a704f71d01b7c09721873c7e6774aa63f863f3a1132aa28c39c7f1df1749286e5fca0a2a070b24b2e184e5d59993b79df7f52c0b1bfaf80b42a01706c1425ccdbdd078ea04e7361bc212070cfab1bbada783eeda5c0d35c26c99b9885d70016e68ea38fe40394e1c77c6b801d9fc8d5c56fa5cdc3ea1979a1cbdce8832dcb62bfa5137724993fa38676c06c909c8c7945cf7dbb59979f34327f66ecf3af64cfef6fac9ec1b5f3a0931efac0a9238fe38e04fcfafb141aae7f8ec37119a04a7aa410fd5c1544aa67433451acf9ca5e3d4a302963f06e7cd8f593d1ff0121d470422561e543cb89cf37c996bb06c623714fdc43cb69d5c8c1eedc705a062538b052ca64bdcfbc28c4af835271bb23c3f8d59fd32c52f7c4120943e19b13c22c1b2047a2279cadc6243c0c7eb66efb4b345f86df99829c257e6bf6376d16c6b6c8d801a6c2581d5af19670f85b1819ca3ade22ec9b3c359cdb716d2cb2032452598721af9af8442107021a99f31f7bf476536d8c0399ae64b60d87831e8ed3fd874b44a1b11261a8e0f2f864427e1f6be5e36be96faf13f4da218830692d07847fbbf0bd17f2dc87868d53535e6e7daeb0efad1aa452354c68b5ba8bca3ef44258320b3179d6ddf097fc5be7f574d3e8c46441c066ea5f452535266451f3c5fbcc2640c99749d6ab4199b166636d87ca11044cf5d4208fd2b25441ae04b871fdf63ea9ed7bfe0c44950f0d0933bd242c2f89156c6a839fa03bf8f97dab1d020ead9ee131f90d8e6f272054da800c6bae849a502d8164c0f86ca05567ded3bb59603603334bff66f47298b1394c46227f7d23105aa27c0cd0c29a62a501edae3d6beac014f96af0428227290cc84d7ea99f6c4b752287f797bd9ed65ca8bc7a7298e3adabba833a9ad886a7a3d6fa09456e34fcdf54eb2e9a1f8a6bfc9bcc1b5ed50b15fdbbb7cbc824bc582f4a2cecdaa8a630c78363312684239afc8cfa26836aa7a7bfcbb6636aab2e0684b0fafba845b7e0895383fd0023bb6fb0cfc394a52711ec8656300b1df40d4272b14adac679169c47db8ebf27b5cd831096941f213a3b97d98102e662183f41a48442aa62410161b59b682f7aeb12b378117f4a9f5e77aa6c5cc018078de0133295dc31cb8c12df99c864ab8794c7fbe69f40f16bfbd87a8db0ba91c66745f9479acb925e7529b5a80285a907b9427ec4619cd2b71b33a98547b805adc66f0353f2944059e47bbcf2136e1d0d1ae48c6237514afb64acb5f7664da725886a955c14dc99b1c819ea755b9a4b35c392f6be96db2aba34d0c48e52314a171254174ce6caf514f57da8ad8483fcbead784f651fd82ce872ba3df2b87b6ac939619ba37e0226d59867597bf77d5dfe3164e3ff1e1eaed44c5f34588dc43aabc80e164f11384d831598f746b6679242343200727ddfd99b7d606bd9002242297ec2edcf694b216f09adb13f9b4c036a22bf4b4dec59c3ded820dc97763305d2afd6762160568d4a9f8dd2f134301e940e33697a91a365290b15922cbd89eb17e26312720c011c07b45a799c8552423d4f8cf09205e2ac7697ba323051f20a9d58369a5bf628f057364c470bb400fb7f37e26b316a712d092e59a7c2959a1b89a78e04ba0b051384d53d15ac524748d81a0fd5733e1379f3daac9129f833f2174c144ca734f2d5a2bb698f2b4ed90210e50bf0efb7384b3f788b8a170a054d8c08771aeac6cc7ff6e4ec95068235c5e5a0665f1c29b48c2ec7750d234475587a8b84a101c800eb386de2a121a2664ec05b26a5ed5cdc6526843bb1b30b09f6019e7e098e87c668c5a85c1b265678493ee6c9d341a5ab7916ec264e88f30fc02644eaa44b15789254fe1c63bc39d5e6f56f8630d6510c7670346ccb4ddfd32e540688f5a544c29ac3cfe79aaff786c9899990a234aa358c27f46ce313b0e2407beec53e071612882e064a7331182efad670d089a6de536b64d56a23e646c8473cc2eeb1992939c91f4cfe98562f896ef460adf20e880d474048fa2da53cb888daa1854ee7bcadf36a8f7b8e23bc05b7fa7c41d16d16f377d96978cb90f84fe3eb3a48ae2c9a5ea6c9dc47044ac2358e8a8a54f7f1d36c3cd3336108e5d977bd0282521bb3d5e18f4b7692c237e7173c6cb4fc16c757f125fdb1b7844eb3302f83eb4846c0d8b0103f17a9504b5a9992ab8d83b4270f03718c7670f228d86319dfd4a1e0bd29a089e3a88d6fcbdde98431536bb1e024071c5e88f1f33698a736c5f0d0d03eb0d78bd7dc797c8046761f3017868daafecdfd731d4f2a2947e46dbe4e0b6efc954457032294afbb755220aec5de70a726313c1d08673117ab0d46d70626634cd12457c99372d86891ce0c875adade9816a86042a52afb2eccd81256d6221b390e91233b32a7d44429016949fc3a9f1d6a6787c7a64b06fd918d96dfb7c7a775b5a10954778ab1ff62da91c4404723a2ec4c1596f970a3f0b0cb34795d62a7d28f2728f378397ab423fdb390;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hbad9c485108c51ac98d7a83961b5cc2c5c78698256f20d617bc1da633632032264996004c962294d54fcee0d1521ce37d67f899e0ac1266a087571c08bb933cae2c2624b8bc12b645c263e32daef610569b331b0141fa931c55407c63f1f540336b73336143744bad3f552a5782493fd69ca4f48793b56a96d152badf25e9cff7277669f35f27ff3bb328ccb72470f68cbca4834dc19c4c5bf20aa52d24038c1bd016906958d5f89477eee6d27cf5ae0cdecca4cd8830f770772c64a41942eba518255c9f45ab983c1d3c8979c0bda10778e7a8da817a63645989ae318b66bc7c69e1194263b774ffe995216526234514b23beeb1ba6225237072adf6502139c0e9ec2652cd4115da6a418611db0796af8e0c817234b7c8c1ea795b7e67e39e8eb60fbfe8bccdb3a448ecb853dd16f0f6bd1e5bcb5e6711457a18f6c54506b15feac477b181b930c102a069af24ab2f25afd69cf35551623716f6fce2a65c190bf23e93b9b2c1e4f73224db0fb32438fe9cc933089dc1b4005bd244060fe29d9f53bf65b43345ffc98b1baa3b8da3d51979e034cc1a517e3eb5df7a2663b89037a08ea0ba8d8e2e50b52d972239b87242f1a308f88d9f670cc9b9ee4392ef159aeab7258aa4a1f7ee7f71ee4a9a9fbcf533c9f508f3566d4c80fd066eb854826eef93151324c3d4499a0972a532c51c33005b9ea464616ee0d12c5a9528c0eb08a077ae391e403fae5e2c19383965af8c561a785640bb81e947c54f4a7af59c004f20a8a0af52555bf9f9ce138a59499a6f57b42f3551aaaa660308f78df2ddaa6900185ade3455ceea09ce9cffdf10d9142e893ac3e4d9757c422bab79e1d53d64bf05acff0a083e02e5545990b7f8e391b0e9aed4819834f144e52e123e0b7144db7d39fd631e107a9631ff3becd5acd8e26d8d65a3c7bbcad709a9b37f335d36add8c3aab7d79ccd77d7777d6910404f00680a25882fea788a217613d67b973a6231d4b570ca4d50fa8d1f42bf616c3eea1514d291291d0e1dd323df867dad27a5228419fd25572d67b19cf38b6f6123cf78d135ee0d51a8fa73c267b20cdbe3fbddfab80407d2c9a4f502701697b0fbe6574e4baea60361ad7b447f08b7977571de3c5b86b00c5809c9115d0938cdffd9db8c254e0195ea731e578c750a456a81dfe54a4b3ab80f3a4d4a3ce8d6396bc1129c66314df9193cd3e3c7f95831e069a7ae1cf76e70fc5e18ac5c6ce468719b0e30ecbbdcc324e130e564f7d58d1908499e3bf43cac1cc174cc4c9e0ce1ad53a2145dacd9deb8de4ed51b2ad93dc89cfe8a5c23b63fee94cedb47de209a6ba29fb5e9f476355318170e7573065576b09653e00b5b0d0f069e9e14e53e97c9674f18da489de8d482170cbb1a341f4042c5a992020ee47fe49e4ad84bc89e90fe4d558267e6908ba90e79b0a0bcd9d52c0aa6a8081f932edf3bb3d5d15f87a88004f7c9400b4948dd1aac59a3668a199690abec35c6de358a7488f27922bc9d8e0bc2f7ff0dc2538eab4ad41ed497215c4146c65a5637540399f99a80e86eecc48e7ea60c23289b9a0d392e78dae1e3dd44a44ca3bd2a9a9e833de446fe39433fa02cd97ad89e50813e585100e0e8426c0864ffa64d17a2dd944e75150c6267b09dab330319e323e00af726e896a94aea4be1a4faf8184d35b5967f921bd19db1449bd060a33dd662b6814f566dc5b6ecf4a594d1c57ed4f3bd372096d08665de570ded1ba30f26a9e53aa0a0743f6d1f61646b533d41f469d30789476114ecda9b7ec19843683010cee1d6b0bfb3f7be7ff99ecbc143f5487ecb0296a13a209caeab6a2a7c09d38eb1f3ed5bc486c92a66b90c12f038a462662d9c8d4bb6fb7f0d9c040373e710655207abba459b4da9a7cc3bc8de670f1bcbac6e9a2d67f694d6440de2773d9652fdbf88334b651b8d7eaa90b352f001e707daa9f07614914030b302d5b8fb1e13ee6056d292fdeab7e4e6a54b4f861bc4914c7af5d7e3fa0dd14d06c6c0a9cd9c7fc6242c00fe221f097823076800d177d25f93f614204beaa37db9763cc6df92724810dd09d77fce5c12868d0f5baf7431a1ff36e5c3ab7556b9aa3bb519e8cd91363a06d40fe4732987f2bc39448593b9b14fe254d99e10c9e61305cdc35811685f0aebe4f08e89ff9e033b877aff8d45f60440496a02cc219951dbd1911d54714ff26348fbc95003cd04abe68d1cb02fcbca42a8e45b2dfecc0d3733c4f1ece5eaddb8b2e734b5912c4071390df584b5ee802be025680a7f35733d9f34cca1279a0a7daed48cf347adea201c8cd5ae178ab109c8b3933631e8ce33339b2de6f09c2851eb7c0afaaed0516283fbe4a9c5b6ddd3f5e4906f393f16266f314aa359e976e06eedee586153b799798d96ec5345bb6f1ea730edefd5dee71903e29b91b0b0b4ae2575f687ffc211a6224ffe745425c69d3ae5906398cb229b201a07f8ec8abe9e5ea6dc3c5691fb7e28eda9cbdf9fd2f2e78dadb7789e5cc3a197fe0459fc11313078af37ae395a9db9a997102e52a37be320ccf23033aaf0aca0fe6d6c35fdc77fbace83326d9af0430e95b86d744c7de00e35bdfd49c9ec14e67cb882805a1727fcc58070d5a1188cecbdce563fcd04585f218fae42e92b3c6c451c8fe9d9759af15528c7f117f0a1bb5bbeb8ffaba14c11e7dccdde22fd21ad7c2ef459e29f976d9b71b8edaf62e2b2bbb439c7599126f9561efda6cb14460fd2da83cef23c5c895eb729e5142a69660e1bd7247f3eac9e1eb1158e2d364ec1a2c4cd38a909e5999e55f217d071c01e033b46acd7e07fbd287e2b1721801b8c21b94b954981febb428e6e4875d9d719bdceb3307abdcc24bc96b0d932884950cc80fcd9096ea;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he1e7b704b7acb22bddbee574d5dbe51028c6341f474a072c1f985d5cc3c209cb6d33034415f699f3f7e4b4067162b966ab53f88ea444284274edc28fc551ed11709b2d54f67fa6ce08ff98f893f61d620b6c0ab359aed025d1c23770c66f130c957ed5b1b925a27ab09f30ba044b974ab1c9973f73827d0456afbf564bd25900fe71407bd7e4e81c2f4ed536f7cfc23e66d693f31773103822469a78d4588b06c10454e06ee6fb6abca0bbba820d85f5931830921f73ac15566b17e0519ef365384eaeacccb9698c0975f858b1ccd818ae8f63f732a27f0998e0f5b7f732b5dff6b41bdd2400f0f1b6c0a025e62b79d0415bc6b555343ebc3b26a5331e73e6d47d095f64e621f46d49b73cb83090ab97ee4d41107d7ce1cffb43c8d1bf70e494a112bbabaef625a5900794508021a00a58e2ed3ab71c463f3f1326b92df77b8af8479a5c9d12f81a81521cecae07217d30ec57a2e576038b0725c76a610dc488e9805b7447b06d7108023db0db15c1a69c3b748c7bd614861bdd5dfdd67b05832e93b074007dcc320fb1a67c4fd32c2dcac292e19eb6a8a4b96efaaccc45806aaeb82d46e14528cc0c24064a1998022c4ddb48b6499c0f52f23ee2fe92da0962c13073ee28bf32944e5901384f533bac4e8e35dfa5c5db1c2e1a4e55fe596f2558bcf683bad71b032ac7944fb5213570ebf0c08c01e78ebb0c9b347a2452edea03ae8f444f30eb6191033a3c124ce9ee570aae7d96367f430d2cca25ef5385aa9debf3611a5657cd2b213cd1a7301dcad2218d9a3d67c890393273286984407e58695a847a2c82dd3edfe14f745a8ac5958c61014b63cd7585d5e1ff451abfaf9269ccf949a03e12ab71bcb85335a782130356104ba0a07aeb1e3f7bf92b107c5e99ca30dd10559b8ff3116a1f5229ebe4a2087b23658ddbb922868575e25b215f714593badc067196800197a65028e3e85ee22e81a9c5250ada4e534cbae8058761cbbd06151dc64d1fa0e7875acbfde884031b539fb0a4029e6cde9edc1b996245782b4d53356582e5c7b6adb41a5c0e19d2584eac8c479c90fef28a6c60db9eee05cae1953ead478627a6fe8ed2e6e1fd38f354083c95ac6cb7045d0b045760f0d1a6aac39bb770e156cb36a36b8515a791e4e7d388687e3f11bbe0f7cde7675be94258c85649f7dc251cc5130b76e8e3c31ca525cdf7fb3d4739273d67897203d57e33e7a89d5560971836af50cab6c45418bbf64f0a0c18a5d58b2d192ab393644d5f8a2b52c2965f34f47014002f527a54e70d3ba1a7479a41e5a9f088f1878b0db9d6a18908cb288ca20a2db167452dfcc8f32774b1b61131c1e3ea03ffc25c27d8a76ba8deaf9591bd8b64261d6fb5c3efb9c0d18cfb9ce9ed47578c81eafe7a04e0095fddc7806853a7517b4ea5da066d8ebaec6709646e47ef32b539c68ecda13fe344a22dcd802281cb4537bdc5f5b714cf702ea54a768f295f25abc1e2ed7335f88530747008d8be39eb520b1442680d1c75de88a6abae438daa7f5d69f8a9cc482e9d891001052c1fb648606c4c064312f5553d3a67eb66deb7e2e87e81cac3a72230bcd98af64b2d333988b4267a82b21e9d8a8a112fe26abae259495f1c6bc23e9b758aa1af5da602b2d0232a46db5d99353accccf214ec4f8949a905f86ce84fe0802745e1181facd3b6f2eea7d7877f3312615f5b28b71ef3ac598f8b7d32a3153fd27009c533330166ea27d5e9d4ea4f6ffc60b8744a3f7f8299ab8c0ed22d6aa1fe445de4c2bd6343284f18fb615c990d30def562b12bba2253879cc74d91e550400f414929a4aaa1448f9375452e424e89c2c52b6b6f22c5b170d5de0f0a9fad77f3aa18590a06722c06467ed3a843474398ce55a5a83f0fd5e46914b0af8558ce3dffb836c2146a9904f5946af58007dcab143d5d2c7eac783815d82ea6866e079d029edbc55e5ef65744c9432937143834b6c91ba93fa6232029c4dd0e7c2bb7df6a1b5237e6bafc92ba59b37578fd77134645d184a3e0fe2215c08cf4cf510078759015a70e87d36fc3e8afc74346db4d488776b76d2a3a3e8b7a95712992a902c5b424d7197aed4fc5bbd1e9ed249576e4c0c2d292ae7f919c2d24fe31e93c52143f1768cca45d5402a46f7b47769b757e6fb24d8374e777d2ba68f778e9780495de20d54c9cb6b48c702ccbfe0ed20165f4fec0fb8a969613ce15dd620fdf4688a0bc79f3cf7037f487a1b4ff18c6881f31dfd060ddcdc108af3580b7e220a59211073b1a4088bf63dd9a50cb668aa57fc394edcb69669031bd247d149db669414fabb06777fc1dbd3fcdca9c758625b264ac781695e3e185a85c63f12330315c54c275624022a158a708e6002b694d50e2b4f47efb3b250d1178e82de76ae7a0d275c3b6f30f524654037e6b7a04c65686d41cf911638b4172c26ac14a8359120fbec953dfda9c5f540627ec09a08edce8730bd2a282137f018f02c851d42fa1b1b3fab01fd99485da8c51b1064d30849c937e3a9ddb3d79ebd57a66d3bd0b3592193d0d872a23138cb51efc9428fddf73b79f45cf56ee899e1528cad864bf01d08e1096600aaf7889e1171c14f4c0f79e2d77af47d9fa7b757aa60643c4606647d6890816d6be1c5978dea505d93aaf6218743a4693ed22b9364e3de8bea6dcce29d6e11e59affeb0497ac5a65efde223835ea092476d326fb5f260332cdfdd743d4c9d63f4f594acb1bfa8e69d6b103533043dd8e45a9d15baf986611a82ec81a065d15a5783045a4e8e434b31f0d804e3474b29cd4cab94c256e6604ca366296e5e9c3a1d6174b7346f465626dc208641e5300a10e4a3c2a3189010cc8cc502ae8be3042c3985e807134480583cd89436a6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5274171f7fde31999b5aecff26fcd758c2c39caa294b58645f74abbedc39a1827fdbe2765fd8437e47c2d0aa9825ed9641b9b3414f20614ebb08897a0371709a561646246aa335d22cad30cdf3fe4e80ec0406622201481721b6fd0326a44c30d55c832ed998ad63ba45d5cc6e70bfd077074ad6581af9fdae51324cf391f4a70701e2cf700e4e4038f971649d5422d8055a2ae0a105d6db01b1d99375c68ed50e99a12c91384a3d786adee13c5fceb1af5ff792c1d59132f4643134f350eb895ac10fc664b382d99441604621462925b60373cff7c6dfd59d48a3df5b603718eeb8c0574776e5479d8b859699be1b939e7d4c8e43a347e63ff576c9accfd4482123f2911cd6ee7d4dabef7545a70c1eb84ecbdeb4286d57a7387c236988907cdc8279cf4eef53bfae72ee35cc953fef4a62eb8c0727734a298df6a34d52cfe8447f90fe917c794ae309d0d4d7b2473e6e8f23d4ceadedb79b6470a1d03b48c526ff020bc836743c58e5fbf28d694d09a33f886f3632977ae443204510c619d70caff84ebbac0b2a8f0a5874bcb65dcd1ab486b2296776dd33b7125181c5692e19cd416984758f5021dfde41ff583f1b0537359cff388a8aa97112863983a5423ba59f6111f0cddcff1c25ac1c51025468a140a64e1e6539f86bd661975059413182257700dc3cf8d9da0bba3e120f07174f377aade2961f09c7ef951468a1a10741ef5a106e68561c6edebd13bbca558bd4ebddf1bfbc61be02221871d5649654c8539163eebf468c742ad8f143ed1a8aef998b79866313d457efdc58291b70e8c3a68d4c714e78ff487a468b42b35e358d8cf1ac5b7674b7b7c1c73c731c123b64525bdbd3c60de650a16ce1b6d07a62c38c1b3eafd181918a45b13556bdfcc956ed01d148bc2c16043f8e32952ad49740121d78b9b7fe04577a97719580a4f17bc30b3be93a310636e9e8d1ac3ab5801c105aa38bdbd21101b5d289d5c540e463ed9c8f93b8585d12bc1c5dca862ca8c61bbe32b818d46582859e3b2b80f3f0a446bbaaf72dce651ea98238c5b2825f71b28ae8743cb01e70458e50714cbdf049f025767210d2a4598487675d4be418d5e495d86b13b9f325aab033fdfdc7dd2405597f21606fb05ba2c060925e579944176ca4d5b4d5aaac8083d4a6d24e2229e4a8a79aab124d3f476b5527b5c6eb405224de693ced4b7dcc47ddf3bbfde877d78dd3a430f22fad6f6deb55df3d30d406f440df46457d76902d8f4a81bca33f1cbd4c02cfd009b56456b7cd7d09e99ba2ab673d4ffe55d28e47e29e346a1a6cdc913ebebdf24af24446c42abaa30e1f26df1d0a4a07eab30668a192acfdad210c9b0dc6c5f1b5c77f9fb3d6b1faed475bd4e62ed93326eadb9a909d5e3376978385486b2222a65c70e9902e7a0cb8de778db35c1947f55830ff951c1855c5c3c50890b870b62f2da565109455d1d1836eecfe35165194b2ae433724384a4f7b2724d22fd7c564e42c0b1c3365435da0e3660eabdae9225616c79c59fc2874a1c1414bd656f9b04b53cfa76c8a3a697ece78584ad80f8cb326f77907fcc51a270b3bf15201f9c52547c1583d7d99720bff74f972044f783cd359e7f7b87e6cde314270ebf01b21e5a12c39fdcb94c069cc07b7a7c8cd08f7a1ab9fcea6a701f0c8bd02a3d0113d28b2fc4e4b57019ac27123473448b9b6a09e3aa379438dc076e30fbb539a32d517df0fe370a056a5c5900dffeafa94c1df2488f40afadfc749e82c2da3fc56b9cfd6fa9921937a7eb9601ca44c11dc62f1cfacc63928978c7df6f67819cc55ceba9386cfa897dcff139468662abf769f9649f8ea30ae263ebf37fb6a7db1b1218d4baa403c966eff2fe26cf011734d4f950d53c93082f45ee5740d0b214e862b1a1996a9edfc5a1cdbde6f5ef0748aea220d9019cbfa3dce2914bad56a85e12d9eee430bbd96305b42b66e41b8af1475f1f248a34277efa0ac2e5ca67c772db10e8715048a714f40ee78c22fe5633da7c5dc83ea6f2e2e6a7ebb7a3e21ff5c7a66f625f17af0d682fa242dc93b548bd2f70d4d9cb023d0492e7c392ec9a92514271974756c563023d840fca73e01056c370fc6e46cff85d702d0108388f90c2ae465ad4643b83de4abbb2d4f009f3fcc1c3934886978b2a84382d858a012d20e152d97bdbd0db6e512bbeee7e39120a67e0b80c54330a59d9749c2217859f6ca2d5eb8cc70c694f634b7b8740efabb5419b591ff532c1b6099be4f76713565ec43a7fac950cca9462d3f5f27999f534dd1fcf17053e6a58919a596600a33faa61afd21f2669303a72aa315265adc71b1513b840222d32c971f9d561cd4d3af70df661abda94419d164c9b42c9ecd048479335a1c30b6ba51562c9eb261d25e650d7cb34145995c52d484cab8fd06455c64607d958a0a60b126aa4be87fd8f10294d9ba3c8a6d0e3e4a22d66eed10d87b79f6484339e51ee12d070ec56e71109fa292190979026fe2bab8e79cc5cf176ab20a73ad168d88c26deb666a2632fd2f98e553e81cd791f91504cbc4d993ded015090af1ca7e83867def718908f2fec7e7a7b517a5093622e23e3458d037c7116f3b53e876d88f98288b37f21c00a384ba287ac187510a49f66b308121a1cbc951b92478426af62e0a966b260af43ce2f3d499a7f24a4a6c64ee6baae02c2b81428edcb24f85ff2e61ffe0c2453196fe48f517ed781aa1c181267a7f35fcd9c07fa6b5e3a36a57d004aec98f366c235b28d2ca749653006f9a2890a2faa9d8ed0085b5e4cb8861f1fa8087510b006eff65a78eee1f5ff3aaa9188483b9546650bfada2a4c096c1735db89b57b9063c5050a4bbcbe2290b052ad730c5d0db8f1d84f8a9289d5b73;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h12b840cd2cfdf4e6148459e463d5592f49d586d02fb65aa11d0d781c51074576f1f3c857af31f59f126389b512702b0542216fc57071242c0b82ffa36c33408baa179680af74cc83c22e3639bbc6eac82909e3a2bfc93eea07ea03624cc3a2d3eb80779e864e4ccaae4fa07e915a85416e223b9642821f149427aae8645d3ef8aae583e0f75895f7c934184bc8496700d048f3cb93d30fdac7025edac91a0c35b870ee8f2d04493204b650ec57a61bc76a135f87a817e3b57c9e189343fef767a90521469334059471d1c4a1e1d8a39f9a16e720f13cd57e2b3079eb1d6dc0d411afe3b9e3a9968e7e194a2b3ffd9a19bd587e2be1278463b732cc26d84922c4f98e7a17b04b7d11efc37db9194a80bf49d6e8b93e9d226f7eb0322f57a402a7ac5e0a265207ddcfc47d4e610439c556404d130e62dfd2872b1f7a4a40d94915a619ead15519642638a6539c70a53d291dd473bc0aa1736044e693959e4b2acf78de2d7057c228b6479907f92db19a7a22545866a37dbb0fb644ac4676a50b1b4ea98087e56f85e8e72b25c5f363fd0f7b9b01609822a19b822bc0f55520d5752788b884b7b01ef10c4a220de9402d3f38e0ee6ead68e91cdd5784beecc1663251a59a3ca5fcaeefc1e03ba193de2a7f26a343c5961a6df7b2f8de5eb8b26744a1a76ab67303e20ecf38dab7372d1a1650551edc6b5c10cdde7e64ab3d283a6390e3f0a959a0569beb00c177ef87082669772c73105044d7f960701e8e8a645f2bf6857435d4f8267e021545ef058dfb521e231259fda0dcc1e1155bae7c4105c49dce61ebb6fe72ee92ec9f42464b67224ffd1eceb133409cc196a55441215269210b5b4df3bf1c0934cdd1354fd48d6fec35e1066ea3c3b22af954e087f63392261e7bca20db0e01205f71fc57c8b5e7de51fd9f8483bf8eebff0568cde400e7b845e44ee9161aa58d7b8cc5e45966cf664494770a69d3b1606822b3a847f22903b6eadc275fa8d27d796d3399e0d8e9b6e94e2e1a43c9f29d39c1f152e70ee86e08e8d1d488a3ee4e49a39433b4e4398f2071601e81f2df0302805e26e03072cc01dfa10679c7213ebc475eec6c333e5fe2ef5d0366914ffce574a8e1cc2ec34a5e1ac4a23014fc1514ba975ef5dc3f8f3dcbe7245e1dc9b77980bb261b221c8c6eb1de27ed5452982fb19e0c8e51d98723fc16ebc948d704dfdf84a352483c75286e4142f80b103e788c6f24cf2bc8ba6fdec028446046ab9f344b698e513935779bc8a11dcebd9c0880386e6dc132c8952b141ec7bc0b014543241f1e72421e1ae0e5d0b116d7dc51e7d16956009f1218014b76b37d466b3c50564184d1f598558a8b4c687bae1c896a9b10594895475ab77e8156a0233ac7f67eb5fe88656e02c3c803712866835e8cd03e104849e05bdfe20918ed204b80c9b47cbc971a68b48556a2ddbc998557e3537041f4b2641b9424f39e56c93aa008360484f5831dbc3e5d236764fc644f7c2c949d3a9754a47af412f8770b25c94d9588ca85aab6c5a8ce78ccd690bdb28b452f094b305212ec366d5eda9ea400498e0f8b2734c1d129fa0531d18f234547f97ed05e7934a6b5964e25da2f83a3419cb33bb98a1b5bf48231326ec081625d76b0fd343650dac33cb8ce121c075445b54ec6c766848a13c34efba4682f5beb53de462af61e4b1eca115d8a6f6b54068b51ac1b40700a4c3644ba65258ecbce9c29f8a0de5c090f4c8bb54c7819e1caf14933d24f1c29e0178bbbbcd78a3501e2cb44ab27744a94e2fe7810cd4ed9d39902c8bf6cfbdc04a6b9d5deeb5fc67ec5946598cd8dbbda114a9c95ca5b6aa2935bff3928c984aa2418539737ef86879fd6068448f23e6bf64c2fff65102175f479a66dd0ea8c401273ed4630e9e83838c54e821f65f494c4ca7b0c4e386325ef53113154ae36343232eda591161c7620a4ede53c3fa9eb638dc158d38d485103df7e6de874c8f0cf33435a2d1d9ea4059b4a09f32465f8f89a6fa18730c642a26d3fc1bc1fd2897c73d7db7065325984188de1571a14b9e1632da1d6cf2e261847c6b0c58908cb06a66ea696d379d706abbee30791140abafe5d3e4df9491c1996c78f60353437830236bfba02b76610b6fd047d4da129632baab850bfb1e8b470e50999abff8d5a84fd8d64d00527ea77e92601f8401751b85f74f6b0a4c1cabf1cf38b4f00495bd6d5d311e380fca25f9d9779d252d8a067c9ffa08e0b97f35d59d453c22669598f5d493106d4c2d1129c4b3985dd34d50a9fe1d210713ed3cc524ae04e9dd999c1ec70d1426c9a6c66abd677179993dde95fef8a8a7a800602fb9c36869020ea014515c54b1d4a2dc8ccfddad843b07a5b49192e8ddad9135ef93ef4450a248ca233db77e0859eb3e20e5ea5d76fc77414356858d6f19119dda04f90f30d80f31d4e5ee6f6e130e784f2420a7788bf2620de8feafc548628d8867087834f6410517f1b80746a24d3d6a912d6549b62410ee7f564607470a125b06396b6b4df4f83c83d48010700d09aa71d0a2107dd9cd0b0ef3603de3a78d839de84b49c3443f43711f8ebb0caff780eef6922e55d094b045b3a5b92036ea49dfb599be54351a4e30718300ec3c72b69e08ee508442abffd4f00c4a32b668478c766b1102f86e292ce9f53c5e0227b3d6ffe2668aaa1ecb0568f9d3935c7ff7d6c4a5af71739603c67b40d3071020f8f94e656632ba45d1959a6c78f626cbbbc6b82dc08fb5fc0d5420934a16e331c7e62543790bc1939a1edb4a6ba1913cc1abeb3385ef418ced01440a94e5e5c15a766ed6ea947a3b40c22a43d0b4260ddcf1e120519c02d0c65653d056d9738ab2dfcf6be125f2ff0eb06ab6b6d68f34dedbd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7c70dadbbec4064e971bde79586aac6f731779047eae2cac845bca5ac67733e1ea050e212e2d9d6039a76c938028f86ce8fc085b8c1d67deda78b11b8905395805726092d586748b5b1f577447994def77175c72bb40d4942eb7686904aaaf892778099ca72cfcf136cbfb08550ab7bf680290e2f81029a8972091814ef7846fceb91d86aed3f84ae3c6c86d2bf43c449250546cd0cb7e600eae5882d30d620b2ee16458f3e00d773a4a06591dc33d84a2d5dff8028553bdddbc559ffea5dee0a691d7448051772ded1570cbf86e0e3168b757337f296dc4da0e28282ae37caab4a4e7c650f8ecd7f3744c9ecf558afc096f166d1d9c380ff0c15179cf11c7aba54651151a0a0f49e1cfcb0f1b9d1fdf5f30c9a7804ef5f65642c8b8b845fbb69c88decea4d3d18f5b5134ed1b4ecbfddab4766e1fb47a9fea86e9c9102406da03e5b20a07a04500e7837f80b789293aa1da5d0396efc81d009256c2e3aa10535d10aa2ef269dbe5fa66f36f6776bda28f46ce4c199bf8e7c001ba8a6129ac0fa4f222084e5599cf1aa6de08c92365e6e8c563b2cbd47f502188188cf3de7a1a852c507c03301b4e179231e1152703cf820b131ec79fe8e0cf7b5a9882486ac4d0cb78fa18195eab959e23864841bc05a1ff821563a291a742cf3952548a2b74e46a9691f0094da4dc28ed68304a781a3a399bdfbf9d2d8ef1fdc7532c9f1f6e3fb13d61623cd39cf751440e4cd730eec4279e8c5d9babd90ef7ae7c85b9bed61c88e17b7f17aa9c7d99d2e73fb6c7397eae36f7908cea2f64c5dba44e6e752f19f30fc380ab23f26e503b7bb08bdd3b669681bb02c50b0b805a7b2d771eb7a849645b7ad468e64c71de0166bd10b3a02d3d8e813106e87407c45a36c18e8a994fc7963d62ae17d29c1958d3448ca999aa99e0d534dbe10d98ab7e1c23d8d5bee158ff08abb1bd614df712ef281595e2a74717b07d4568c7befe5237c0c5a482810a933a9941a922d6074005e96ad5134d8612b62b554c57b6867734ef117b10354ccbb5e4fca7b6d8887e046a289e4a1c48cba381ac1b914f45ebcffbc53354b27ec28ff2f7f98b283b9cf5903a08be857d407e3afc81689d1f4ee340b1b70e2567ec5101610851fcf527db5a33340843bdd544d7488233f565d9a05c479fabde38a332729a0fb6939413a5d077a08747553c037e56fa655f10bdf1b376667c583b06cdf1cf27d6563b912bc3d00f6db9bf97ce36077813d80b4bdde5b542f73626fe55f7378a5b958147b35599129867be77932034da0e2baffd4924b28644c41b3a25cf67728166309ed068bba9763e55fe37a214e7e63cceff785de7d561ed15a1b22dcec4dc7065a9618d723f15652192959c04847cc2a19a2ddd833a3603d05e0903a64bb77d8e131187c0e08d4d5de87f17aa37a33c5f68923ed45ef348d5586045f51d7671ac61611496ce87bcf00ebe025acaafa3ad344114ba9f2b65ef569ecacdd5c644903eef93dc7110f6a8ba9f9f6a5bc386a07621fec610c411d09889d17d9cf8f5f33ead75699fa7306720ac2361c99b3654e1ec4d239b865b3dd48659912d7f6f51f59a7e152c33b832beebfc2f5f7708889ceba4c49f871b519b4f0be15dd808120563f3b1952bc38a4f20be5a968012b6e07b527a170ba82d12552a95ddbcb46709b8948b2940a71e9ad6772d7d4de02d04bf6827f83ce96d951cd138d4b8ce506f80f3f4045da422752296cd23f988c6e0c1de446aec62f2820ccf10e836a24d3c12d45948eeb561d1385f1651d09e85ae68fe75506e24e1ca8f891d66bbdab9fbb001379f34c72c6b72b2d55a729dc4c065a28fe97485d4c29b345b76e208049c804d1a5df703defbc9cf72272553520b6778626af0858f92a9d52d0e18fdaa470e9a1bb2791923371f42f742876b4c5210d259fcf2cd37a54278b60c68850a5195ddf4f93bfc87970e7974d78a8121170ea5e836654583b90448f01b0ff940e83728e6ec07e6bcb8fdc7015bab85c306d85380452f603f9ea3eeeb74e070e71a419e15114fd43fa2a2507b4768f03ae23e7fde334f9b437123263e600a2857e030c7513ac2572f71eb9dab83e88f954a9780522b42f12f5aee54280821954be52aa55b0cc9ffdac0fb1e7eec2e98d5b17551bb1464063652c50d74a1292138f2fcbec815bcd531d57bcc7311cadb5cce1bf154d63e4b73a60fbf2a2c7298f15b853180486e6b04c9b5114f5f759e48e5c4db4ef39a42490db4f353708f62bb8798cd4be3dabaadac3f773cf1d4b9d61aea202ba83aad224a0b54832578455a790b7b5d55f2aa11a1c4459359b983718c7317f722dc538262e868e9bde9d3331ea0e38ae524f95326262ede986ca7a8b872325150a80fdbf771294b372db7de499406ca0a3b845310dc26f4bb51af7423ea220278d697db9a066a58cf2bcd86d0921ac15b9e7b11ffa09e1c0efc7d59030341344e0d712740d4b39d70fe170dfd905c5cd0dbaf34c83c51bd61ec3590862d5d764a30f1bd6200d2e537e3a09b725d62d84c0b383f1f3a030ee66a539c2fbba0d6c03c675633ffb0489ee971e6152128e4aa624212dd2dc4cde3c0379a8d078b86847d71dc98cbcb9e613a7ec119d58d549d09b540af3759c3a207e9a25f2a16f5c612d9beebdb15d72c1efa84d2004a617a3af54e7ef30dbf6b31de77bdace634a9ffe0d42cc3eb101ead9c8c6e5f90f4cab5d1f8085f2d0a7c1cb7653e10c55f605ca38adc99ff0c9170aa3eafdf4a93f54fb43ce09a89e337f85896e730790b8aa94a7349bb1d1be720aed19b1f67784cbd435e434379a3919a90fe50d31740256aef284c24439e4624e051a9ca9d2800258b9e14512480d373559a5cc801cb044d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdc112eae60694a123283c3d140778930f89ac35f7dfc29243d9121bd165b629145eeb3e66ee82f05bb2d72ec03f92756078c1704113ca27fd2261cfbda9c3f53920f3b8cb9511f15ddbc5784db061ce7e98a68138892b5ee60dfd5f9d39c45bfd6652fff74f70d90d7b53b8efcec83ea94a190565e27b9b131fe615efd875a6f23e0d75fd8ad29c6076892dbe84288b2665fabf2e5dbee1392c162cdd0b5a51c59635a1be4c38965b405ed96e59f7ea060388549727827b82fefa3a44e91d683f74ba19695f59b3b328ec84c3e0f313cf33bf975304166c035a2eb2f17381391f0d8e99521dff7cf0dee933b161479209d8d746447999d769fecfe52c4e50e919fc3dfbfbf7625a493609f1a112062a7148e757034c68e5b199cfc565a8a4ce33c5f0539128b1ae8ed366057c62eeb360ee49b6f579dbe34997735e5feb1ab8428b8e120747ac130fcb1e71613b4a9ef452ab273f82f24376cab0889266c85d7257993f38982f8afe5c6b5854fda86056e5e0ad7f9af257fb05212e8d9ec0b358a32572535cc90032c0d3eec131a8be690abeb49932a12413d97a190422102674d5f00781382d26091971ac2b88bcddd61022bcebea5e531ebeb00ed17e7931f61ef03cd32e55a44d8af332674bbea0a1eeaeaf111c977ee7a96a1a3b211f677cea0be1eb2ed2e3026eab27adf7eafa14d519794a724ad514149d0ddebd443c91aa2825b9a9587a5ba6d128e7d5de1ababc85cc7cfb5245d6c3415de62b465913161c2489faef1908fde659ac321b43043a01f8ec1c6b726bca608b33f87861dbe36ab6815ebc539aca1270a57862e2aabc9d72a99fd534114cc52bf3fb91c19dab153e8dfc0207aea1bfdc7a56baa7fd63df2cbfb0e3b61a3c9cad2b4cf7a8b4d363f6f227c16ecd61d0d410c7163141c3f55d447854a96639da6c897841901cb75e2bbf7b6515d86b894909f465fcad3e1c25a3867dfb86ec6d68109fef428ad348e4b2a8a9b3867d0a4aeda4aba2d3d077f103815390445b04c399aac3955b3457270a8e4ed3836a0770f3242d27b05bf81ad395b5b3b3acdb721d5a6e49874860e2025c77715106a14bf8bfa3b5a38f3aced81f1e8393bfc81c50478899187f8572485516cdabfaf2cca869b80f9c5d3c0ea901f8842f0705d92ed64da87ea253bb186ee4532d704587d0de08be97a850c90d57ab837083e8bde1446b4e545511f5587208377f8d4a6780665037fc0421472d3862765873dbd95a788ec4222934c7cfd1ec3460a7155ad832991c6a2c7dfc486ee49cc093cc1e62e6ea0939db2d141392673f33b82fb6717e0b00c33619a32c74c2d7f4ab6dfc0119678ab6ffb24b934d7aa84c09192a06340de2165343b67623334790832e66579b53de1ce0a33cc434ff607ebcaa639235ef8f3e0118937b95f63f68b5140a527b5fd698b83c7f343edffa55b4bd492e8df9f63c9f32f494f0b9b2207faa4a13c48da352e9f97fd8b5570a692bec33b38b1f092d4172c07c630bb59e59ecbd9258e9445077137755565acb4be41f0d27da59c690bf94f3f63b70a026a2371377239126450c2421e812fc7c8498e1a3ea6db5cf5d96b43437916a145e24f2551b8a22184dca4b572a2590f47d7f5c34ed3848d9b924472b22660218a7e8f0ffcafde5acf281e03b0f4354589baf0bdadb20c69ed8dbf4c2225b2c5afb55163e2a0682a700251cdaf53ef6ba3a472f08f8239a27db9922ea3c141dfcbf7fcb21b43005f8b784a6f0d5034176ec7dffb866ed171a27d9ab9ade8253dbd523339323c5d4b81e3d8b8d9e1d0b131dc92eb215c30225a61595e5a7cda859a2ba1f5c0a8fd8e261685acf20f5042df77cc61985033f788a4a4e7c179b0186bf5b0f59103074efd3510a7508961244fb6050bc2b4befd2ffc5015f7bc6f2c608fcd637977e92e54f46e84793f8af2fdbdf8f529cee1a151cf7e42f16695906b1a3e2bf552d572710b062d6980831739756cb93db62e56635f25878655f130e08b1b76c025f733578a174eb03f263eb393331692f534e3daba87aca2433a063baa84fd80f7af9e646acaf5994a676b1fbe652da87dc03f30007485ba0e99d1191c150cccc49b9ef4fbc4161aea6fd477344c8516bb88b371923b3d58ed16109ee1b52d5e3c48ce9d1d377436e608bc91b0677805054056e8ea09deddb6b2b7d55c438d7c63bcdf5af0b56b3aed5510be42e98a29b4d722d4415361dbf621100044e747b9b04ac85a3df8f5706206a1699d8d511e54f235c448d99c5a852ed1367df643ca29eb1fc262d1c86d0f6c050146b3674ea3d6690c5160ed83680becf2f04b7d46bc0bad6637a021bf8ac75a724bd2b78d8abcc8fdd4464dba083754baed18f007c2a6a3e195ad303cc0147beb81a9554c3b37acaa6581da88acb6425338e977542a2321026b1942ceef61a90aa28db5d6c823b41f3fbd87eba182971265210d99e950ce488c4f7378d6fa03679b909a3f6712b5252196faa3fecbac8b0201ba21031720a2dd929c4864b621725918e3f19028dd7ee04b5e8f8258d012d7538d9b155712dd78f657ff3282886b83deadd40ec6c0ebe1cf0c3e1394eeb090f9d1912f9f0455687d613439d051e27e525ed23ac5e13356da4a5ac9e04113bb8e4d844d6084a8a4d321a4a0732b58485f3e1f775bb8d7f4ae045f9fed4a75031061914d6fe7a40e877da78b6c05bbfd18cbeeda8713aa9e3f5156db0575f9a4a81c0ed2f8a94c1b8456c556e93ce40ae6fa8d157edfb5b57c3acd0fe360216af08bd6fe76e482245a8fab42b271caa7c7322607101456b594550c8df9a9e49e6e82d61e0cbf07210a4d266d7cb6f9ea0ece6e9661e54190f40f039a7049b80763083f450f9e8b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3557dc4a20936f88abec774ff365e16ac3cd7d83e4e7aac049446bd9ae5c786f724fdde4a1ac1878f8e24917514e7863bb187c1c886d388fd7e46b80d8adb68f4c34b82a6c3e5f7c167288376f917182b206f3c11c0eccc813d92262a52694425ead19a6cf4e29edae0d4f632e0492b9c7be365cc77a6422b13b2add4e7b634b9c8153a9e6919d3de99f81275a41392d84e0c1695d48cdb2c3a5773fa24af9a2dfcfec925cb6328deb1abe5ad127c2fc7399cd0b2e5520c608aedc9d789da4520ce3630d9530f2881e6dfe80b2f6a4d2d16073dca4b94e9da68b850bcf69c904233f8c904cae6e0fa91eb806caab1d168d72908fbbaaa75f94cdd8a27d21eb6faeb813991ad735b0866d79e3a1afadc481cb8ed738c33a130728999f1cea16310521cb7f3f29037f04c406207fb32b0edbfbf454f6680a27ae3afc32822982e692ac72c071c5cbfb9b675fe8b3cca432031262a982ca8baad77d80cb78f1814bbbd6d7a7cb04e9748dea742308e3832c816ebf59e1603e48de8ded0bb7e201b29b6e5d10af47db3959d0785bdd518c11ebd6070e1b471866265494044047f61e66303d2ea5483b131d202b1f04035c71c2e2830d58586a53ceb4ae502d23baa7b1a260b3fc2031cd70febdb6c1f2d8d81fce66d1229639cd0cc912a9d8a438b4a796de44b8fb190b3a02565348c81346d78344f0f73fc7a9e4f9477dab6fa88bbd262cd7bbd37f487d8c3c001a7ec5df55f56f496c8477707258e846bb8d9d472c943a20dca6971a93601397fcd586a28357a050552af988bfaad10eca3014efb7a2245545fc8bca18d2ee7428539dbac996215fe2ceb536dc9673754c9adf04d094c97143db5c43d0388618fd1eb05e255b67404895306941075b2f7914cf12843fff218828868e7b45f163cd26a1a4dbe56bdcb7e3b139d5505d49202cd08039a603bdfd1bd9926e7b5bc3bf95df4df99e2766c350228b2e9f95abfcbbf028faffb6a4c626e79cc26c02be36f855105e7285fa66ade3198e5673edc878f2692e78538120ab099774fdcfc9f93d0b2170894dd995987d2b28b9b0170653d64199f4ea114e7d6586ddfd97b660f95de152cb792ae963e026165f32308af1519c7658f256ad512159eacb859ec7651c7ae9ad8f10accbec7a546d5b8d5e2babac338ab7370934a58e1131e4d19e4596f2c9eae2589b4327a29759b849607c26cccac2b955810b78a6b6ce514aba3d15431acb2ed199ac1ea09ff90d383900dfb6396b63ebfa67879beeb9040d61e2a4e526b19cf3417b78f8cebd8d6bf39c4718640b38691e44ad35199d8951db783ce38d6d37b82eed57cf70c724cd7760b7ab3a3545a6395ca24e63b42b4c01569fbc36cb385f83eff3e9cffbc9188fb092af8938feb28a3012424f579c4f4c46dbfcff9c830e71839b8807a81a668cd03ef105697f93813fada6956d63e542b1c62140cd0d54a905ca339e5cd8cbef6d8052fbf67c715ed00fc73c7efc79e588a8c57b07ef5a765b7aa8d9bfab9f42a387ec485191959c894b360a7507f02fa84786fbf32ee48ca311eb01096e9dea15d0e2550e17bd6668089e92ec0e1edd8a45ea53564f817b4aa86979d62b91674bbd1e475855e7e175161d2e1d8a7939651cf6d9cd4b9df99e751c39a972c1c24d941b53216b7432b8cdda156f3ad95af687608b005c0a4954b254cae1059a33472fa137934dec8daad17e350d7cd9db030dabf08adf10b82bebb261bc369cf3118af29a1b3d05f31799b04fbd8cb3d546c71e0b7b9cec99727ee8c0b7a33701b6a3f6b94f586581a1678f7d56d47d5e373d012fb0fe6b88c68082fe0163882d7b6d7b1ab95811669df427e8df37852036e94eccfe048414055b5f1ade0759df242c531013c0b242c252b509c60e1503c543ce3573dc00108ce68fe3df8e137cf2b9c60e23ab663a0799e0a783fbcf8718fff3d06e16aa53edcb373fbd5cc6e49373371edada2af019b1b0f5654d16e3d6249d70f34267853d39069706ac5053334bf3bfa7e9c90a82efe561acf5bcc5ba9f56a2daad0a7fa43901ccff4cc27e70c1bc31a344f11f499826a22de078320e884667b08d521968ad1ae8da0fb7501423569d93f802b16f5e98768d2df1a294f29e7f965003f206817337f0171cbf1682505a82e63337595ff0ff9c6bd304aa5e92829b56788b428b3f429f07fcefb7d9e9ec192647ef96a558c91e7a7b1edf2735dc7d6e3e7d5ca8d494da669f94ce0d5c34fdd5012dae4bab540d10ccd9b5955e6cc4a3f25cd585b4bd676516d44385a616962a6382347324040ed1fd657d29e6e1479839ec8a75860d04ab6dddc54b4230cf2f49dded4ba4a7c75dcc2ca498d7f9968480422cef56aa9084d7b52c68da32330b4b12772299500fd42e1f2203b3b493704cb92bcc297eb89e353a73b7d690fc53fc7d60126ba593aed1626458130277209575ac9421a9097b8a34009260911e6a1e5e7bfd4ee615b64959b7ff550941acf81ff2db6c5cd56cbcdcf8cce127ab74aa46a1641abb1e08bb3133cd8a10e4c26cc1898a82770707978674c26aca943203f7ff8e8a5777935fb5858ccf4ac94841d148bf55fa5a2fe4a269b1db3e02578907369d6f797101482e73dfc3811f0e3cdd857b14961c90eba38b83f5ff52a932148fd36b8e756510d86c41644501b41b16d311747519919637c83db4b5d9155ca58c0667b1e82785db9c9eb740210de6b67da13d23fed678caeb8285397a3b4507b020eaa97c754972495ef30d43b84ac2fecf6c3ba38470098d43f3a64e91ed2b556e4e7d591c762148b8c3cb63aa8248bd0776c6478efdddc25d2f7d2f6a545bf76a84fbf2a5e76384ce29f4ab02b4256438fe8c4a9cafb164be84;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h75f3b988bdc6554f94408961c1bca8bd68564872cc1255b1bce901a43473fa811b45a31a82bd23fb30f6a4620abfbf0257981d1db8c60d47a3073b4cc7b360b5c9757e4b4a68c20d6bd0e8a3e185a3ea029bc747f80125cc6e231846765e3a42601ea80754ae2156fd4fb685ab961e7a7da44a66a19b50522a86a80f9d3933317d04591e41cd8b72a788eb1e38ab6fd75c48e9966046333d4f4eeb01fd2fa00af3085707a4570eaa04a7e98f55c98952039843fa1152b642599a8f02802f4dc22a7f4392cc168d45f183188d29540a882460c50c660b9b72d353a9d01406d785579d7520878f761a3c0e2ef52a1d7c895dc48dafec798f350fe945fd81b108166b98815dd0865a77853b831bbf81126e5a22d92b4a3eb8b8724967b804e048e331c7769cbdbd3f9d0125c6ccc345dba83a4156ad9520bbe41d56fd1dee208afccba089a80043aaa08cf936fb90c8d1f26c0b560baba8c218b007cfcea7279de5b17c96167689830a5376b2f5383039819bd50b015a1e57d9fafb5eb3da2788e708f85c3b0f110001a369f9f1c1323ca60ab0da9e190695f8ec817bd740c2ba6455105816d3f6bffa9f08ea6fe13cb9370733b243ec89573c705d4bc4abb626c357ebe35e6cb2d6405cd6e4a272f61eccad9006730639f9a2fd11aff81e6ee8fe3a52921af99781aee46911ea4d0a612a9128d694cc510264d87f1acc7af3b719962993fdf93b4e4849a2ad4f54201fd91c016ab75a847ff202e2e64fe445f4989da4eff81de84cca9da4c79bfaa7fb7e44177aa4c2f268c645bf72e44c67448e083d985686f0de9ec8ad4bdb329f6ec210807197237e3e0eb22b3540af26646f2710c11a0f476ce4b99c01174e39f4ecaf060d6a809cff0c1b2d009b1f3b63a203a93a5351fa389693683377c68f767f51881cd65fd0928b65dac468f7d183e31de42b5374047aeb468d7d792254b0547cd23ae17731e7cbd791b03b3c125d28704a54339e676c5500354cf0fafb2c4c9e5139bd5cbfb8fea0de88f1d5b0cd70dd9ee8212e04cb527133c4c07478c0bfabc51a262cc1880284080a16c086f6dde19b588bc6e7b046e273816adf18f864a213b12c9ed5d9866bf80879fdc7198454d65727b6a61985ed401fe01991847c7a39edd60cc1a02ea17cc648eb5999b75e1b5dad7199bd82dd7bcca7b82d69ad8ba11db22c0e25f7e76f88291d28ed9ae712311bfb5b91a92adc477ad28506161a16cdd9215ec4c99b658b2f6af8bb06edf5cbad3b8125fba7aed372d21cd5c6160bed3c7fca0c0e7b7feb568511c815b04235f62826e8918daf1fe0a6b4bf5b5a56c2e8ff1eca07150371b74912a97d33613aa47ce4b75a8be21127740a2c22fe90331e020aa5be779a1dd30f9b5cd682fc1c9d48da925ee2e77225848118c29d07d3705eb6982a933f3f348bf9d50710861dec7c991cb6fbf6e8756a2feaff3fd83cdcdfb2725a64f5a1c4cea4d334a0660090763eeea4de7ee179d9cb3fc6e047319cc9eca9436d6d2d61d07f70bdead3d699273cde7fde1fd43f34f50a5d736d98db5b7a9536de61c230a5e0396f6d6290c791f0dcf13e17d8ce01fd6cf1780c5573ab11d5b07a59fe9d1238686acaf7a67940f49c3c8127a677fdea057c5b73af932121e0bab82bad95bcf39508b96b01e2ded43fa07fa67f42934c4020a8f14e59ea736d27fbdb66a76f7108469a7af383fe46909a46125fbe7352da7e2fbe2c5159740576015732fc02b6e02747bc2e37f2c5ff34986ddcf56153694d3d4ef26c9fdf0796bb34fa19e661200115649114d7be10dd9da8f2fdb9dda36c965ab5c4b57b3eb1b46fa02088fae05da709aca00cd377aa7cf0d7b926ea48da565975b3da50fe2d4f001913f08fbbe06da4bb51f22f71aa472f2ae1c5f7a55f5ed7adbc97cfbb6789a14e6918a44b2091a0bc2dce78d41f7fb1e11178b289590b35eeda1729068923dead640962434a21c5a33d1e361117f613a5b32246095abf6ff7778a19b3e8ecb11b7666bd3374743b4464812092c2957ac108fab792bc574bee94678f9d5c7420611aa7f9d716e4db1f29cb71d37bd8c361d9152258f612304a7f3b6ffa6c3052bde150f0341341823aa56b1ae9f174aaaf29ea6ed45744cd50b818dfbf85a32ce04ce6f1de60e677d5d0066e544ac91408a8bcdfe514e603c39f2476829f3e2915a4b561c9534ebe686a68abe3fa79c99a35b0150eaa483fa29dc062099ec0d8ee981ca5a59ab619e8adc578746c43f86c4522f5015f4796a292dd59a6168d494266d7786440280feff34c13ba1c04abc98b2aedb3df25624b268691622848f80ee332b12a67d0f84a8ca314283f86cedbf708a32d6896967c4399ece077743ab9d785bf965dd98b6163c0e85f91f39f194ced086b6b62c5df7812cbc3ce3dcc9eb39c96dab5a710db08284ec842793308ddafff4227388d8edecd03665fe3e79fda768474ee60ad2d6e1ba002bc30b1d3462dc0c5b9b807975119fee36a1d413ec1cb4a988e012c0fec323bd41996cf07db300cd1c7da5e28ae325171828ac9d69a02d4ef7d9eb30ec1b9fa0f7c335d87fc245354a848b5a99f4d9388feba546284aba47c39092645a75c41ad86bfb27489eeef28802d59b6bbbf4665c3abfdb915022f9048e7bc5c63fe288310040b004056a069eff8fa71388e6037deb241df66f66df08fb3fc943da12c7f094030b13cb6bcd705c5f57c980421b325e998c8c7e49d983810039456877f523ae33f0d9015af83b08be00885c37c5b1d4a9964febb36736eccd06745ea808942b56faaadc699c821c7d1dbe43fae532263f07bfe2fe275939cbbe6bf3361bc9d918b5252f5a9bc7b4f010ebf14564a270df4eb11624e16b3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he16358cba851e30cb342f5479d2be3d20be4911b0ec6fb280a560a8784f541cead44c07521f844f214f02a8f85b59ad71cab881a29d324dee96b528181fcd302062a6d8273bdae71d02559dd12680fa64166ad5a9963c0952f0d83b25cb016f759eff8439b349df034d0006a960b33fe62142eab21cfff7e345b6021df37660f86f8272714ff2cbf6f936e18a32ff7217b72a1b0bd8d5203aa9af55e0402fd8f872ff96a47fd1d1233b20532b6d244d2e47e54ce8b10473bd4fa19fcdbae4acaa33bb31e328274be1114d1e58131c18ae941af63cf041f11a11e46db61354b21fbb656f742359b8211db3091125217dc6ebb4b77cbd0413bf0f1eb94985ef7af66e053728af31ea932d40b0929e35f2e9d14078f575120a1f3c3be0f3ac20b1bd94031009627a31ac84d0d92b4d0fc7de884327fccadfcc203ad402791857d40dafc4104bfaecb30dc6eab11f29f91a28c8fd423dc10f7afa13e2f1d24ed442df297e64eea781956510a25e0d93305e86316d66bdf9208f49446f388b5cc0f9e1b83ff26a6eff7915e2610b80701cb8013af98ee0d4c4fbe84c9e61128f05df1c0ec317e4cbda95f1d2cd94099884db8c719efeae02250f6d4759009d5f5f4b55124d449e84bc7b743f511f3e62d5e14d52e35fce87ce91d2120753426560a438f6b7d746c04a5f250ed8aec5194be82a733a51b5210c2623e6eaf4a2e5794a19ba206e65a24088d3361f329d7ff711cba43868d2e062ce1f0ac252e7781dcccf3a5209bf95f22ef0d07ab47535444eb7bee2fa6d0a641e6a4717c47ee3f1c648880b58732448133fe4456871952732eec44cbe2cd00014202a7d37e6e9a71eb65fbade77e6930bf11ad79ac58e8711412acc5b520fc4aabd3444ee5f704f21732e429ec243c7d52751fd54675cb73b9041029fba7da4eea1c9943abaddf0584f1302be4e2a9f5aa1fbf7a4f48d76ae81933ee153815d22a6bd4bb65b93a5161f0cbdf402592cccc9f9dfdc3ba48c6d23af9cad9f90c140756ea1fe232f8080f75ca3ada91fcf89c2916412f2498b30312e93f3a94ed171c70f3bc1954e6e9cb9a3db7901f29b534726cbb494f9e4a951a36044a60f2bd62371cd3074fa24028035e88e811b2c303a08f42a3b04c34aef57e3ba80e2287b6d4102d4bd903d06696e26fae77fe2051659a0ba822c2c9a19eae2672a759838be3636b3801b4818eebddeff39a7d03535453d279009c44c64a262311433a031ae5e236c8f608ad4f29e77c63b7ee2b9bb5731968dcae7dd800d613f3c2363b48af5e05b0e6cd43136e21de6933c977ab2745497dfe46e4a2f0fbab09b195b958302beddcd33ec6ce9cc628af9c25d6746b47f85d2afbe41fa547065da5d377127224ae368c44a84152ca361eb2e58a9a87b4605fb6dc787d58040bb8c68389bf514e9ebe971d8a5933414cf602754573f0985d594edfe42b3dae1da920bb84be8d2dcbb03b0a7156cbd412aecca79bca28862ccfa6c80d7672855e1f6e7543ac63697e2fa421da28d874f8d35d912033288a7156e3a134102c8ed80b36719c6953e10e03fd4b3dbe7e7930e91eed407db7a041fb2bac49fe1e35a300c0631a6a30af815f089bd01258f029d392a261e3f8ad3350f265e17cc16b2c5931e4d2dc25ec5d822eae451662d09838166ef579da8465eb8af6440e9a570c41a4eefdd02886afc1929ee1bf4183f919a9b53243491e13368b68d0a2a9f74591ad121e78c3bed59ce0f6bb0f96deea4d84a582afdb7e7d593d950844efa14353422ad1e8cae1120a9d82d7969476df011e6e7caeb25e4f3cfdc5413523737f0665e9939e7543ababcd840ed88aac715c5bc8cfb5ac4056a79687809d4327ebd14ad5085868450efd6d4cb2d9d205c8e4dc5e77e4ae027cce465eafa53623ccf16403d46615bb93bc77f8b10ccccd3598e0e29c9bf00e4b2bf4db0c555da229739fa01905319c26854291d7bf24807c7459e8e1d54acf522e13d68340d41b1ade034bac544568ec01a0c81949fa8b4952df9a043e1d21d9fab462c979b19b060f5233aa1b540ec84063a57cb3a79cb8594fc145ba4f30e76d0666924abc33d05b3333ed35a9bd6f940737ba7a29a2dd505c9440aedf39c7911487718453264ee288344bcea3888bd0665a8a7b91315a4bc6cc8e01a6d4e7ff66897e235debe9f6f04afe0cbdc6932bbb044eabbc3746e8cc9060e0a9fa3d79e700bcbc6404f9ca4fc16e5f9a342356424fb6e6dd17a9e4d75338b5e51a319a468f2214adade1b1f1771d1bf497666cba872459da3a0049773f6fb9232ec483581ab5a1902a28f3a1824d9fe77277fa23c20be530a8c5fd268a22f568bcd48956c9c98c89e57dca1cf4af2133d8b7881776f9ceca93dc2fe0a94dfc5748274775c2d112e2be7a4cb06f2d7706a86cdc949c326e97077d339dc7f928c77c7f89f8e2fe0da4e8dc18311165ece6d1a6bcf22f1259b05ef14e0c3dd90fce77b700388ba43252e068856bb747b19f18fce8a54d7dc986409fbdc6cfa7514b3eea1e6b96a81fb061b959cf8d5bcb1533816fb21c3f1d0fb21ff121100e2e152240ebb7f37e5dca910f39a0ae15e51df53a87b3a38ca89dee51f5afde19eac865e430da72fa42c4d771088a8e44894b8306c51db1c9bb2287d3ab0487a381e22122ef27deaff6ae42d957f9e45eb7578beca468dbb56d7166560e9f180108f21f5c866e98b440fd1c68941f20d078eba9a12cd6e00187cccdfcfc73dc1afc85f77c3b4fefe3537f8e8ed7e77bce5bd13fd1993ebfe199f256f78bc9e061c1fe0fa9b3312e724f9de496c0e085517aa1bd8f7663b81ab956639cf5bc07ed35f53dcfab99b958c78d35b64ecadbe74eb87fe5e27ca84844;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he05a78b5d57371e0471c7064dcda4f7242c2e039ee13173d2b528adbea93c5800afc0aa98abb9dc8552cfde94f372e5b2ff30fa00f5190f9c5001d32e9d94af72a26f570e07eec564b9ef4e96d7e3685cde657110faf8dda10715acfa5b924eb47dcf8dd8aa78efc4b2eed430f7d7aa331fa500dc53abf18beb3ef6facf9794b7bad73a699b676c9853974d2dc20da862dd94919a8dd662fb626b802a03b4118f5298cc22e293de6a6152085f8a9c96ce3ff84957f4ff44533ad1329e608d739c1763178158c77d1243fec3e16025485f37ddf295eb2e260fb2d9439b8a61bd0ab9d952865f848d506c9465a73168021e2d31512ea5628fd4b4e71d32e7b00a980716601e285685884b1ebb2c7b12b55e546ff326f75b1c60f21656c3efbb26909c3f286e36cb853a667797f736bd4e1688328101dd0067f20ab22e6433df30bc9d4af833bb967cd483f0e6371d4f40cbbe1a35d53bf9af3ffae48ef4a710e5780c826c3eba044dbbf5e953fe50450fc3bf1d7506d8c19308b6ab67e1dad00859bb072499b0d1de69df2d402bc721cbf7b44ffb1fc2c1a2cb66937648b63d8e24309b64ae6546c94bbbbba567738736dedadac6f23d0243854ff65279be836c1bfee1a0c2b4535f73754dbad9f6764c50e0058e1fd853e1842e9884816edea9e514f6c14393b76396ea209b17de3d23132d6143683c4c92eba4803f767a51df9a9f81881a7716b0b4e78db7da27800f41539aec63b6f0d567cc7cb70416c335172cf3c1614ce6c8f8b54147ce629cdaca4ed8def622cee21a921d2d2d20f330c3dfb32bdfa5aa19483d93994e5a8ff0a379d083d307d556873637e8c17fdea5f9dbdf81006fbac5f808953b9965379e6219cb94fdfe14699a676a9ff65950bca6124ab899193f56c44d7269f9d2cc79117dea6ce3c28364d1e7283247501b7ca9011424a686a7e4222266532c9b78e7d9ce1940b2e28159d04b8bdedf0871057a8ab6dc233523fe90ac9ee0adcb2f548db11b7abea9a594e0e1ae4a8a79cb17920196e804f3d200dda47bbfde4b56f1b8e8457cee7739764fd051b1a26db77a7f4cbfcf2643bec3278e4c54a49a5f54b7feac9d9801cce12dfeab548084a33d044f6553d273f329f8f7a1e8b9a06466ff461d1bdc31c1c02f799de96927a6d74cd67a6dd669bac21ddfbd9c5b63886538f920dc6d276485af3c7a3abbb0d888d6347f85e7eebc3c254794720297dc852088e623539175f390666048fb6f764b5795255f0175a2498a532da9ae709e14b2c6e488d61ba85374ab904f83f28d504b8353f05863e70d8879688e07c9ef0412897695f4af56968594538043848c5597354ba19680da327ee45a7b76e58ea0ba1fcf95e200d2ff82064a2ed4f4e405e9f57a89e8eca86f7babcded5b723156e95eddbfbb3e37dc06cda91c673bde7306a243803840816734ebbb2fe6666a0fec55f0f61d17f5dc5d75d42a9ca33c7b72b70b32533e9ee680de100bf8b3aa5a9b34892a073665c7e2220b604573b5c3154e5b12877bc430ed45d7de456183d47870ebf803bb96385183dd5bba07e6b31287eb1133c9d59b47256e5aaefa448abcca0ec78e02a24dffe7a702a030bd81d76c628e1173ad35c06897bcf61c029cdda52883c4a9277bb14286eaa6fad43ad014247d394a6d5901380a76e2dc4a096bb3f9df51c5709deaee8a6af456987fd7b266663a85ee821a3e5de0c4ecd2c1c859f6481341e198c766901d0c3796f708012e1c1075accf43d142f54cab3ae398363bb3c180361beac48db682453face5a63093f1d8713b464a27f7a8a6305eb1ddb894e7a8e677979febc2c1403dc3437a51009e0313276ebf6c06e84552b9628e567e6791c43b75cbac1c3ae1620dec7a7e1ea52c9388db0b5054190711788939b9ad119110f48719d1164f75b29da7c07fea9d197ff326c8ed2da2d4bc0d02d6de50fb75af1736b72b6052103702198a1044a63c265cca14b3a6c113b382c0daed262f5aced6b995f7d6597dd221e4120530532ad0285b032da5f5090877916ce7e2febd8d5b5a2612aeb7c0ce61e03dea246aa07cb526727ea99ea008b8ec58b3437523319567f1d7e1641bad77d1431fbf6943026bc422f02389d7fdf1d963438ec9efc9fb0ecaf9a10f3d1092c8ed7d3b3bc7f9c4bcb5c8fd783626ed4fb069819b10a4f0e9383f37d77055653fbb6cca19306697d1402ee0ea0d62434ed8a4921c564f45efe7a5b59666d08f3f8f385ebbb151d559266de98d34d76df7702040dbf59accd416e9f4bb9255dec9899197aa2ad609f72af63d9bd35ad8869b5ee0f5e151c00e242500b30f131959a98a616d3974146f4811490a56c9b6b357e682f62e268218b4ebba03eb161ab411f5f03a17d8699ef52f0cc884f430e3e113c111659557bd62b3c67607f2f8dd564e8bbcb5474ed92cce7f0019afb07f411c47a8a414df1c412f22fa68bdaba76aa4809237531d1ce86c65c933242cc7cca8c98b46d55fac1e182c79829b227700666d43a696d9580ee086f4ae8d06b7041457933f26c28264559ae85fa0fbc9bb72e65c013acc7546aec5915baf6e95f6814545646794a59dee8bbda9e84a695021389ec4b658d353dda638d70df37ad8e08962876dff3696cc89c57a5219f5cc45381fbf56905a9854d7e11f3b8c64a888fdee86d6077c101933f7fadb58b9c7e86d120b16efcf02fc4a73098ea38ea4dc7f6d7921866071d3ceea6198d0053ddcd029cf2d16f0c4d2a1b483ff0f099abd1d64fc80aff1a7b44c038d7deb321f5915b0c63f28489a9fddd33c17fc5882c6ec8d6cf79dc11769a81e264ab97eb12ed2cd83d2283b35fec8a893a0da53cba2e3ba64a9cd32f3ec871596f0e0e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h62669112d5b3c25a142e0c4faa600bdc25120d540a4053129ec5b6935b443e889f36e081bac9d7d6817d6d3167f5b0b30aee65814534fb626ce3cc2c6a3e5ce7bc716950a3a14c6de3ba09c2a802ca79293aed8555bd8660a377902b411476668511a4884a31c7dd6f32f6eff838eae97e1776a36f1f1fc73b310c188a9a599d22012dd22301ca0bfd87305a14e7c9b0c51f40df0b38ed76566fa37692ddb369ca41f40d2a60370330fbf4e390e11fd79b3173674a9c8d9c5354b50004a933c552eb6cf1ba581e835cfe7d0c96feccc95b348ad5a20c2166b80f91276b484007d2fde3740f063459504ffe1c0ecdb923e3476d28cadc3a95fbfdeb7f13667cd93d1db28c42cff927866e9f9850a939d26fee70fc46447b57b35dad49c553e4a9655b90825c07540bfd0adb18c4d430fbb91d6530d11df2143ad1f8489095190700c7663c8909a4bdb1e3bc467fc18bb7489329fce4fd193dc1946d637a579880dd4c2609463b1a63edd17304a91ceb4d757d0c7059ee555ebce81538d76c6c76455197633a18f5df89226d8cafb02bfb1bf8f065545efd3ea60b03baf917dab5774d10fbc1112da12c179ea973df598e90731f462ca3c5f5eed6fd09581e1d5385e36fe288f31bbbe27fa08b9197d1e1fd7c8fde097748e3cc0c078c8eff23513d111ada21652f3add16d99346992392993ec76f7f3a9420be95408f694c4d9465a2009cd5c3eb65be6926137e3e4dd15d04c795158b273f369b840d6a8e00b973a445642eaaf6ebdda26e7b1052feba7350b15a8a949216658fc48e9dade3a1990bbcd109b0fe4e996f3d9c866dd821e61506cac45eb2857292201a7f2d33c5d9a6115597a7a83eb63cb0391022afab687c408250eb61e5e739e964eabdae4c931b48a71606050021030bf6e57cf4641fb320635ea8c612b09642023a14aa76765b99c097b2666f6cd8900a7cd8e2a2dd8de7babc26794677d91b6bc1a7963256e8a9bbe76a30f36d369a5ec124009d698046518bac21e9bd02c83e64b3e87784b32c4bd1b4f5396a2d859b20bc3e050be1d90aed9a4a95ff8a27b0db4bad11086a41e6b0cf452faec62505c64707daf73fb5c7fccd7bc78462582f4949c24f9fe56a271f8c54093b591292855026e174ab15268b3bc2d64f19cc505273900c6dcd6257b540e01ee342694a3ab96ef3b45a7897985936226c7726b291732d291c67e4ca1b9527377259d00ab0bc10f5f572a03810de24a317ce6ded3f2b1bebe29bcc408819c241e84201cd9b6112c78a6ce0a4c32a44aaab7bc1ae3d34a8484d11e40b41fad326e43e7427b3f7c099ecc5c0f2664db226870d44a72d20cb1bfc6eed260cff08f24ce01d65a34cc41160ac611ed875b337ba61dc710a9536e6349d3a8948422da1ae044991e19bb626cc4f91a6e1cb1f1e0e73f2ca17ee62449f66058476935ef7a6a184fe56739a29eac25febe2b7d90a20943e91c22e0f245a266a59016d8171716f321f29efecd6ed2516221179ae08325bbc219867e0abe9cdd43b64d062b1e3915679596371c66d8c3e931e5034420ddd10e20bed05e7064c93f798a0ba93852cb6d81630edc19bd61e46d9edf029a98f2a7f6236b52f53d72601323e24e11b3c1cb083dffbcc084a8855b53b845a27ec903074ca528874845eedc649f1819c3bb3cf098ee3a9de25a116f50225405d91925f335f9710cc55679de8f9cc94bacb93066e0f9cd0dde023f06969aacdeb438d24e9401a85fa17b88971f489f02b4fb3f11c2a1533aa653839b672ae999e938e362d1545c0a115f7f637af49e018c36513ad4504151c836003c8ed011726a8ceb07e0b55a2fc07a81153ba8e2f5256752f3be535b9d2311975acd3ad306b3d1d3965a01221953e358215c1c2a804942c0daec00d40324babd63c3b9a39b4611496c13933f15890483897903f4e7840f1efc1813e6e2ba88c10a3aec795b0c8c49eed876d59f6df4506bf0d0d74b42a742a0eb62e07fbe27e71daeb7de3721fd42d91436c8f6223561f9c5327880014754d129f0b0f6c676553d866a232e12fa8373f2e951a6041c2248842331f2a246e214f40a4de05bc85c3c249e1c35b5c4402b87ffcb737ef0857f7e0b5fc2c6da587fd18a6fe20677d6712daf6e367ec40ba487bbca51c0ef6be4799f039f019b7d5393301f4f326863b5f4901819dcd264963d1a897acb1332bbd7324846b0a8dbfeadf0fc971bd9f95b6c2f60c19a8df44a54313ef8cfb60f6bc392fac462ae139d5e7d67779ab9ebe86ff1f753d3fc7802e63f0a96911bf0e13526aaf1808189d791e1cd9d1452c075da60b77306b5770e834d0804a758e19fdf172dbe21396f95460b23f657713c47f142e435b6e6cdf685d17ddc28d2c314bcbdb1c0ab16d2a1ec4df8a436acef8005120e34bbfbf0f12ef6bd36955a61aea3d385ff603ed4fba1429a36943b5e8e760d9931e0d722106b8e75447f59aff8a4e316ae757f6cfa082f6764dd4940bcb954f719bf869f6da158428d4d7e925be2f4c702b8e5eba387b38e7fa4e55e52b74f81b7b4a321353ca04544a47441f6f39bb8d2f390b34f41c5add37b4d2cee0bc50dc0c4cd00a40d6b7c6005f69a18b4c737f237cc6f82d870a70c6426dd644533f47ebbc4b09fd1d00339adc6f12e5058e224c021667122605d029ea1973790d6423c39d45cd0aaa35c524da5f69717a53286c0942302d2f96bdd71d2484dbb46dfe7fb918745dcde008f98b85790927665390cc8512656d27942aa745ca6a8909e601beb8f67cc8145d6f8e7ae087d2263f0c631c6769d8bc02df93f6844675967e2ed536dbe1166e6dc1088a1190f619dde217e0fbd10e0d3fd99853c40475ab28bd548d26c3a2711f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h402975542e7a2b94bac3e9bb83a21aef22e8a4e95b9d1b4db8055c4f05c85e6982be601d6b656c55df70b7a5ff51da4ea3dcac0c77835875946d011df5b401d5cb06bb48c5589aeb2575c482463c90bc8333ff505ac3c0a74cdac1d6dc4e3f2081f618e8c957b8842f3d3d847e38d55922f32a775b575bd4cfc5d299ab1025a5111fccfea2332558a0798d80d214eb411048d6cf804c6537b95966a951ab852c221497df788b9c635f19ac2e8f166daf8a309b784a794f36fafbd14bd08d37e843df6f3bd5dffb962f5a10e011511936ee36c5700d72c80d690c8669f71e858d81855f11bc315eca4ecba17af55abde842813a9febea0d6396f4684aa28a32f8bae551e42db4dc726f08fddcf85960e4a92b588261968dc60633ee0b7d90bb7a9db83dcab1357dbb11514cc99f7bcd935f8df3618b4bf55eabbd2fe9e2b58154d2aa8556d6aefa026ac51a3f05f4f4335d16910d7fed653f1f59e1502c64578c9fcfefdf308315f9b203c4099b77e0229d7c2244f0d0062c3a437de24078af24d94633834d12ba46b46305471e3a98a1d8fd070c5cc4b8d3ba64300b6e179b7c4658d94f4cb83d4530f0e151b2daaeab6001e5d8f830195624ef27e9703b5f5419dfd320ae49288a055d1f4d21f7a327197331893aad5d4be682ee3c6388e5ecf3aca8d900be5b9098ed9331257b5321776ab263b92472b4eba96043f698c2298754e1776e7c803bb4018d2260757acc5197c6e8e859d9deec9b7cc1e08541988ecfa7a5f01b1b68932d9f52ee2d67da9514e6cb6b8d7aa170ef3611aac010782ac428eaf7ccfef30931134c5e1f2bd5910730875350e43ab53b2d543dc41e00b6413b2b29dd8bfb490ccf2120890c38c96997839a1dcb5906d046e874bbae162fbf6578bd85edb6d695ad02eb6ff3c1369c397d596a928e68a9c7f698d418ede5a95dcdf5d9ccfb0d19199e9b59708019b31df1b6929d2f5fb68fcbea9492f20093d8fb90c6e1c4ccdb4128a48ef5e0eea1c12029f32dd872dc63a0f7a40828081a76d7c1962ea81ff6e17c3e0351ddd11a08e74a63a473230cd2ae95224a050de52139cfcee717553ce0c7ad306fd20c2d89f18b43a673d89602e2e539ef0f28f53dc379d03b0945d42d2acf83a5e48a6bc25cf6bb02f242cb4c5d2bdad8d7b4bfa8c59f043646b27efc191017e518a4ce72e71b5a925b1759685db4bcb3aeddb397b7111cd1cc783c5e03e3103dd8699ad25b04d8f3bfc7848e9ecf9444083385dd2f0291163f3f32245527cf22f3946580f0104b959dec30dc0885784407424053b1352cf24cae0b290fbcd17401e4e3f6430e1ab9f958bb18c54f98d5f658c2c7bf214214c632f20c731581a6b5761819512c1bb72353ed8acb3a2d1593fb01d47851c24eb36d89627610ee65f2014156458f43ad5498c7e206fde455fbb52ae1d5e4a93a4c351e56bf76d4b7f3d8323c74c1ad8935b1295056741c13f980a320182d00add8d658819941aabcef32c1cc3f9f47c2a7049d092f257993f10335953d19fac185b59214c94d9c7937bfc133a0b755b8934bf20f9e70dddbd822351cc81b3448e083d9492907056062f07f0360d79c85cdde73d62386c20311501eed1df62e8c50d8cfe3c7fab312b6b504c8fae7d974e105e1e61786dba27e6eae762be5f5d4a29b06c3de32cc38288c172bd7b8d399da089cddc0b22296cb555dd14eef9c7ad13084d1e1583e6a13d2c9663a555d4927740c19c3b055554e8e16f2a4ddfbc0b50d27c0a60ca64f17d30ae055b801c0af804e62d05ddb8d4f6cc2bafbb80a0d3f1c594c201d8d88fae2b777e72c9ed6ea6ce9b332dcb04a52ee02c4452a66abc208a9d280dd8828ac87012318378090edb2fb9f8333b5e73277181071a3f5119d35e17b68dbe7d2218dd35775c8463ab10d0dbcb30dfd7c04aa48c6bda5d1b2379485fa1fc1af0de1cd828f547793f7c056adaf31ca7826faa6649a56ef91cc6cafb94cfb35c3266098173c018e93c7d80da9b51d93671173512a642a64ca0f0f804006f5f8708e77089e5ae10d859fe6e5a236a15d02e1c6ae7549b6e3da1b8fd533107b379f57de78597640d41f0069a10514339ba7644d1dee7d0f23964e92e34690b347a1e4408dbe21bde0b9ef24eec062f663553b2eece4f9b8d3109dede96049cb00c06e75e4723412214977d12634bc1573fc4f62ce36611613cc629eb7817f53fef542d9febddde5ab81b543bfd8ee74e8612e8ceda1ce8558bb9e91b589a7d514d158e55f07ec652685dfc582c5248cae68e1edf36d4f6bd39dea5a3a017f82b6a6455d33828c3973027fee994bbcc6838fc66212fb6779985332f6d6be83ab7cc646653aaa466de53e4683420c87c8c648ddfbaf2fcd48315e12d4e15fe6d43fc19ef471cae96c3c76f1446fe75332e52e4d9cc7a5fea096c1d80fc45ac3f5c42004ab372a6f06fe3d99596797af740667831c3df35d539d4f44c0d45cae49bf93a83281148d976393d7606dd896033c5d9b77ef2804e3202da881f3c35c5607f9fb021853656b690428fed2238864c7b21fd80317be323d23bfa7c107270a0c9c6808e6dd0aaf28cbf7f827637738a894cf619406ccb0e8a49e76932f1dad6632401c0115bbcf1523b59f51622b166100ad4ed4baf75e85334a3181493fefc3c4169c079cea8be1f836a85d72d3dbf75b016733be6dbfe92651db812f281c89183be75f2f98cc82099b60452cd24a7997db00a7fb5fee5971d45ffb14acd34ca7fa7ae7bf5e23ed16649c2b79e3599777c255d1d5f1df4ce42947eeb9ed6b265615cc770101a6d30038f34f0ddcbc04145935df7a494420b774b6452d694da0082513baac807716d2c1a80995476316d8d97e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h41c7effdce48c236c6defa93c3b4afe5bace7f904caeef1915b23a181cf620c34822557911c47f691c60c14b20be6d29bde48fe66c4ddba0c13ad63df02098587d5ebfaadefb40b4e3a5969b585d45d5f02555f0ce61a20372ce3d884372b8e8fab2b1e6307afa2fdf1cb2d8f23569b9b4abf2879e5529f589dc928b6b56e5362ea837deb83130a21f0adae4b8bf57030aa30f9367c3a7d83ae2681962a5137dff89d5321554cdcce994b778c06a8de05d04617ee0b4b9d5ac0d04f56832e549e3f9f794dc8175b37f6562211761ff3d864a1d458fa4547c2641f677545e4e823752937e1019800cf8af6ef4d06ddc2facd5e00b2a09a62a754e95d971a04b08ce37b22bb82c207c409f99720ad73c267239f1f6ea0dbe4ca0c79d5ddd069cb0487befde7fc7895628f111d6ccbc25e52ffc7e1cd3565e6701dbb11c9c46db1b50b724bd9436eb0967df3c07d1a1bf652662022277be170ebee187afc742ff42b8b0670fbf9b2f260e49b647716d515aca1b5fd1af10f0fdf08a0daee9f560a30ae54335e076854a13c3a89b385c0d61a0a1d0083d672b3e6564cfdb67bbbe82726397751b716b4ff21b98c25ddd60d76f9272c14e93a1af0ca2506d565330f07d16d3e74df77432d766d48ab84d1291cd7ed2c31e2487b7333e1cdf38296f89ee93ff08c18015579aa72974ebe55322772011fd507cb5ab39223d2c32d3f35267067438600080f58a00321889a97b09856679ea37ee8feb23f3ee1d76da735ec08dec49cbb1e9b1a4c063e3edd34ed626f60d756e621831b352c5c8cdf0e2972816ee538f16b420c1804bea08b6b47171f4f129322b7429b8826a11c7a402d5241c9c9967dd1cf15418a64d05acb1131eed7b9bdb4529c65fa72fccd696f4b1562aeb9ad5de15509e2c2be683b240bbb89baa4b645e9a641abfebcb35997050c7392f61de151ee3e1bd77d60f0fbaac6d994b16dc3c3207bf79389f29a8a904462f2e3881f88da0d4e5a59821d904828559eb1b22a5b226d33805f45b7d5a41ab97cec9b90b60bd468847da8068c6b0b6b1de5aa46d1e2ad4db9ccd05a04aa6d16553842b9193e0d053da77b16e5c63711606eeee0213503f9aee4132f9b390f52adc8e50bf6880aa87dba1bd3300c8e4c16a5d942548df887d10e500406e550154d27a6d2fdee10fef2cbb64a74001b6124d9667c1898b85be10662f11fa9dfae9342799168d62945484e8e063b6d52ce63e67c412f4997d7466811a529d3f2e8a6204eb8aaf12b48e4139add9a25a0b89066b65dc4d389b03a90d6f2ec165ebb347f30339245910172742a471b5ea66ec88ed64da99fcff89efb2f365d30a8ca0a62d1401f8ef191a44613427dda9b773b198774ffb70b7e78fa0a44d987b17f8e4045894df18445638c524067c789191f78033019b1d2bf995fdb8a4bd41f345a8d9dd805292c9c06d32cf1d922695f4c3fed834cec6daf6bb586c3bdeb5309dedef130f0cc85e445db260d8766b74a2a1490b47dd187695019979678b1e71b41b18d72249db807b5c34f11b50cb4b70c5d39ed23d8e82f62ef303dc2cfadbe5e16195ec2138f47611e269011f0463da62d98602cacca907aebab06f5e495367d393f3afa9a6352902af9f903698cb115d58b696881601b6d40de516bdfb4a073da61d9d6f4f234e59f025cd7bb13335d0ca6e402e52c943eff54300c36ad0d8c4ea886b5029c228da7c1e1263626e2c9369caba4337adcff30c1a63c2af98dcfe50e7a16802bebcfee5031a4246efb8350778464dbb78983cd90739923fca7023a7637ee8b00eb046953573fb67b33bd0c9cbdbf1a144bf5b5a685fabf4b55e49b7f73b66ef91081d6103b57d056fbaec344b067228b50370e5819d68449c1ed2826ec801a9b7b8a4c7f9abd0b78a0c277a5e7abae3ac69981512d661ec7749486c659b568bef5a061be4bacf0026386a555d87516c891855deb78ca1d05784a1c6dd2a4a1af121a351ed261c4c57f8ea032f2fe71de2609f79eb69a6878b2b2470c09ac16cef6ca261b9553127cb36f555114697de1ec04fb355ba3d652e32bdc8f3f75bab7555ffb5a59802eb531143a9a555e41992ab4ac5c2d58c1d5d222b48e282b0e4fa8a51f89800ddd906ac3e5294c51a6276a70fd4e8b03dcb9a84bbfdad0927a9025fbbf1edf994230121e4f85a3d79534a0498a2606e1ca9e8114d16585161582bc539ad1b0a4e5c60b55e35812901d8919e935e1c0ab65d74cee02a880602768c0ed0f82e545c7032a66d2ebd8b528728020ad910b3599b2fadf6a065e6165e7741474cce0e5dd895feda64df7d3767c1cd75f67f482e220df8ff8b48260b1bf818d7bf41e794de3572f9b97ed1379bb5fd305cc356349ee31dfe50c3d65816d4413806aa8b2c4fd74c545822b32c355c8146c8888bc978f936ad4da32d75bae8847fba601c2ec02debfac562d9e29aeda0cbd71f698fd3629ede19b3a03f8d2a52112292bffa367f8602b03a51548287ac8b4b956d0599d2a58f535b570f2ce7a98d87ce42eee86f98fb7082fad2f608294f9623fa66369aa3b48bd762205577203e7f592bc8ad1a16342677cfb42a337cf801e54edf533df771f2ec786d1ded88fdea7ca863e215a33efcd2feabf6d278aab3a23db748d22803a103f0fbeef6b963f8abc6f8b9bddf141fbe532674c3f663da290f06dc1e49f0ba635d9a3716ba8c0c07a1170dc357daad14bac3b98d64ef44a92fe6da967d5c08278525afe4f53fb11cceb10b27ea5cea542c7f12d649907d57e3e528bb08b6965321e854bc431152298f7035f87b5a79598ede0032a15cf1bd2350072526c058400c594aee0ae88e4a7c2e8220b0b5a893992594e0e6370bfa66e12f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb9f4ce172db74442c448271b22619ac2bce1f2c09c5cba59c93c28f75f81494399c476646d492ad557f508125b92412d7dc3dbbe9a909fb5241d2f934a8b9beeaea8212cffcedb958c3416ab4de8b9aee0a3bd243c0d1c0db74c53b0f1e36e0412c2d99a545f16291b955a3440ba1d6a92e84c83bc9532d670c4bd93a8e2c79590f01008ed417167a980a867239d7d1d070c61cac9684d772863a5f4b4d02dfb2f2c4381f7c3ce5cc388e1371bfa5ecd9c95637bbf92ba02668432d9c942ac35bf8c892d871b41cfcc27faf929533151efb120066aa2cd02350149202ae37be7c29e51b0039808f2f6ceaf9e444ffac3d0a89f2c435ca8eb024112dac0c315c85faf2b1e7b6a462ea47f9fd83c2aca66385cb7313c4361cbac91270e040eda8f0f4f8a8b8e976460629e11552146c79cc6070b4754452f100c0ae10ed12ef4e67707bfb37febfbcf0f889f2bebe23fecb44589d84f7fe59c184adc0584bdc9d36e334e58912c36dbf8bc84adccf68f33303982f53a8c98326571d96e549aab87b88ce3933266f5c60064f95feffdcb025b475872ee7ac7dec9f1d9b8ddd8cdcbfd74f92fb9fd8bac697b08da1306fa482470ebdffc7093e7fdb2c9d2a873443e51cd9049657424a6b627336a4ec2e0876118c07d528e10f1219ae0686c0bc74e4a1fcc7e4e7eaf6fcda691084574280f0490b63654e47130b70275f0e39607ce594a60391af65a02165ee5e04c8276c81e17707b86516b1befda5936c7eddeb6c1c96730b0a44de230a412162c77100b21e1701a98c6f17e3486361704fa7cff0b005aa795cf2c47b759ca9c61a52420a8c09dcf3eb02c998745e7aa58767a7a2b49402a23c1925d511446e070914d8f3031c59f1fc293333b8e1fad91782a9ac16ffc4e37ae94431720dca9b58f19c117687218c8d060ce3a65b2bb36742ab3fbfe3f44d40a3d1adea5267c2ec76f17a8e50b204768dcc30156531d972efa54b8789c52b796df9fcecb9652ac7c96cfc069bd7b73e9e91022ade82e94b8e15b9ffde3dea065160f32e32a606ad7d3ef9933816223664f9053e318c72eb1efd2e41c157cbfa3d8cbc8bb3ea423ff9639bdf128cf9c3ade1a629088660d8d91db943e3a41e556345207371435d6253ea3af13690e5c6770d901188e63953e65cd3d4e76e2499729899ceaed046cc84cf4b7c5c932c870544fc7cca8d9ea0007525e993a87dbaca279a209200a35284b2ad7c3b7139256afd6825ece57d980c6a07023e0d4f4fc6ab436a558ca36acdf99f1eca01d4e1e7dcf9763aa980ca4a246f1254297b8ad707595e0d35c54cd9c77449dcee67629a3f593c330855f32e2a336613fbf517e38bd519d035b6f8d7872713be20e0124d7908ba740a597f2a2e07d531eabd20293c4d7e9168b8e2a49e90e5afa4b7015ac8293f2a68333c67317e08a4c8ed7afc48d6a2111e0b74742fe6aa77d423e5b24b0c72f00046a6fbc7f44ed7ff277cd7ec7a00985c20bf7ef6119fed731e79d89699f5b6c19caaee2b407a36fb2910392e31d158b4609bb23026ba15badb44fd3b4c1fecdffa35a5bfab3f5a0aa0dd338527237a43d5ed99cc382b5e0484c353df8ae816cd2a4dd327bf06bb559812b7ac9ea96c5875f91048008da2e5fa3c6fb1e739b08056228ac7a671a377f846bd71bff0fbcd49a8a02cb9d7ce8c40bfef243ebf77834f8357e87f10636468e42d0c1040d64939237eb97aeeafaf0795ecfcca51f1bdd3493863aabc32e05745e70e34556b1d6bb63e3609812db2533ce397182466ed9a8b505674378e28c1c4e35a13d2effa3e4023b9930b580d83b98590169f5f717ba6fd4c5b3de905eaeb06bced39291488d3b6c50f63819c40077237ce415d76b695ad7cf5ff89afd30c177ef1a521e19651097a84a03bf4e943d723184555548953efb9efef37e795ae247ef24c41fd27b1010a14b1e57059dc32a466cef8fdf89bdf61eaa2b2658b02c1f89a27470f107d4d11bb5575d95c273dcbd99a701dc04c31d332cfec22dd2005bb5ba99f19bd67149ee1d5b4a7acd044a6f6a2bea5ce9e624b607e7d74460e2779a3fc7b13f5299ee5d43a58a0311c1215854746c09efffb32f2a04b8f467334e1edfad5c34f9379042c449e9c7e358d9efe429703df6835f7e6ca284b7b15fd114570a541b8128bbb72d1527bee368b3ecbb41413da0d678a79d7d3f13e122ce3504fda8072a63cc07066445cf9da94e7ec068892abc82762abf0758a85004b047139402d9c18e6b3fe1328f4045ecf012a8d274e01849707e4db2bf67921e57fa1e44805bf067719c3fa8ad60facb2c1207ed35d3e4e6a40673fd38fc114881e9f4196a96de73f975de8e8a48c09b03957d749b90be538086e1436c2a6a3491fbfeacc8a3c91af00b52c4c198438ae6f08438e3bd670469316fd756be9f3931323b2b95a036e19d243ef6ea944adbc1c53d6d839767dc8ae22b37444272c87651614d8d89bc3ef0af89700a826957f5e66bd2e79ab1c687fc286004f6403f79ed7fe3e5e4cb52f49cab9f6e1da983f11cfba75868cc40c6cc874bf4d73dd9411b7173aea42b8681e3d7cab9b5dd922a4f6d19502d407b6d531923b0395dece28c28d2324f1025cc7da562d55f948bcbf4953f32cab9057cbf1afdd40100dfba6a8586029d87d88c414946697186ce104cb0ad8efa5016dc01e43ab57958ef8827a7f7b49e857dce57593ac323672e4071ed07c53cdf0447cd67f0a60f4833d7e7b0487a45c19a2d7fb356456daa67938f4c9bc091b6a9fccc1ab334257c62bed43816e8050200157d14a7f9c2184de58e54402788139e6f8a64dd7276cb4dc0d51aa6a998237ebc9d20bd51377e30403cb914187749f5d73b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h504c2ed5548277446bc81e7d99817f6c2131cebfdfd4f464d80b749854dad2bcc00e3256f14f43c9ff81e2a7a3e915f077d27f94a72bf3b1156ccbc6518d52319c1e6c944b6909e304f378151862d2900e7eafa259834100481737e1702d25990cc764c45e6bdedab314f6cfdff45ad2fad77a94a42940d956b8cc7b3a3c757476406bb59b3a03170a707f5960a4d38f40deb79c262130af80fb7e3ed62671b4f5e9a57a2bc1c012634acb89c284dc01f79798c348e8993636279cd7f2c9b010b3e818aec1858b8ecb7b08028df006e9d5ac1dd3474d51c4663961603d428410fa2feec1a673d4982a857e1adc554708ccb9f01d32878eee69c8305c6f46ba1fb8d3fe90a455c20cead9b2de3ed38c7583cae73853c0143d66e79809a2791325fa64a2fe79649768c40145013a94c0d991de55b68927b6273a6814ac68faa09f09413e53842a24fc552e52056c40e64a006609ba682831d881f89ef27ba59b678c85d9cf8dc12cd8b3718fa3b241e83a0f122bf1483c17d5426d11b06a8a8218be35d92f05d2c2fab9c5fd7fa4f080e79b1665630901419f0b083deb68fc3a64fa8ce6c68cfe7042a13080963ef91d9a79d056e179792a55273964b011f1961a58b69790c4e69bb6a0d77155aae2642643a2c8450893d9d0a66b5d9d8a80f96ab8fe7bc7f78ecc74f13a7cb2f2438e82aa2b04537a8a9e3a44c505baf918506394659273906c38851a8894262f3abe95b4d897abd4569a93cdf53b0f92da231e707931ad59b9f317fa51f5db6d3c499055a50553c4ff4d91c1a3fafb5c161a968e31e2c50b1b93381bd7c5b08f2b667a1bb6ceb40d255474b559d486841c45e8e6946483836b9b2a5472341abc882071eeceb9d938c3e49f1f89651a1d929ac276334cc47ae8169ffa8a9e6034fcd78f9fa8fdfb6005fd1bf9161b5dd7c150070b3c91d07eaf1418496e0af1375c14ae6bd69e7df3a70bc8ad69af0571ac99d1f3c13d978e7b835e75d9ecc49c93a0867322a1fee1adbe60f6bb85d8f5927593a917264f978c99304a89fbbb453caa02a74c52999fcdd4a6d599ac826b2525f750f98dd2c596fecb5c9f04d3f2d0ae6bffa5d4a8b4e26b84ce1ff46c6ceadffc90f69ef5dfac19492fa7dcf93944bf100f8d12e6562ea1eaa89b75891ea8e14ea61bb4af173194e4c9b44aad639701ba3adb5b1d556843674c92015195988c2f8d23f455e7891b31523d851f8b22af6bf60b148916e0f3fcb1861309c939407dfc14adeb10a65f2449a95e69ddb1abe5a044d566eb32da99308f228749260170206266625739887e94ca6e7df5b87dc51a7026d0fca9f07fdd470d0da2718d8caf5fb5152cb30351475d9964d841c7985dfcf3c46d95d31f7821a13c8e098850b83b20c3f3fafb8a3f1ffb5069de1b8193e950b393539f3f9f8b3c919247cf0510298becf5b492a1d2d615931af0a79f152b24745f2b7106e2f1cccb8c1f40c7d14036af19a12fd55ca22fc19be29a1f1741cdeddc1c91d37499893a8671d15128c215c0033b135239d9c0dbd332ba07cae861ff28496cd966291b3bc0a1c60fc3fafcbb4dac3bbe13cf223caed1fb8a9fc5114275324465b8430130bb26481259db072da5567e0b56a20f54a0d27a075a00c76c36884c308faf8f861189b6c26bec8b01843034594bd07b0f38fc6f73d20291c26ff62899ac554f6e75541724536aa80c7833e1c5c24d8daea4ecaf025821279b35e1921bd3273b2bdf459c468c06122830c85148f7fcb62e57c9a81a601df52db63f49a48a92ae924b30b4acf24b6eb565e61f22319d4acb5c0d023cc63062139b10cf95a22521a65b0a1a53dbf39437e1890ad8115959d9fb937b0a687b521af69daa6306f9155411ef7c36a8b7f0d51bf652e31e67c4efc520f90eaa5ae530357a8c89135f81f22bdfe9f6127def58b62cdfa3bb2132c8c32d78782a8634717c8e3f0eb7330b82ac779a09c86982d891a8c882c9d26eff0c0957f95af8b6e998c54e63ef9f9027a5fb9438e1726fdeb973e7f6ce731c1edca0ec9204cac5bfa3aa2e538ce63814e8c9378ba556b8f20aa359468765d3db1555a83edfc58a16ff1cffe886803a999fcc1f340f3b9f550abf03def0a688be93fe5d36fab033416bb21c4c969108a6c8b28a1d7eb129678b07af726a6a941fa5c7ae2aa3db03e5c9ad3cc5370d33dd56b2df96eff8aa2c403f37c4f161d27f4de6e657c6960da09e20fbd29848c4c550ddd80964455fc48d7a34a7e69b159a44f71451666aaf27989d3c36f36ebd57ab7158d606ca5f5bcdc88191aa21443798cab969362c8d3cfe7f486d92401495986893b93b6d5912847f467fd632745668ddb99ca21efcdcddff5b4a6d671cbd01bf09d08512399f32dfa85abc0bd788bfa7e2c214e653496312528661609ecd1e98e5ed0f20a091288c5889383875ca3468017a69b5daac1769dc24d8545c5d01f007a497522ccc53570d1ada19fdbe00934d15d01dd3159d99c48eef9e374512140786b33828eb5f4c507117b176d6e405b84a942bbe28429f0bb3e069ff586cdef4ba0b9b39c5c5bd309af5b40d31ef594cf331e86b9702f686adda05c67bdfb567a588cd2f071e3fa39d2c5c2ffe86a53791cd490ff0b7a90c679b6c1a69b495772a936c8482c6ae1a7c0c039d51fbbaa1e51de11eea7006d61d7dbc2bad1e687775b67bcaaca75b776d0a11e51dd73aeec5943c9cd98140560cb01d289e1327a0c4c8b7f3d625ffafdcf88eb90a0a8039726362d8a8db85f2ff2f443c0fbc5f377815dc904a0cdcd464ee0d8989a49afa53224195a560fd2202b91a473800662341b19af7b08c4413a31ed8bfcfc61d9ddabf2402d793a631616905c81b9288a12d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hea1ffeecc738247f121ff3185f66c5fef7bb55fd795cb0435433f6e7819f97dc409b3afd80d7562bed394829831426306b450f8ff829d880dcc183392b07115bcaf4eb56adf8299650984f8dcc4fdffb9803ce289a0c09aeca01a756b754fa141195c20508d31789051d4a1519a6ddc1f2f3782633d12612a7b61a3101148f9568af23e02b88e73467441810d161474bef14bdf6b5259e5405d93a53e44ccec92112fe7b706c115a9920e0ab9dd0450fdf72fb2dc3b9e21334ebc4b5373d6ec220fcfdaede8d0e5d989016d6ead5da2f5d5eb83b137c0d181e5f9875275751fd4d508fafd6670ac4865141ded363309978542c73baa3e4615b64014ccc4b6b240a34c4b9670533123db4fd984c7125e7ac52a1d78f45a0f53db8183d409c4afa164575bab9a0f3e7f02d221a12682aa18b12eb78112bfa1fa4e8d5e4a70607df8a39c9574580b38267cf1cc8fa0586f85b6ae73937433f23cb459a6da71b71e5052db06f02d8352840b934281a94770dac21cd6c97e81d98420c6d3dbddbee054c9a4753972fd6fab509a2f30ecca1869c98f9580afaea1c02d0532f577a05ed7b419b576254576571d2b3f742d74774e4c5c7f39d50313b15bb055f09eca283c45509efd057399e9629dc948796543cf4acaa7fbb91a4a981c0d19d804f74fafc4786c452ffe99012bca6cf7524132209850f696808578e0a8cbe257b3143e6955d6a7afbabaff833caf2f0c6500a0d991907cfdaabf72aa963f0fb68f2d5e7699b9cde6d673db81c16a3cf8211d3bec286939e430d6c3c460e37c87de8193dc4ec72c2689c2c30e512f6998dbe7af178d66322f7d8f2c7181fdeaf45ad8b4c30f3b04a0c2fde0c4cd7b6ec2f82ce5d0f4825a0a0ab8c6bcd3961b678cfd69c47d3465be6801bb5c7430380b713e3b904f0118840de76626bb93f9b3e6ee6f702d0dde11eec7581563bff6cedd6c9a4fc30d41b2fb9c8ee6dd063a4228188098bb964515007ff13edaebd5beec8bf53e89c318a974e21486475933ca87d48d653d1c49ff8b5d503b4250799d1103801f40823dd8adf978d8be3f35b1cd73c405ca5fe71716d6ac8ab3a0bff94fe0105a2bd33e7a9dd2a89048c3708768b34ff1f3b3bc89144f1118d188479d9eb01ae333f8af704e5503708fd087e25f1838311cb5428b7ca5a3c03482fdd84d2dbd27cbd05224820302a63b6d5188583024d6ce644b211f72bdd1cd88bff5aa1c7e6fa75b05125179c0604c1e822ee0de7da293ca7cbc7b648d0e83e4a7c7cc69db62b358ed19e7f501de66e2084f67751ae5c986a58b8b7ff45d369622e753522cb02fe4088d6a07fdc835aa8a962e6fcbe3de99ab87d3f1fb4d1f6d24a95e56bd74c51a76844d2286330b62f432d1809a9efda62929fcfa6fb256b7b38bf26e4de4f697b422eb47650d7bab6d49ec2dde6ed98d8f887c1f931ac83037e4400192b0c642c2c8eaf537150f8c1acc37dd4f9015ce472d60537aef7a30c23ae36aeeff78dedb846e5f82fdf29c5fe5b853a0b8558ce60bed24185d5631fbced4578f927cdaf6055b9004058e78b02283f728f500e7f75fe1f515b526f979382e8f99081ab88beb104fa6eaad8155f4f2765b748fd0073f217662f847542af5c4673886e3b701013e350a6887ea9e654c31c0a3eb32275eb9cd227c056fc76cbb96f810b9007ddcccfcdfc7a8e5ca4ee04b53052555608401c4c4d50ac8128e38032954968aaedc5630ddd2de5ae1ebf918da8c021ff916c0e45ac7a388746397af4cffc8ab5f9fbcc481f22ba0e0121ad468823dedd92c969f8ab63295375c4b1263eb99135f31e82152e5de1458f01550fd65f846297828346b407b756f019dce06ba279de0a7f3762b5e15ef2e8b861007e62a40f939baed232dd02a0078ebb17164d05e71a0b773bcf344dcbd3a3bf3cd799ea44ee445a6ad6fdde9d846dbe5ce5852e7f767905d0286404f2fd565d68f52b410fef1c5f27f985905d32241392fec441c6e8e58d11db56fe225ac2eaef2de4c202e499fd6f396eb00d060a61c82336afa436d017d0106db105d35473c9e427082c714350b64106071b0562718c6d34d4ce33e64d5c8de81e951f070c19c9cc0336eead57e8281d042243cdf6b1ec8d3757e95c1cb5fb72d7f7e58a8d33bf56eb3450fbd67e59adc1be783ba3d9184d35060c5839e66e0b1bf7e36f674476b7d3de4faa1979a4815b7b17f856f6d0f8ec1d8bd025391e58720ca6851572cfd1d19e51f43977767eb37d985ad1e680a5a391f3b71f5d486fccc29b774b75fe846d897b227d95980f81f8d353a14482d461d496327b0d47c3a1b0871c13e671c9b6759fec421f9f4de334ff3810b111929df95d8d1b1a825611191f219ae64699a503525caac3614733a6bf124cfafd86e116d856344b87b74edefb5c34d1ded86035c0c5d128f45c29dbeb3b7a01ae94955c33a3358448c898f28c0d0d2600bbade39d3628f18e7f0830a96df62daf9ebefa657e08d5b4b622e0600afa436eeb94793a594d1c0d1556e6b14b5f5ef410b28f716e8c409647551edcf5badae301e276906fe54d96d38863ae03446c6f9274945647398fdade95afae9269671c39253687215d53a80e9dce677c6f49b490b01932b665f2401ddd5822c391c3f9d0f2f7494e3a0ec6ded3378102802eb2e8e3cfe2e1df92d4049467af95fddb389fb51b96733bef928d316ae8f5ecbea4974129099857ebb8f0f259c5c98c706fbb7e7eab9104b5537ddaaff512b01d42003e3cce7cd2c086ab4202e9d4672f468af25b62c5685135d18f34a02deaca2cbef4f3cc71d810625923c81229acd78da25bbe63b851e9796d613e6597532459b6d740dc28ac2a75ad13f6071923bb63;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5846446d4d675422605bede89b2195772e12960700b948c83fc109ce9fdd98ec1129574975774785d085c4928260ccdbff4403fcaa8ac2b74af817860de1d0abb58c430d1acf81a60d9c46190f27aab3464a58359100ce756ade0e4ebca6b862b6cf35e443a171c57212593bee30a73208cb7201f6ca5c3bb1dc957d6d276c0317e9bc90d4bd95beafc0e30d38aad93ac7f4202079a9f7abcc970c5a608484701b9acfdd93c089b9553cc640ed832c176b4e37d7337983b12a9c17c98c26e01d8a4ded21a42f58ab4428aba4cb797f3245f17e5268cc5950488af043b3ab907aa185b5745d6d90d073b8c5f680e0795fe3aa03e15bafad814064ce791b13e64c7e9800e631b79b889ef41eca1879454166da9937f416f5af4bd030c84c85198b7d6cbbc29cfe76027f07641b643b38fc23dabab3e53d7938d2804f1d28bf2b6314e599823ceda814619880886cc825effe7b6e506cc8cc70a885533d3279deefcc7270ca4396b0e77380bf4dfc45ffca3e39f382268c0255af1ce061b2ace33aea93d019c2fff85c7bd1db72439480ff4202bc84ef8ef12639d4f760ec1480175cda8173f8f2b55901b3238d1eb7c6c08c07f1093f2a98eb9db2b031850d95288b8b0b830b554fa9562821f8f7e2c0338a628cafeb4bfddfd190c5addbdadca57f67fbe182d302174e9d3371db32dda088b081c6916dc428b19ed704ab6be08d4759ce7b6c66c969e461ae7a2cb669fd3a9a365e895568793f807a2b62ef71df1ab93b2194f96c0d8be1bf940c54336c97572e5efa06fd7d4b02f4161914e3acf552ae14a46024ddaa2972c99c59f83e5379da3097b996c82cf1f5017db840dd2436332f5ce6c995c577de0b3574ffdf6c26f60dfe524701d882f017743b1b54deae22e4cf475e1ebe36e5c7f8faf299d82203c9ffa87759d877746f0a673c3f0f43f85d86ab4205fd3c360ab8838f09a54475b8584c5579f2bf1e49853eeecb35452aca24787f55a8317396e0f6d1e11c04523d77576ff3c26de6c795d5460c014c01f1f8eaa13b5b38eb03f7089c1d262fbc10c0922ec2d4b17e6787cc290150be2497c2f8a9491dd003ee531dbe1a7492a0bd410cf8be8eacc108f1391bf8704c078665676a49eb02ca840d1e84f21ef64401f1f4b7fc54c479c3b43c66f58ad8d2e6f86a597683a4fd8fa0753b6698b21f2f1beaf7cede5fa5fabbc38e6989c251b1b4ca7284af79944060194fe414b00c0612efc321b6b17dbda9ecece39184eb56e6a8561b5d0ede4d2a9821cb4b8539e6bf90afae92e85100e1eec9bee3ce1eb96eb203388a2669f41a47a16dd17f09faca214b917a63b0c5773a68d31f4ad03215a7139c5bc682e42c991a8be99a8e2f98ae78ca141e2074d25d02b15e0ea43a5d7ad3234de4d1bb73a4e12f4d0e4143efdc445d25b4cbaaa88fedbc0cb6d7b986fd71a373411d6c0ca94cecf410af764d15734dbd2613dba575df675c91b7aae2ac89d686d16374d017396a336d4541daaa261e1f7f9feb95365bac0525a1b881ebe7e42454fd285b6a995d8d9bbf51aca7a6d94cb3bfc3cc43045f6bea83e78cc7e40a5249ae6888db8590a3e982c765600ee3bd5d96e48975d4a74647129a8513ef6fbeff6eb7e7c9fb93b7f7720c1c5d90ff301b2b1913a1cb7171e55baa742aa6e93d59d638a3fbb47e20672d499b8f8dcc1d854fcd23f60bf084a6563c4c74a7462ba368f09b53cf37fe86ad3d8263cd93319558783fe5f7a6c2e42c2faa465b60acea44b4fefb9af49c4466fdcb41dbb7a1400762e95f2d4de8c4df2d702718b3ac18d8d94a68980e5848064e0677adff2998d01b03620fd242b34bd3869974f5864c8310bb0956746b3dbc3504324de88661ca6c08698636690b3444d30480b342e1cbfbe69da0cf67758ecd78ad1d9b6bb6b6f8912e5bcc6a7e48580227364e69052b534110487acbb15fdfea19ac267bd9452e79292bdad18c2a53732cea7367b33ec826947abe54fc948c56cd38b08ccddd5edf8c51c02e5b1a24b0124bb8cbc6e7b7642b6cb21b1c5743139fec398f844655f9a5411a537ad7690e07a05253ee47e5f96ba0072afe6fd18f37ba8840a33320f960a450b3ebb309ac437abec29c36b0be0e1be84eb6e3dbc8f08638a6b0a6b0241f2c2602a1620cc3bfff7c979967bea90fcb16b5ffee45d7edc5aa908226964bbf5e15fb22bfaf3c4a4fa043f2ed4daa51a60d1e16f86a5d73a36b862302cf40441835bf4a48ada7fdea73774a45c8420b70ad1536d5b9aed13f41d8175a0c235280b1b957bf361d9f01746f6e1244aefd33a1264d5e8f4858f83e40ccf58cf67103bf5f05de504afae2603070ea4904a7e41b5b63117e9c5052c914d64404032342597ddbcff1635fabef5823aebc51c7a4977b86add79793a365467565f6dff048a436d7ff3c08d8ea205bfb5f72ce64c95e9a592b02b9e2e0ecdbd7dcb675ce192699f618408d67ac76ddec6a6cc3d822c5500a8cb573eec45e7bc5ff19d97924f3eca35ff539888039df7ec6b2b2f48b15e9dbdb740a188c95e5d37c357162d8759feec4a4de9959b898930fe822e8fd90ffe1a1709a7679aa77572280d2c391e56089f737ad73875f90928e4dcc4fec0d18d3f6f0fb334586264fb1c9449a5b8d3471e280813282c3ffa5b193a8470e534fd8fd80a0ad574ad1013ca595b981f27ab2889b3df3897ca5beecf3929ea7e548dd451e1ea9580f5d93dbe161a8265ac8b65154bca2e6f0c099e45affa759a29af74e0ca1b64493ee11aa1590af3fb0c54ab1a72ed2d59b97bae2381ef006e5e2a032b86ad906feb428abdb92c4e74ba165e7183ba68dafb26ffbe4aa51f5128e87028d88ebf8942b874c56f4519f80;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h703e51660c44119ee1556e3c527da53b0d9a6b00429068b1fa9816d5f6ceb47aadc83001aabe1a3ac3d41555a940d3bf71e14a0021833a54967c8eab325521c118bea8b5c1f0ac3964062e9d7d05a045413f63bd218f2f609100664381c360f7284a22e1401b6698019fb63f1ac44d13da6c474c71eee781f03b084cf079af255189463fa75b7b28c237f1d4f6956f7802e76469e947c3fb45b871cd8408af55fb5bed69f96f31fc4fc9546633bb8174e484676b4ed9c8bac110bcaa65a2fbaa4f92e9acf873bc41d738a454c42f4359f946e94dd90d4bd45bd0d5335866710a29206124fdfda50a29e7a6f3b7fc0d1d861d86c7bee3213c4ac216295ddb8fe4c466b2650950c03d87ca36e34c0277bf49d38317b82fe16f6c42031df9e75cad97ac13e3b00df7270bb12dee4edd82ee2a81bf72d6dbbec73086aae9ecf165183a36fc32ac771704f9e5debe68d642d849713e5c7e32a9488891c291b719f397a65a0f96a40607438a7472f4a5b622fa8f651bc3b565c0c643f1798784bc156afb0c5483ab35e0d4ee41f31ae4ba4f25b9d1f34d01396e0eedecd7901ba16342a4d21132ab5d76dd2b085bcc3783b4e430b040fc549263b8eb2d454bb708e830b1acaa9a3de9a6209e882ed315e4804fdf4c02c2dba0ed17c32e1682cc7a9333333f20c63598762e238c4fa1a73bef2d44b49acd0fa929079d0c3b3c7db043bd3009163d8594974cc8b738fa2bb02eaf5f46f0d65dfdb4d3c40f050c1809606aef6e1c1c69fced179377e62f06465031cf68fc6491c9244aeb2f6c8fb8567ed9477abe5533ef7f34ff325bbfffcefe19c02d2ba63e367e7609fb3cf55725a15d9d750959c05e4f17014561c040b0052fd890e7c737f3906ce71e5682ef9b160fb25299664404fd39623f25b9dc9eebbf8352926805c7c46497a814b8a3b2a7ed00f706261e33af26917b7ccc87bedcb97c354b923e01420a23ff93ef3b439a6e996cc3d149f6932984f6e87143e45805b56195fec84233bc52fb7a30e5cf20d634ba9127995666d35f4ce0c4574ddcd8f18970d2bab70ec6e4aa870cc91f844c976ad794f6162d97019bf862313ef001616e63afaad56ff75f77dfce8114df4859775b5727f7b039c3f69838d91bb275b75a997c3ca6bed12772ba187ef0544991ecf8f5f23d8af3350e04e26ee56b1f03409d9d9d300e1d4a5258e4a9a8c84db50dd9a7959606585f6521cdf9e56cb1532706002d08f6a3f00a1233e40512cca7ae8d25212a09f4741b974663a71898912e4344bd27ad888f7a02354b1dfcb9348beebbb932a1003d55a5c6a866e407fe57b49a3018567f3fd32f5aaa97642b970dd721f1505f8678c3794c188e281c381cbc84e2efe2f0817636211cafe2936a3adc993381383b4c191386baed22d19e66d015ee8842c060902973d27a17e5cf70cc1fb8fe571a82909c5d72c92787378117d1ef2c1d3da8319b3ae305b01b543938983bc6f327a705d16c7ca283b38b09ef15bd21cd27a671ebcf4109372881cfeda7bd98a484e2d1480ae8b5b782e26be430c6f615840e82e7c35328c983684c432c20baa83f9976b8cc65eafe00999638c284ad9ca8b223720e4709c949d2dbb04e0d26b973c21acb4d58c1c5e54cf03e99d5b46009e0948258cf949388fbdcf30b8df67e94528e72da06189b4eb27fa475588a1d7d22eabb0c6698782f05902c79063d7a5c9afb477d1fa40995a43bde3416ee85306d3ac28aca81ae8514a3d8e385555470fa94d5d77f24206c364b5a69b6970de7611e49c00d2f04ea5cf3223556ffd13c3293e7d4964068add03dda894ee2a5722d71922abe8d78b46e62b0fec807901b08a1a8d9680768692be0b9c49803ddf2b2e1287102a8f5cf68a813a151c330fb4071f84a67f4308d35a9ffe0d8edd19ba34de3601f3a696a503bb09cf021f9c5f617254928b77ca1038d4c114c7d259b2d1aec11c5dae9bd1126a0c1daf53402d80bd70a767306c567a8df079f0b91cd691803952d338f6f533cd01155f83aba4bf022b023f2b218fd4527ae4a8aaebb2b21ac8969bc7de2b736d8a5e96102e84d517da9e7e04621042ac147eca76e7c8326e33808164221395883e0b7fedae780747a3700d27fee2cf6fa7b6cdf2310e488cfa67f2e894d4cd231790760bd996a177e10d4b2b74a05ef368cd5e188212c4149c503f9320c6aebffed7427d9ea06f5953c407d9eccafdf2e70ffb5d911b57b1b0b415f4a9c7b112d587096c9df8e7b5a8215fdfbbfe5f9447953bb792e3ea7b777602aabf841258cb096c688cb60ac50c4557acff05dd7652196cd7484cef08f4f85ee61dfbe5bb17889f40ccfdf7362033c09ea95ebe8b2dbabab5c0d43250e892d3970e3d37ac08bc1bd762c415a94eab23c1e8cded07bcffedb8d6e81bb501b5e851a2fbc05cff44eca4370da20c0e481077a97a4e34fe64affce2b898e4db8c8d1dbd91405a212eeadd090c225aff8c3bcf49179590216517d74613d95bce280918b9078396564e30b091ea1834c2161aafd43d6fec23246392e2e34f23d5e02d62215775b9d7a46dcb23832165b7355c04031dea1bfec0d53c927899efdd54ba73cdea4fcb20fbd2f27bf1664d28208719c8a7ed0aecd51fd6719a73fc15f733ce3e2e54e3197066f4d309190c5d9180b886e8a7a8c3d9fbd9cb58817d61e68636b2fcdaab0b9ad02e6fbaeb87397f8d0c3ede333c81f252cc393f148be12862c1ae825eea01ee1fddcaa3403f7b662f749e23695b8ec80da31d10d8511b8a867047a49639c166440d1edab34dea64e345c0ff916fa9f4635482099efcf2986d726ffe43c379b5f4722c2bf6d81f739880321cf5504029bd80657adc088a3c66e7dca;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1eb1edb3b81fcf0e50d60117609290eb73764301f32d7fda6a30434f4c890082c5294a526dbed6ada829ada8bd3d8992c719acd465f42379623e8f5d037dec2ac9009156ef50a1af3b86acbfff56886fcd06efa880d37cc7eaeb36f3401785a4d11c42a3e9590e4c19a818e759db634fa223a4b95f92a0d3e2ffde84216710702408f1fd07398a5e3d26cb92496c9cd43f96564afab783b8702296d0b7ba8ba2de94966cc098c78e9f38b8a50e56ec04a03d06829291f139e69eed4f606e41336a1bcf68aa90c08fa5825e06cc8fcb993e24626368e193aaaea21bd6437246a5dde3d411a8d44fd6232703ef3aee9d05861041e25854bd7f93c4b2c291cfe0182769c056902622d6cc82aa5d436d29ced689a5ff269fae489aee0effb1aa2b0047adff094cbe8819128f8706374293a3645b6513a343af412cde5f35abcc83cf96b5c144889b4ef5cfb240239b86b12450fcdd41aeef6d2fcca0c9125c2d2eb88df0a507dcb3a685d4cd4e417963dc7fbae02aa38b077a0ae6e427edd50df4d5ea5c12a64a359a09443da5d6e378ac8979bf2f43059d6d2c395c025f1553b8ec00033506beae0dd634f6c2cb0aee8dcb970b32abbe0164090d90b47c6ecdda9e55be3a73f9a0ff904fb9cbaaa32798ce75ec785817d280d67a8cd4092483800d06fca098edfd7450ff8b5dc3fe9bc3ef03d947140e19e739408113c084e7f1e4ac57af1871982dcb646a5599fb302710e662584faefca05a7845e420b638a08027529d66f9a42169abd699b512efe077a5c0074aaf3aa5f05b9309397bd856cde35f2e5e551546ad3641725853b724fc7d11338d93dabec1adf8c3ea38057d2e76e989dee313721aa215a206bd7e63b65716146358b7fe3d17f2145138061527541746da7eae94ac3cefa195f6f72cd82f3065bac52d0fd9a74aff2861964c7d55eb50be0354a5ebf380b54165f569a9a19f435a916ecb63c159264e335c95c6b315a723fa8a150ca3df2d3dc33cf1ebb0bc1438a8d771512a31573314546a58f84e98188bf256e693075d38a213461c413faa7b0c1be2b6f426236bc07b48f86015cca8df4caaf9baa35ee175d6abcf53d63869d92823dbffc790c172a7b298762805f99546efb838e41b1ce80d8e9e846f06f376ba986f4224eddda3bec3b9e554421ca06348101f69b810918639acb00d0a1a171e5edf29177d11d65c0f1e38209edda07638447c9f4b35cc279f8ccc3ae725b40570a744856747b05ff24b94611c380f117b925845aa16a83900c76bf0f5f99147430e16657adf07e50c7cb9ceab31b77166b035c27378e6daf5b9cb5728457a13cab457ff8f05e38de38ebadc5d86e802f67a9c8f617555ce3950cad129ccbe80ef13e7cd874a505940c1ac741960d7cbce66899a904dd8effb11055a6ea6022fe98f318c81fb8a685987175bb6a99a90c26c10450e0a6decf43cf46893ab6d52cbd6f66690dc6353d995515f80dba274b7e10b27188cb7c58667e33063640d71a0848437ce33c0847e9519e7e7c3ed8a00dd30587dc636fa2c317e79a3ec92ede21f8cd6ce77a5a366a6746bc3215fa31b933d83f0e55004c95ba78e55e3e85fc3c7ba9c6b69a51aceebb46fbcb81d5d662131dbf5a6a2c5add25546001095f537933b77fc31d9a4653676dc26c411c9749c04eb87fb30de03a0124cb01c878c6be59d94be850591730b7831d296f2a3020514b4971923a3afdc36cb65a69807a68a24b66397ce9ca6de17eca2694ed570be3888d363b5fd649db652d0bc72db829809bd45debe4f0bd57e31b9567e8b00592f4f8e40954eca87e0337634ae62e13f6604350ccf5d3ee640ad3ec43761a8b87045e33f0751539a5ebd1f713c4ad6a97c5ffdb3c901bd99890f7c4d46c7f477315cae4e7d9810d9382357f5484b70e0305d8b82174019047c4f737e0fdab49636d8971bd56fc69c79e1f8ee3fca69e7890a1bbf1039beb9fdadb09611aaba19fb3118788e9098a66c126f5db0a811c0f8a90eb03780b42173de561f3a73d592825f3013ad1f4d73a00ee41857520cffaee793e2e0ddd65aed74e5270806b4c37b9c8cbb867af9a71883493d6b17607fe5e4082978345826c0d01671ffdaa5a3460918daa2eed373d707185aa2446e002f991f6a533291d5d4649c84468d5545d5fd606255468256ce7020cf2e8a4eff76b554d39674c97e4371f22396859e904512744ab951092ee552a85878e69981e45899efd13fc1ce188672e4cd10ecf7183c9dbe9e8c6914cf3270be03980ca4d7bed28b2754497256a57b1dec3d530e388905d6a522fbbfdbb3848c615be301ccecd9c51ec7f4432e0ad676202d470c097b145d86b997f6487266395e29e1588a898ffa70fbdccd882fc2da1c3af0059a7c4721cc624e5752e7c84fab8a6d9f9def4ed1b1fe1989582b19e263a9d8791b0f4bc5a5d591c1166c5edae8e2408ee31bce0f6e34d4a8799f451a85fed221d05328c35648aea692d48077e124e8a3df59570cc0c26abe1d71cf927547e475316861f8b16b3f4e085b5a8ccf299a085810acc05e8f5316930e2d0400acd9d30d707b1ee739a3547e2bab747e7881af4ab33efa5e8f7af178eb8a26c76a203573e43a2d08fb800d84cf4b2c8a7d2ba463619780c0d4fff07c5261288b4fc7cab51257f1efbd3de838bdc25d8d236b0f250113241cef1e77690a4dfd06ce1400ea481fe2f45c117fe4b9d098e9edb501432ad4d6bd512078dd1272477c848f1990e2d70e81d58ca45aff2a9d593f3343f8c84e1e897311e4f2760dbbd1b66f838e688472d22dd3ce68d73e7b33796b14faf215aa4e4f4faee9abaaf1d2d1119d30301f3efdb0d40605edae2ad8f58da2746a92bd82a4cf64;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he1792121c2731fea4fee38f41461670cbbfd4d897f011a183c278728014b9c2290241ab8fafc0f84d1d84ef528d1b682daf27e2a5ede521d9f8d6227e97cb9a1fec58ffe9b69a49d2b2d4400aedd7f37b38dde8e8b68fa4ab04d0cd6a7344d638f3eb8e92f286e4f646d0bc5ae780fee3462f3c06990645302921402ae78d47510124e00390022a05cafaab0579f3c271d547267d6cba07ac5fec2fe616210ecd075111c755af9b453101c25331f14c644c8dc4d091a35f151f3ed29b85a6ac9f953b19a72302b3f754187ff8edfb39953523a5e204f188cdfb47dc78db13e651d5d636d8c0273f086c45457a27ed419d0ad232778b61f104ed5f9249f8d68818553ce50f9b04eff5cf6473c1bd27c8266b0e5e3a2e0ac3ad5705690589ce5dd4010881650f3e8bb39e6e5f296cbac50922fd627ab878645155e32c7e192bee62ac052f873cfebc17074a58625606afb8ad85121f662032ddd268d87b91808d715bde7cc6441592cad4899ac3c128c7dbe854c545aaf046292e126b8aae49e42248dae5cee5676657ee7054be001742dc4e8792c62dae616a5eaaa3c27fb4b48a912e815e15c6a10b2703804ee8eb0c04146d14f5f45e611cff085542c21a11f4dea8dc9267348d4e4e7a2131dffc570b4d4c63d209d3f0e3058f33965853f02986573ac31ff716fad9dc1a9c69d362b54c09afadf926af5b9e95c0e287b661ccce2341d2acc906b93419bbb64f21dacd7d3257d95bbdefff45544784ff9317c74a8df6b4fb9c85d65fbe3b6c4f7b7a7e26b6536a32bb46b63eecc29c0bfff855f2be0c2e0b3d4600d5990aea234a080b2c052a04aefddede4f26e95be57f447067eefe327f6661bbfd7c70df7f491e30323e7a882f515399dc7032e667e090545de461d7f153263c5cc473daa83cc1efa72936cfc4324a3fc8b24fcac6d3aad8ae8b5c6cdf6171b18bc29eafeeedcfb77582feabba417da88338aad9ebf37d0b32bd96995df0119d0c39859ee644c3354017b0292b1542892ce68cadc47126adbe9fe6ecca8b81d64b1418afb3ec10c6c20eda1bb98e09f92d82d53b8eae207bd1c40294c64c710cb7af0713075df389b1ba1ff49b6d34127e8394a63250a839c19a32fe1d9a0d2ada1c801f2f606b68e44c0d01c6a35b9a5b604a2d115b85a434859d73fb2432903f0d1c2accac4f0d80b9c4869fb3a36bcb918d847a2673c8ec913ab80fc6e891367c1bb283d1d31af8d4e07159a6718d21b2d06a7c19a8e15aef17e0243adfa2537b8f14e9d1554913482ed3229a042bf2a846b7b8555fc1bfc2fadaf91f99406dd429f6820696cce0eaf6eafdf6827c5fb96d607280545f139b780e609a737212d742a5e228b7e3f18a5e6edb796e06d301e5ad24ae07ecec792cf8f16b36298415e0c03a59fde68c0adfbb5185941ca378c34a8be081e726ea1cacc3c3c3401956058fbeb7b193c3dfe7b1337e71bebaa1797cec15c2f4c13efcd91c3849c43efaddde11199466f8efa1f48d21cae8c79abf03b17d3724a171b063716488af4205c96e99c2176b06f8af273b77a6d1773b1b17e691a8ea2adc9c6a7ec9c237559bb96933c1708ac5d55eb5690b3a0e12e0e9be4f0f7e99f69ab8d21953a2ab8845adfcc648658ecbfb63d3f27e3bb9a6c20bad9a73843b247818103795ad9246c0e534de8bd3ec14d5f7b5f398f80e0715a3a0285c7f8342832e283f1123fb38ce3f0e68ea313fa8e992b046f5b9679ac7bdd7a96301f825569fd05ed5db263a070f196f05c8795a49e0d1b0a84c5ed2bc507d7e635de30acc1ecb066c5ed6b39bc950b375b51f1e184ead1d0b62b873f08af5199265c6b256e86cb67d39aa175d62e480c3ef807504e97326d45296621ae872cdd64a05f4ae45944923010124069d47af122bcf1e3871ed7d57a4fb1b792807812df86d83c514b56142921cbe3d2f4310cb7d5922e9e19340d20a5f336c7f704bbb1e0508bdbbd266b07efc3c6baeb10542784602116262323e27bf69a96c20449a7301919164f6f3bb31fd0e57a220a4013cd877f908ee1d4e6c3ea0af19bd3c1cdc0aaae181fe87a707d85848e00b6fbf87a711f7d8cb3091b4554eb0a1a532b1e5ea4ed354751c818c35e36849eb361300f7af7e1bb13e1074619e9b8da8c23780a4ddf43f1487d739443daa58004ad39171b70212075f3f76f5a367565d072d504f648a26f92d1fdd3701ac7e2ac799a4373cceef2d8f80f6f5de94ec7789d47d0904ff244bdf96c96a281657ebe9b5c2b6acb044a93a3ddd9b900619845fd22dcfca3f5ddc7f507645acc833f16d30d56e2a03ab95516f9d364b367189a42d65043109cb6e928bd6157e8280d8fc4786f217a89e975241d2baf10bbbe526cd7b874ca4284b512acfebbeefc3447a48c1d103c7f1e8f0bf7e23dd4e43b6f2ae66b80691b8112251fd2fa93742ca4aa8fb78dcb395dd52bd6d0d1feddc990ffdd35294cfdb826a1400b83483a959a77d4cb6fd36ad39cc5b9adff3a7709fedcec44a3f4276de03a9061093a912d760831c52252e31b4afcd8cd183f839fd5aee6878415129b731b9390c94cf4b798485c83979919b543e609ee23faad63d361ec230a263c33a34659b2104016d57b8c01da8dcdb814de6b040c1309fbcd2422c83bfb0a5b07f422e33b786cac821370cc26994b6f1c4693a185fc6f0c2ba85e349e7c0ad51fcbd6ce810d5a907bce7cb36a03e614fdbc513c9456afeee00fdeaeadea3b4c4d156ceae8b4a4d36bf5725874850e5f33339e93a3fbdc32d61a1be29f92b0f29ba283a70a839e0f1176756a1143aca621751d6d57f92c6be0f8945702eae5767a881feb03ae3eac3c5e3fda94be84f4c8bb23b1fe36408f8f3305013a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4545783ec4d2cc4eb44caa4fe7567ef4bae790f80d24603684b8d67b88be6f35756838eadd54607facca80f6d15aa764e3feb7bcde83c470d18eb0377cfb3635ae94d1f27fac4bf70e463b1388e92f2078a0ed58c8b0cc1798f2a91ea8f37f5f3eeec3bbf172451b201661acd14bc00735081c5a65f0d465a71bcc91adf0a35b4700191ac3bd31d11ea242edb04d6086acf6a2d3ca38dd0696331395d9d47a462f8436f21894d80d274140978fb0f33d7120176aa5b895a135cd4c3f6ef5d1445de7da284cfe72a04185b1cd8ee5a32ee28dc1bcac6d054dae64d55ab10e83a834595aeebc0c557d835dcfbf5a1a8843e76c38e7337d32a7a2f9af8f8bb3ef2879d9cb03ba1d157f04fad7d9f3d93a8c4ccf89ed2c2471339215fea3ea45137fb3e9ec204805927e951cdb0272357498c81e66581fa6d4190e746c6926162f6480545b2b5e9bea4ffe6c7d4de7cb30c21009c4e80592c7d536805a14571d559ba7929a9f82f10051421ee38b2f62280f775a8f9b3f087ef2d305ff380d4c6bb46b28e401d3e8a1f05282da91d629837ed08e6093208f1ef882e2945041437e3e931119192e70c0401673c4ed8afda3b09b06410d4bebaea0ba024065871195704c1682ad1154fb311e0bb76b0364ded1b19365ba7df286a275a28a48df43efbe0ecb8d347dbf6f4275272b0a443da1dacfeac3b61e10f5f06e2f133f961e3ffdd9ee495c7d1bb266c28314e11e86e9da57af9357bcc72906e298e00dfcd4ecf496a58ddfaf5fc774e7e26ab89efccb43229e6382aafd31ae5952a49f5828eb59953c7e95c96e40525aaa47e97c1848b37e01fe6bcc6f23f825382da05ba98f9cfd0d7d6d7d4955b59b56069e877399a43ab91fa6b16c5db1e5eaaee53d4a2252f1b1452757118aab0d968a5dbfded524ab2c44823a4611d4cea7fbe422a2391ecd6651241e8dacd16d386fab9a6883315e2ee2f1d44582d77e1285c820ea7308ac1e36c0450fd9cbaae5bd20627cb06a6fc43bf04e92c30b4e4eea37cbd1b65725a153ec347a33d7912da4d938119685c21073f10e6fe6d0dd122660991ad51b5fa895aa66ed86c778f11fe5d8d89fc2b39f57601db52e44accf2809e4644a23db3ff747922c80408ce7cb68c186af91dbc220a8ad53deaa49c1945bb89594a2841d94c1ea5ae524628a57b7f3a048a0e92ed7574a07887d9a4ad660e8caeb9bc4351dd48d9c54385edc6ef6bc30cb8fa6fc51e664661f2d3da6ecc27c10cb703aee3c381db0b36ca697b66c2fa511d259bd1bde9377e01863687a16397e350b4532b2f4b7e8ef2b887f4998f9b0d8c296590c04695a8341e33b517432734738b563e907ed2b5d32a2b44b6e8ce2a81c204bea8fdaae64fbec069a3ebfe5aeb5fc75e76e4a24c0e6f727046b5f58cb695cf6dfbbbef5c23de95eba5229e8034f055f2b831e1af04e9570be22ed336d7f8620afe3c88fcce2ea304476c3460cc3da11bc4a864d2c82d05cca0fd2d2bf7ac5e6a37127c92a8b54375ee681da36610125ef0986eccb47c4b60016c1d95ac83d35421ff32d3b1b4b1c6d037aad185a0e7e265fc85433672cc165c230eba3ad0f4f9cf6c1931cfb15bf455063868a369125eed87ec759d77c37a29058d5ca1987007a8eb7bf491993687c5ec88b93c1277e20b0dbd08e1a53ab710f8f972c0a16f26bbe5370fe9af71e7d893f25de45387c2787f57c21bf21f475e0e0131e883ed66c4b2b2ef36307d142801ef27a88b8896841622e35aa05776897785a99357d2ba60277b5d1fc260a1a4eac3de5ffe736a071750fd75a7306b0fe368f6106b81558c0eaba64143adc5a284c9cb7c1ffbffb1cd69291a05ca92c2907a70f06f39b2c198e035ebd22735601c3d238403fb875abb67a5dc0de09af8954a96842cb4e9cc175ee2791f4af6d162302218941d016135cb72e1490451a1bd24372cf7772ad3fcc9f454d8dc1669dd603f911da11a442e83cb0c4b855e1879283e053a9e684de044491370612f8ac913324808c0156cccaa1625ac91ba348c670dee19df398a9cafb398848bebf40e2a9ea810950bb1e70ed709ca0721bc5d53668c2ec3aa1162bbca40db95812be5859bfeaf3fd03648a13a3d04b60da8cee471241a05690fd455a0a70cc03620e21ad8e70a98ccb888e3f6ca7a14af3d6c14161a5d2dadd8be2e0a0c8660b657f80cece7c28967ca86c8fcd132c467cae9366a5d26b23a379f2d814ecef8ab0a5a2923ebeecb2c4c9c384fd9a838b09d235aaea8c6868a0b882b191974e78c6c5cf74c16a9b98dca9a660877cfa2385db798f6fb7e1fc5c6a76a80fb0c271f197d4b1f0b43fb8ac8754a6fb99047afaad5f5ef84da714f41cd0d75218a1d7dd69da3f4e417a6456e8d18fd1d4b7e0f2c43613461e329993b062df0c525e4a3646301c0a13f2fa4c5419af51bbc9763d50622363281270f2fdee1896f9618bb0996751c66cea3369be117bd92c5b57b39319bf334fa81cc8c543983709f86b5af88ebf4d462999d3a6add34af72dd7c2115c104a8933a14ae34a75611865695efbb1864672f10d66862e72ed639965031932fdbc7895b632b4d7783cfb0e81d25cc4863cfc8b8383bcf4fa2d4d540ea1f40999226d44304bda94b131a93ed7eba25646b681473fc35e60cae2d31d3daad39c0426896affc608002444a687dce82909559c5786c8b1dc995d0abab5dab3d140fc3b27dccc7063a70553acea5ba41d26d0a82fef7b5efd704782ce62abfebbc7e67ca73e6fa2c0df2d5aed79189f90359e676ff71e851503b7f505a957d01d3854c34c8db8f1daf7b08514210847b0d2aaab8a86eb623de79128de752d1f3afb5a87abf14edce4fbe242b4ea77d53058c19de7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h20257d37cd3db4678bb0c8af4daf3b27a1f3034a3cedec3a4f1dfd3140e1feac84c94533796a76669071ae77c02fb811158cd20797dda00f7431530fb6d1e8c7dffc64763dececa13d3b90bed000f92d021f7035ca1fe02c42daa12968336c209ba23dfca56dd6d6bb83132e9dc885755c55bee86585bd2c332425ed9e257c1a3893408bc7daaef3ea7623f51add70a1f1ecdff2d4edacf3ec9f11d96ab45a209be1109f4086167116a04eaf58be3ba04892083ac464f9e879319b0f7d90c23d858363749421fcd760340fc3d41d6e0ed4404c7fd0c0adfbbfce407127c16265bc58129ae6037e8261402342a6725952595dc8b2f69141c7ec30559ddac1d1695eb5e7c0edc7b0ec9c463f5b159c440b06066d7ad7a3c97bbdd82dd618c9a4019304acb1145637f048fdafd589f8c04724e161293f83ae6e58b0c100d90cbbeba06dcceaa6a64e3525f1cb3b30bcbd74fa53dc60573bea13321c5c7f5f633725b8d64463bc2d4896619f048058e2030579ae4c0f8f6f308ca7bca915230706a5e04c36efc112bc1808afe5e218e0ae4bc92585d455156bd2433e704c8c713d59dd127d4bae72c96706094e8e3a2acc55ada09969fb1067189c7000d386629f344ce02133b60119cbada2f28442a64bdd0ece1eeb6bca6a9efc78afc347f35fc0a99baf8ecfe4eb8b0c813a9b32d9260e24e17e581b261f078c678684536ef7a9d5fea3e179da9a70ca12a909399f796ae05e524bf440180c6f0a9251ded6b3ca1c3059daa0b1b0f928789cc26618049d5f9135cbc1a9d505f5246b726b7c1d422f012305f2d29100f2ea5849ca6dfdac30a7b88d2d33655564b3844a36657fecfd9a97047d06cc307033f323f6d183da5da2d33413e9cbc7e327f23d1d27d6ec0035691783c357f746e7ca9b01b93197b5ae27dfe985edffa0c65c872e287bad5eca211713659d35141327e7760aad8857af9b19a119b4324bc02f48f54cdbfaa90bcf3c8d5a22e64de35e59ba5caea8c08837baa65ddb675bd8e31d744465d794b3c9023f80fb38bb73b119eb6ad3d1307e9e0fdbbb5384c25defc6a587f701748ac3557251685393383066def8f6b177e29fea9ce88e7454eae1d23be7bf966074fba5c41983d59ef828bab31ed2bc7080e12039f066b5b397d427369b09307f4153d7769acc4030a3fbc44b517556165497fdf0c8ccc6bdb0d1ff049befe051c26d9c460f725781743a9dcf44b5d8a28b84ba57518109ac3718c2ade57408152dd32ed31a57819296dde6c408bf47aa378fb6a7bc3631653617b3f97ed55d7a65929c7d3320d5e85838a4dab8513f9e30ba072a50b3755eeedbbe92508d5866ce51612ceaf956ebec9bb27e5ce54485b2064201901c8e3db08998195901cd14ba9c78810faacbe385e016d6239f401a8815c60e2122b456bd4939bba32bfc476b2ba0dee0424ec7da56e46d6dc9181ca89246cf8673e4f2ea53e81ee669188adcdde574c79ffa79fc1b0a269bc17fbea26d8af87fdd8fff61aee451e92e81d57b3d9381656d9e174698fdee2ca2d9f506b21e2eaed00013e6e98789ba86d499f9d61cf95256b2faeefe8542a8f840f330dbdc477626b1b1cd00cd2df0f6ab687aa92173d35458d7b2785611807d621464ff9d8c3db12fb499a80ecde70547a0929d8d172a372aba51ed30b03764e68d610e65990e17ebd767d8c4c3b4697cce1e8b40bf2271573cd300f9ee6d9ef86319a6fdc40da264beed0c5e5790f6f522df0bd93dbf76dd3ea3d381a6e25bba5ed4d07c941f6c6d03bc577747ec56be913a04e1a94660ce8263a98317d4e0dcbd8caaf5c56fa8b8269c77c4cdefc62c7fdd4b4430818a6476e5f382c4fb3fc8d31023e209aa1a03f03e65f6985b0dbe2d502009b297d64f9f43422fbceb2424923467fc03a215ccc25e31e35c984093bf46fe609c1fa80ba94e42048f0ea64da5dcb9af2d13da6a0fae89325e2d94e8d620a3d8d4aab5b7aeab34da8a8d6c602ddf96ea5b465ab35c9ecf16507c1f62c59218ea9c2d8fdfa8159352fc5189d439f5d247a6b3bac0a1fcb0da18f8d0407a529864350bcbf3f29b78b2081f4b80ebae2bcc4a6503499a7f3705c0709487b7f1117569d1f8e7ac2f63178ae48926c063f9e005681a927b769732feb280fc6cc43522e9eb6cc3b9df122e7b4b5fb451fb4db208d8abfdef5f971983b68b4ded99a16eba9d7d71d4156783df674f9e351f0b93f0947c2695fb1c046a36cacf14ab0b5584436f33f5f59d120b86bf09255c544cf9f0471c7071f3d9fd83763fcf042627d8946aa096e107cc32b33889af0d572aa3800f1b384657a47d1266e65d04795504f6e9ed894c989091dccba7f55d151f58afa70694e3070e1a2fff17cbcffcb2fb64864e01faa5c5f11ef60ca0f7e974e06b79a66e939b0f794ef27f75255ed1973784e21b6fc0056b62fb70aa8a203cb4affb19e4789fd06228f13d5dab8dc5a68b7d13f520d053604e9b398f87fe8f3577e924e8acef20a18d793ab5f6f25e4c17b575d46bb9b554a36943cddbac22dc41c231a6775f3e014949ac816d0c789c777a6abeec3405ea20e69a08205975d2e90cfb5f7580900d5801584cbc3c219f087e3fe2c732c8a5804f4d3ee2ca956222946beb9f40d8d549447c8405c352e788e185308d9f62959e5dec6eb0f50b7c33d9548788ca9a1fe49d9a73a9e261fdc3e94c6d11d64b82c735bc864340faf51056734d687e8a57a21861fc71c557bccedc241f620688eedd37d84063ee642b6cd4a3c9376f3ed42d0603577dc3ee9447051044876fc9c4a3d0e2ab58559527d8bcefa63e8a002ebf5d7b4aa4e9f12ab32b4567eced7914dc8322c041cb58241cf33f615b17a4e5797d18;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h692d6eb72cba92e401f059fedb2c1e7d9f7f2535477f77578896d65d0b934e573b87bb5cbfe7c8221d5850f86862392a4913267d7b9f939d83ee6e2dc723ccbb6575b84e183f21f01521727ead77eec816dc48e7bf3bd19e8cb359521ea2602a71426747f1ef548ef2bf193d3f3ebf8d1698625cb43adb00463a58f34723950a2e4f1d3f391685e7f8f23e0172142be4da0b79b4e15f13f561e7191bb2e81de2c18c8fbc71ae45d6fcbe35ac2cc28d43d262bdb942e28120cabfbabfbb93326d3696ed554f9f7d9561e7942a8e4c1502615ebbccef7247f40cbee0cdec19bbc46510709fa49944dead31875387be574d8249fb83076e7320924d8f878245b72b32d012b8bbb787b117c862ad2fa79c349f6c30ce92096594efc6d001f3c288d6e310b00bc305ff1b33bb8558d5848eb02f7a399bf26f03fd72671da4141878c211e20d53f6d0e3f3cdeec10da7c0c82ab92f42441bbd73b4e8da913ff59093976d85a4d34f8050e735761ef7f4002ee2383d1a56429682a5d224d6401f07d0e990111d3348ca9ca164f113ef7548cfc00c6ab56c7a05e42095f760dd667257267a84de887c414efda51db8fd39113f8d3e29f0002d07a0c7233c5d260cfca22fd795ab31575bb372b672c7c700c9323e5ba2cf5b7c2b34a2e55e2ebbd787faf3039e4049fee3d13e17ae6ff95c02b956d966e9344cadc60fbd2b60a401aeeb6eddccfd1cbc16b13f7e81b72c048f37fa83dcb90e4d8d57ff1b8a9a9217a24bacab767593840e88c23b83a6e675ecb7140209b4c0111fdf913ae64fe81b5f1371b9c169310ba312dd1fe24d7ebfad3fba4e4c8e15334c5e745c73825af3bea22c264665a4b9df107c50bd5bdc0efeeb91da79b604f7be2d3a17775dbb220ced8e34a49329484d74599569fb156baa3deefcaae48b8c38b1654933a9df4949aceab1e5962e1750d34e692af754df2770dc02b32864ed788077c3703aca26feb585fdb239a8df48ae1992a79d2d68658c3e758db565c9cc3bb6d2914cb4eec13a8430c2e1b2faab6ebdf1ce3c3e5092a6d32361e624563ebf5f58cd188392ceca7e4dee380bbdb2343020c3fd2d49f37161581f7dccd0005b706479f8c954c88056dcaca9bf3bba007e3d6bac6473302b3a04a926467b9d4159be77546502f925fc09a8c61bafd7296eea56d7dcb2df0750736152931ae7e4861fcf219ac7ecbe062971b8d905daf6b44d5eb108db90f1f4ea0ddb48edf2150286187683918de39f3c713ad65ed3ebd9104cad0cbce3ccaa998f1cb638d06e737de34862e1252f55662cdaf07477b3c94370a810342130d2dc817ae58a921ab785ee72f0cba20385525af5f9cf194be9754b9d463354ef01a8e3f5b7fd0b26bbf9e46d263bc99a6da1e2d9a7bd037510e118dd03cd9e9d30c6792694b1c8130b0cfebf1e09b11bf8a560b51bd83c12eca801f0fc3c0ecb3b121a1ce300ce50659c7dfeed8b159603989152945eb230d5baf78ca9a0a1d58d6d91c6a3f90ead38577a531c14901252e9e96d557bd3e1caaad769abcb820a6a6095d7c5e03c9118a16cc48922d70e3fde8a8f3640dedb8f0609da46aa9e54a71353adb6326a67de5d88017f1ea8550a318b261c674c493e657188958799987fa39e2fe6b4b0e54ccfbec8ea248005ac99520a9dc429687f75e06c2647336e7f91d333045d86b40931d72c811d48abb517affb81076b98a68815b5f4e47d7e950636fdb36e44bb1cb206b3b159148d5753a860f63b50351d0d87a8b55470e8dae282dad079401026c440ef5b804a72c9cef7e240ebc133f017cdf6ff8f18d610bde5d368608d407a1e53113c4b2df30267c53011f862ffc58e132844179d6b0ef9cfa97d43c811f7412430238a36352e5a95de67444043bc50c6bf46b76f7b285138b45b595afb366112bf62240bdcd0151c588de62645717f2eaab6acf2516d68a6c1ae04385917e4a299bbeb3ec87b0dc5a1dd7aee8a19b18cc3d60e8f5bc72fba657beb9757c9efdcb851401aa91ba0fd050af69afbc1cb184a77172cf1b693599f53a0a64c4da2f16797830bb0726a94241719a3178b7142d46814f0c9b670ffcb806899d11d26b05e867fe2203e0c9a8860790e98b3ff637510bae521a528160b1e33a5683306c2ed72d992c90416fa300e1afe7748e7bf492ac6aeff7c64d7fec2f17f77365763c5ff82aafc9dafdf74fcdc4fbeefc3537e30dde9a612b2c651bfd931eeaa4efa8c1143ae80f50c6ef4c7c4dc0ca9cf5b181354bc7d7dbce79dd99f6faa003db0c154bab2ccf700c9a0bff837cf16abf7ead9cfae54fdfc022cc1980734d8b7206b060c40653e7b48ddfe98fd06189e666cc9f76d502c86c1872d29906793ac0ab7d9aed596d8d646f0901d83156a6728e9945864957654c9db236a5ab4d68509c6ed8b52c3ecdca3845e179a98f30fbb0fd090cd7ac7232858b3bb2ada14f58b360abe3114c37f25e722cac3e6db4f9108286c75ae69c4c8499b9d5bf6d98ff936cc268ee6fcfae77f750bd117e21bcaf57a574f85ec04dbd5c64e640f21a46a0f7d5d4417f2526ab4d27362c3738475759302194b0e3a06c6cfd5d07c69231266d1367e94f84153de499d1408a2ecd2ab4eb69448aff3e828ed1277dba10c8ca5f9e8afe35548a069390c8cdbf2dcb09d021f03b647d4bdc2c8bf22bfca53975bd8720ca2e249f0c665937a7a62b749a4f03795d4b427a28efd19bca3eb601f33273fcab09d9cad4737b4e440d1071349eab75ab52b4b51b669ab2516d9348ad047908e8da39733a6b87152172384899ef93b9144fc5bb33733b87c8b81505c5ec8d1738499cfdfb69a0fa5e79440f9129150619e227f9fe98f8e70e01522227faa40a7e4c1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h264e0ce204627b4fe00151a1fdbfa023c43b5358986a60e072674bfe4e53551655c16ad96feaf0f4ee7c04555bee9c5d6cea2d55b3c4f260bef7958fa6b46ff88ecc0b2130f358ce930fe28b09c9e842e2e5f4052f598b084f82e159e7ffd89aa1f1569be0ab604d270874c13e27036968f474da7502eae34df28a9cc72ddffe9ad7c5dc445758b01ebb9b1b1763f05e328d2b6f2d7c7e7e572bd99c313b5f46218f4f974e97ebc9197a1be1762044534b686a3e3dd9ec4140faa604a6986e0d0b9d0813be9b294766c4e987d03fce009a53af6763b4a1050d805f93254443d2305e6d856e1426cf98b2ae8201794468ff9c9598e2cf74a52df5ca20ddd4dbecc60ef986820142c793f37a84678a510aee56f3a10c6a0832d27287c0b22c495f4b36bbf212c16eee421d58f7f4db9d07aae6a10c43cbe4d125b93c128b5ff3303adb3724f3ea510a0312c5c5cf71c66b870368894b976c5d129af637ff92e42f01c50f98cc01d129a921fcb7f7f11e19045684c1e65d308f87c335f20a1e0bd51f27131413c94c2e7851e34e1813282afb772e6b6de2d535daec1e0353ab70e87514f55c1bb568a524354a3c7ce5c0bcfc2e49d8b73c95443bba9a3502b2786ea9d2d395e48f88b2ae0ba4faeeac963731cc72988b68317ff41ccb1e9e6a68052fb76447d689dbff16869feb0a8c8b6250fb91cab7a0b2908d18764a8b6a1a0118ef601b820bfe391c14c851357e3f8c391e73403599329ec41140a40a986cde941feb6f0cf591187ae30219616ddf2217934589379257a7341795e34e9e87511e6206cdf3f3f22e252194fb1f0841425cd762c71fd7729ae11fede95b535f6199be6ae2d1ad90d6f0d6f932f679b44b9788e57302cb7f486091941cc1bafa9670b1585ebb6f63244086e889b7a69af0010b57a66b7f870f33febeadbd165a727a083893ad2580bbc07821d91394a59035e3c3f328f9793da4c680319b20aee7812207f8540b5d63e3a8efef4b55e66b70f2674c61adae7cf10bee66e37b49c91fbd5c498d7272eaa570ecc159b1183dacdb3fd8698b2a42272fba223cbb011a758a48493edfd9195613dac40e4fc2b58d745cb49c0aadd4a7a0ed172e3d899446e4817de3301b5bc2a4f566d6d64f93b0d215553062aa9b5756e0677e58a4eb41b4b3b8d5fcb356dc7e9d9f9e08e4f598ee9132b210d0f847055e11845218e4e48e2851fb3ed12577588521e4b4c584e8e774551b2edac1374c12b129b1aae3febe017ba110bca018bdc3581de870bf81af9bfd53dc873cda8b53bc637bee2cbb982553c2ff9288ccfc886989df2f2808489f5cd5c5d62583c3a9dcc174e2f2a0bd615cc57848d3f7d3d8337cbae9cb0a8f42938a156d73eabb464ac1b609977bba111ca762cbdd7b83ad82df05ce574876a9111d68047e703dc10606416fbd6418571b4c9e4066e5654f07a8289d8b2e09a174ea5b75c32ab08f391600f3c647290dca6ec92dee817b868c0fc80a6c111d76c3bc49fcbec98a013573d74a61b75db377ac9279d306e25b3988fd9d78ab23eaa6042b6b758cdeafd4221b8adb38e0e5526ed8b79cd2bfda905796383738391551aaa09fa45f9d1c1c89696e63404e4f86381e6b3e2fcd07f7b0f9e4b04c9023fecf048a92e06c6cd6599663932d29e2b19c48948438e13e4e01ffc401ef3349419929ad32e5dcc1c4cc9889f57947aec91e912defb0de9cb82e1c4c04ad1e2091d36bb86347b869be3ecfd93444e3bb4e27f0cb019c1b423c793b61c566d33d66d56089ed3b9a0e4bdb99fa64d72f8fe1e496e791d2b7ffa0cd2d3323de6a682e5c366166b783530ad569f641d066366751817e7492359c50ae6b68f797445127401b5e7c4ac8c6568e7431a1acc8b431a8ec1ec5e0844a5ca4484f783cdbf510134b61cf3bf9b15d7a0a846f6fd59d1910ebaf4006434fecca0d676dc61e1154616b4a240cbfbdcdc9c70faa1dce726630f47bda87fd21ed547fcf73fcd4553190d0e2174cb9b42ae98157245f3e2cdd26bbd609362c660644a0832f28cb82d1e150dc9318edad23aba1bc2ed1a20cc0d8fcb0955cf3357fb8308c400214279d167c3384a27664acc2d8953a136c1fa86781f93cae768aca15510ce9f9e9a46dcc25b51fc62302e8efc9fa20c1172d64c795d7b7eb561019c5e466eadb6a2d1e53332e33a4b02c2a482274aa504cb506edb616cf25774d21406fa1aa3cbe071870aa74a73ee272581fe455901bbb9fa49a850390618ef4ee1264d82e63e88482473d9b3c985536d493d5126862f0e36ef9cb5adf5886ce4fc0c97756cf014530e973f9e582aaff01c9e19ef01f7311acefd58aedb0d82bb628dcf2663530945174a9e096b5557dcd367ae5cf585c5f8401db625faf812db403de46e2114bfb85706de6da2d5c3cd5848eb8a89786594832ab94205bb7b72b53693da3b4b243e1bf0fe5b45ee2104f41aecaada9460c0f2f4e4b02af128a582a1fb8a13cb04062181fa749198f1a2dd2548f19af458da605dd415b7e4cdede9864107851ebc38ff9bd2ff9eee14c2b23a44e4d6f00eafb84bde4326a6cc2d925f818d800a1e93f6b18fff5796a1179adf54484fca5005c6fdc6b91d16eeeb84c280ef087f5d9637b200359c215a4b186c98e51a95e05da4e46883671790f7b69053de0e9d8e1bdef7da62e063e77a31e5359c9384c9f00509a55adc18b757de9bd6e6ea3104a948e5166135c1170b4921ee66d8ef6ff64188df0e010227b136529665fc85cbf6112426328924c873c8c91118d163414af85caa32192f6218ddf693ad20f7ea3d1a52b05138ae02d8d5d4d7e1fd13cf9d2f1f7cbec0db9898e93b80e573a6ae16bde0dc3b0e8b17b49fcac6f4f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5a8f83a195b2930cf7cbc06dd2c121e6c03442157e6f7d238621e4bea7363d8013ace6fb3ce2c3e9c7b5cf77f3d49e062e4d3ea4ff98a1ef3605fe9523d1a6b394e23ccc1aa760b842ddaa4e2d76db6b77ee23fdd566cff576eb5096838de830eb7fc5d6da8497d7ea7ba41ac905225ac4ee31ca737c2165b6fd017f07c01bac0cb609a25ac8a1b12b34e1ea9530eecbafe8e4f620e714fb2db29e6be44e847c1fd04620c5b1109121e1d02910cd44fc9b28f79f04ed5c0666d6e58df249642fb22988cd73adc8a0f1ca8025813e44a21d87963b7532f5dd8e17d13b05518aa46dbb0bafa926c98dca4ee0775c0a92d1fad928c462251a22706675a427affb90ac6a52f1784786ee538c9b6bcf94820053c72c84ec069e7dbb598e8fd777f410823b7052aea8ec2d7debb28721ab3792d073eafc69d99d0a82285a407702031d7f1f5768d293fa8efcbad47616f890409ed48ee571c7916469a3e41d277677d866e208f0f9ca013caf24bad46e5006dda578befc06ddd2d04d1d8e34a0056a58f09cb39ac4327cc7c3d15ae3bb34f102d1cdb4ed6f87441e2afb344202311df980f1f1824979f152e3fdfbfe0f5ca538a696ffd818881fa79371896a7a7ec25b7a308c0ad516a9d7918e67fae8a79e73d2847bdbad7b365b531537a3b6de8ab03eb3e63275c06775f92d2e52c7bb947be36799a523a4caaff8098271c1536b7931007e042e6b78a9025ecf47719bc459554796a458fefb678026a311bc8f286bf2dd4bf57839abddc2de41b9e9756ea8b17b52271959680a29d8ac60e87bc2c50916923c4ab9b92686d0a738e7019fa849b7bde8398ec98d08fa459c7886e67a8816c7362e652e759b8cae325f904365a725d9203aad8aa9784bec23f800ee714f7c1159b0ca1111ed36abd20a615af41d75e679e45fbe9f3f30cc581fea0f1142619c634253581851dd8dd56c7797d15ec27f6e43f0f156f9a05aa98147744d2b7b473866b68cc4c1f78c60c04aedf6142bd5a0df312e4c95d0332deda7e924027ee616af199e9c7cfa18c68afcf0846323f5944037badb2ad147c37144afda52efef93b17e0f20ca6a56b500b41963c5b45d2e7c295ecbe104faa5e5863518d63e1fafaa7e248947346e80f467dd9a5095bede0c35ce757307a55638b60f6dc225eea625c8374cac5d4f20cbff8a91ad10346dfc8a4a0963d80bc847239e0070fe3b5688b69f8f5df9c4b833645211f9f1967dbad72227f40f98a0b4b34f7174424a8393d03901740db59c989eed88d7018f4116b8dc811f028e1ec7000d2df0266d7f09bde0ec7a349f1b4d197b530320ae163f842e2e08bf62b2d07b89c5fa436170b0ed60d5a8b0429ee37f4aad5dfc79c3f9adeacb1632e36ef94ce7b6f2a21ee492af36c4697731721fc0fd60334953d10759b52f1e46f7d8783598eca9e6883fd82a56f547cb164f4e66ece59ec53200da98a86b8d90ee43b4a9b576d3d4fe3e74354e73cb644cc133011b0a1dafcf0c501a3e18221e975642a2c2be52ded820a90eb273b95560dcbcd8942499feab4855c6179fa37eb70db446e81f7cc21d24dea4c2ac64effd6a9d37af6cb2ff4d6905c931973ec6231b8c13b91cb045d6093a4580a95b9b3ddc42ab7dc177ace8c3913601543813239168adfdd513e9765924bec8ce524bfedda8079acf71d006b814566cbb55ff6fdc4f493ff58a1f16931fbcced28947ac9c1a00cf9bf5deac0e0f287f8e1b5e51fef2f8f7072d86fa2ede2bae4b74ac13c5fc6f51ec943f2ac5834fc8ac65a5502b2c7baf9ba16dcfaf1e792b544e6bd70b64fb80da75bea51310066abc45faa5e5cbff1268e071aed11a3c03b73799a6e4cd5d3101127952237c7e882797098c58d475b2db195fbc8f6c9908a6188c612b1bdcc3401c8f4a36f86657ea1ea105c91b2003806929b8a4291d916ac9e759126a2b041b90b199d06959979c793947003776a48a600bfc62844e8247b61b0748c24acf406417dfe8284e1dbaab1c8f7ea0e0dda7e432b666d2f51bbd55e2c84bc423c138af1cfe6900f50a4a7665192ee852c55c1a9cf1b07648a702ec595e16802a3eb77d0dffd4a4dbadf4c2511a55c1c7e412d19ae80808a1ad719abbd9562b43e869b71c62884385c379056e0ebde34c2fd3e3a908ee477baee4552d45ecf7f38658dc8c844a4e1db10112dd68600db6cf492ac5f613f15806754b3092d848ccc079207461b66fdfaf600379d2872c7ab91f9ecda4700be39e567b365157454450c31a93ccd81367d24e5c5e416691ce73dbef9132ea5c73f8e16a5be0b290e62cdfdea010c0b6af57272a8de4d35789a84c70aa9c0ad6f1c0cded61c4267c5f94a63ee3b0273a5d96f48bae9e406b85fa6c085720d5cb7480524ebdd5ca9c63f0591a5f374b74a2aade441d58f3254c5db5a6c5ce85c69a2ed85d0945180a49d5ab0b46fa2e32bf68443b3bf4fa35e896959214c99a87dda55ac76f68afabdd8a6bc366083697983fd67a2425021f73b3ba0063d47c28c0a86874ff11968f2727287870d2be2d8c59f4cc9ddf778bd149427f5338074e946ee8e320d3ebc290f6c350a477d5c7c74a11b78accca089e16c70e7c246e7e547ba1138cd8ceaece93a2b1e8aab909d2350c74e3d83075d9220ad829169ca44bfbf2334c9ee7badf9e796deb3bfe96b982c195d9acbcfdf3c1b059ef1f0883e90c02a25b189d98b615e7a93c651af7a80e03a240bc392064bc4907a9df01e696a30ea1c38fe1b8fe3be5fe405f28c41beb2efd5b38bbf969d356fe95dc253702af9327d51d68514f197462a614f0fd4c970a88667ea2937958c678d7a69b99ef1002b1afbc934edb52a14ec2282db5f4fce6911ed23792462f30;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h10818f0be9755234cbfb6372532fd08d2e5a89b98d6eb6d7652fd3a2ff6d281d951f0f6b642e9b58ef6fa4eb7cbc8e6ace17a796f3f7a1d90fc83af7e2c306699d01681df1ef8710d13a70675cbd393218012f993eeed73582ed2f5482f467b362cc9104ba4fbc1db0cabab6c035997c20fc6660ccd0c550676fe71d42d4dab980e21178d97d0d3d890e460f1d695611753b0ab511b4cdb9feba19166549612a2c20c73649ad747f82742375d7f160e3d44727a4fe578d27c734fd7a308f218d3d7f07341875f23d8fd132fa8df156f9cb5c1d78cb8a113ad206ea23f9808b80b3221249f3b681efa57d5a986bca27bb081cb37c22c395bbd109d80077116a4f7e61cfd329851fe107aa2fda5f78736d281135223457284aa3fccc6395cf478666d7c6d9a015d7a1f22e54c835f871cbe07002018562f827c249f576276744c4be2dab5fb9a9a1887864b6bba13039b4b8f1db2135f755d5848cc57737e8f5592761fac6279d68d6ac9e98583c6ecc2d758f3a2b377d3e51c04dba255bf39d514c8ccd09997f747db9cc7cf8f5ce70b6450328783b6a99f28c1fc5993e1721fc09919ea0ed4190df0bd248705dc0782aa8a06c8420201bf7fa7a6ac2b7b407195750c6b5f2ac41cf226abb6c510d3db85ad14a058362e9de9850c7ce4ddf622dba483d2beeaace0f4ccb720251c0b36dbb3874e412216c14dc76cb906bd0dc801ed58093d967ef3d729cd8a9af4007d3cc8115589324744891f766ea699af8dda30d4c443e55403dfca98399fc37fc81d4586e778755deca9b5300254fd176e1a53907befcf1829996c4b820d3f2f76143f3f933d73b8a6b422d36c5eaa67b5ce2cb40eb142a20bab836efb7523c3641e42f78b7e791ed76da7bb894dbbf0316d66b9fdc1a7f98b126dcd5ac182ade533a7138fb5d457d980d5cd5b645dca84a4dd8cf1797b004b7395657e17538c30fb77d30d71e98786adb1b0c20de14137a759acfbe69232f2185d0c2ce2cf14ef7a5ec35dcb8e34f44d033f537652e736bf40a2566f7a231f35ab022b308c22cfbf3804865aaa13c029521c74bcbada79d7fd128a7511779b74f3ecc85c19f83f1aee1559bdcdebf572cd86bba6b90222294ca4f8053357cc8df124176099ad468462904ba47b5a4002b22dac1a0bff8f23015278cc6f5115d17e3abb4bcf063a4d211867851d9c3dcc43041447730b8f1bff5cc6f5748ad3bc5dc0386fa666db5916cd40cc51a9a0422cdbf24667996dd3fe06d3fdb6b0a436a7301ae790ef967aaa82ad34dfd2ac174d3dbbd23d4bf1a93e7908d871c4eaa77c1c5d2b513326501b62695e9b346843d20c984ad99d2c10354c05fd87ba2390ba0efd355df39bae658eea571a9d85ac7c4e1fdc710922704f1b777aaad4b51f2554bb20bcc7365984849a85c50c8caab1b4462196c83c392987d622b6eb8983934fa3b1547bf746d668ef1f63e40a8e6c6937398371f9efffe64653643f0fe6fac192556a8cf28ac63fe545775dd0868e9f38f5b79b1aae5d14da9ea1c24b467b6e0a120f36343786cebda8c91cf756ce333ec5f40230daf3b3397d250fbe00611182779911894fc4fb552cdc7fc9a8b0d33ac16c961afb9a6b1e3c42ee116c3d6ea0fad0e3051286c76f2f068bb1357ddd50dfcc6cf7ee06185f8aa6d4eb3667d0aab945c044222aefb935b99836dcdc5f6e5b9b982dfd132184db7ded0a68073bcba870300594d581d993b735dd3b80029cc07284dadb29156cefe04c8ede5552aa0544909c65e31884dd88df94813e2f6b290a813389a150bb2d29012745290591a9986585843825b7f6d3f22fd640f6b72a8db1ff7438a7424bb86187e6efb11533e65e557cc346f1fe23c4d71e71e6392eefbc61b7012a2c454a5c3dd780adbe506e35fee5fbe2ab0671fa02e14969d34a201ee76dc6ec5074e99cfa4315a9f8e9c5c5d55ef9fd038c1e09c6c6916ded5ee790b87c6b2bd085e7da40ebf8fc9f534a457bc83e32c9062df4fefa03d5eeda9126c95befefa7886b1d6a8f3a70574db7fd22d28f32ccca4e9e30a4164b59a346528f2ad7e80381dd697f77bdd631164548a128f65b93037ee2fa33a74bd717152142bcca342742cb3ea769f5b2a00c8e7fe60629178afb5585e1af3b20416354a062e7a0f760d55148312c4942e628329822ccee6a8b8bdae3e2fcd7e7bee26f5ad20906c8cce75096fd6f5e79534917256c4a07f8308815bae511d47ffd374b33cc7ec9f086f4a0d464e94b08acc9d0db199de7ef427e106820b68886c62cbaea974044494b76661a75ec6dca7dc5e9044fafcd4792e887d1a71ee75594cc534ab3465d3184533ad2ceb44686f1b89182c35884652417fa477ae3deb771c95bde5c7dfcb41f165a46aac40d1adde6c6057e08e4bba70c4649d071f50c414d10860b33698fd7186403ca494065802ec30ce3cd2149a3d72483ef0ba34932f16ccf0e0c22012b1d868afceddf583d943e80ed4687a621ac4043df1b1f3692c7b29de59c4846352a8572e8a78fd4e0cb0c0e20fd740d88d182e76bd85335aa30bc7e41120356580ec4b3e07a3dde7f8aee17b69a031d10698804d807d0f810b4df3b30da515d7021ed817454338d2809ba4834de543ad9d96e28344be8c1d00cc68946b9235aeea15ec1279f32b184f83c0f0a18d4fe1d970a25f5ef91f60f209ff7f3dd464158840809a41324abe1723a2f49a465f3e5e3b49f7d711dcb833706806cb2ccb070583c98568ec324bcbce27a1422f3ef55c41e9819451ffd0a08aadad81977fd55e844f9eb6c22251af309d694ae2f67dc5e53b8af6a0a8c7318e1a44c57357a7a2e2caaefb98f47897affee386dee3fb980d9bda42310c1c024ccf7ac3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc33dbe8f1f92d8bda60d9bc492faf24cfe9c1e6182444ee49e368cb9abcb6948c39cc516d46e0ea71f386d6e24952f0b8054f83b06e6fd89b30752744c0ff2e901a18f26790166299fdb501c69163cdc02b095d706a6f31ece6a9190fbc131b407307fe08fe03545f6105f17e71c56f7ccdfa0abfe2e15bfc1d92b502423bd141fa8a714acad2f12192aa191a5f7b32bd6093e878ab02917a52efdd09f68a4c031cd0b05f11c579482f43a3b58e7f6fc0a5facccdccc76f89a267f245cf40e3cd5efcbfdd96f6dad6fd7c107870ac92fdccc370834c0321ca159fbc6071fa849bf1474a1c2fdfdab97c6076490c57b3c5027db7902bb07caf02afefd57fa10939a2facd22702e3669efe92f867320981127c037d5aac85d744a65ab96a1795329a69d900224caa3a7fcf9d7e9c204d553c00db5acb280127c2e854d960cbabef04574d131bff54220292933a1581bfcff12441484c61492d90d9d2c27114b5eb9476aa9d3b79aec77941d7f96713dcfebfd28589ef9224cffac19f5bbbf9d7185d35000ed0b1b1fb76d25399fc76200f410c6c89d1fdd6c33b71649d19707fa9b2eb5a8f88edf749238eb693a97f5b027f1401ec20168f35ffe2e31f333533baa76f138719ed3e28ae06f41d63216ae24a2cae02f8be46049d763851fabc890d751551c9d22f5cb9e20334195c11e0f5b07580dcf50bfecf03c5720f58836191e0ce5bb39a19d2e70c71cfb7dbac043b934faf549b44d825b2b878ba0df12b8a1b0ffdbb34b552fa3babf47a27e755dc6d463adb044883a8c9c843bfcf80c89a46abaa2047155e166f3f097ea7a374b3e66277995cd4ca731957fe9f4f7e1d5692eb11d1fecf9166d4aefb275080c3fdc1e236835d672af5287a7368d81ed35c5cadaf0bcc5e0260318546c05bb10204a2201b7d6dc15f8f252b0fd1480de3f503ac1c5389e77ede08791db37f84182a71b0008bd300002e65510d37148620470f48e679a5978ffc81fd77ee98616179e2b18401b0f4f67f0467fccecb5069c5eb0077092bff0c211e977e24cd5ed793e14ef82ab31c353007fa26723d337309beafc5d3b0c3196a843567088a758722b1895318e3001353869abfb263c44d0beda9012dece7349a859d7e0004ea0a96ed1db2b32a399e45a83d0019edca74efe671100463455b9414f01b2265320cd656404b2eb1edb1b81d1bae96968ba1d1635ff180fe38de4fdda9df0f994d12419f279a0e60b60dc714d5cf5e0792564f9a1428962d9db7f0f168ae9f0f0a67e51077f33e2185abd6a7284dc34f7c166267336acde06031344f817559bcf8dea2eac238681da7fd1c39511be8f232cd73553bdfb0c256befc4b38626af401cd487e4bcc88d9471ee16916896ead87dd9db2c33d8f292e277d71633b1ce6a1364630f9671e2cefda2b718369cd955ab11a5a2b69317e6884057071e706683ae0816540caa398802a83b6842065bd6d2ed6ea43c0ec740c6cbf71e1dcb99292a17529fa1c174f88544196d16ee04c17644a193cb22a740b5c38d5e737f82a30338f44148c4f93013a91ddd6190f765b8229e2735fdc28387b6d7c8f1389d83dcb12e7b3106fc497908982dece9e80b47bcee50d61479e9e2bd4f89d75ac605936bcd86dd3029120192a88ac05db6dd801c90b33b6dc543b590da9649d19f90398ce32d64645f4de7fc1652751d9629a267a8bab16a231115325da74f3dca83862809744e0370d267fbe19e476af95d6b218adec184c307cb87387d1d46a1d3b998859c29b8a525d11ae128a54dae02050e53ea67a05fdd1580768226058a593a32a8a7b5a67e96574b95c3ca06d5a56ac79a73c1c76fffb648886dcdb1787e37fe9e0df07d283300bf544d1245da249e6ca032b322570318d0008cded2ca7db58e8eb3c60b45b103cb2c032d82a0cdb7ea63d884ddbb9a1d8518faab05ea07b52dfd91b890a46c20f5aea9483a20aef4aebca1016d9ed3db3846cf8eafb0dc0e7dfd911a27f9993aa0a6568c859aef9ba6472006552a5f07a31a719ef28844b6625a57d7fb9eaab2bdf2a4a4f83b925dd903ac3d1418515de9c27783d825a853379efbf52f00b584d85a7e41d43a98d03d9f053c0494f7cc9c10aaa5b701fc58232f0a59fbc62284a826f5a6b3c52d2f7e1f3794cb36f650c40adbb3f1f97c6244be95850d2acc71bf72ee13c89d8dffd2de7e060315692ecd6d96305c68cfd4ba4d9fdb0bf117aa39fbb9b1397394d03ecc9636c873b5b3a9c49bf883c9a08e71767fe2828eaf44269524ccbf5220b309bfa22788a876bfa39405468c05aa2879c137d4be6352a07722eef80225deac6d0082f7e162a11189461bfee2faf404662cd86096ae5364908c9ab48748af46f5ddf25c8d6ea55b226ddbcaad23207916936381ddef618121dcfd11aeeca0dba84b5bdd78746b871517ceecfd316e790cd85553d19f1add92ee4d9de8ddf672238a2a0a63724b215ba1cea73103a43b7f6346af33240122ecb986b0c8720f129cd90582052580623aa287ecf8237141bbc657b125b9ef3da1990c2432480a3ec382f2b12d6eb2835acb5ee793be9c62138c3b23272d194fb9b7451d7405df3284813d3d32055de75adcde5918c9ca37ed76a7e28ba7bfa0108cea48b2038712b8dbdb5fa9ef26d3184c8ebee239f2a604d731b06d8ad52e27a5bc8a39e0a1a656192943b4c6146c28480185d526546b1823ca58bcaa8aa280aa109ba0c545ad4df19db2296383cd6ff4c89c2ca9768ff50aaedb7b1262d24e4333f2d33f1370c069eca6734844e2fcb4d3dd9ef3213981c14211c8c630b8f84b758bf770c0de02a785b3dfd3288da510505c75c56725ac40fd870d2f4b670ad920b909c76640435;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3ce9c37c2d79ac93200007609eaa0bede32304aac619d66e092859adf3b31d29b4f33fa98a3462ab22df0e4c26e74b0fba7ddcce9789bdbeccdb8760bc02e8e1a49b0a2c922c2a7c9a804750f475aa3aae5476f4bf6d70fa6cb7921debba9d10cfd49d7bbb39859f74ba25b3923da7534e26838fc7d22c9785c9ddfe0cb4212a4ed34a4cccb58d534a3d92152ae29111ddfdc92258fa0703d9fc3fac63e787562013a9edf4ace2a341af532f2bcc81523e4547f2db56279134ad1e3d67a0c2be3be8ebf1ca0a66833cdf5c8bebfaa91af447fa10dc764d706492a2ff318f9c91f7fb223dfaebf14f11f55056f0dbe685a92fe56d1df404e77217c39200b46dfa5a4695f9999d3f8946b998c2e55e83c846f9cce03a5d89f42cca970f3b9588eb886dc031792bd55424de4eaa888c0517c0e3bdcd1c0cb2074a28683a06568bd2fbee3382621fdecfddee8b5a391b56cbb9e1b3e5216d4d5834d6dfc86e5b9605f13f41a16f19804a3335a2c69a29554d29dd5e7958d5d87c4a1bd4e987813534885f41d1c783d78136b0e9c030c744831a43316748a1d9fe27b33946c3639764a479e3f61a32934ddbe9feea1c64ae2b6aed57d1023001b0ca0e99f5824a41fedfb4526859555417e34a50a0b2bb4883ba35d9602a7e45535866ed04b62d6227d6f87ead66deaefed592942d10a7326008734dd9ce986b058891d59f7f6446ab9f3a57818302571c9474562370c179c55dfbd6fe5030f7e872ed0d63d70c3ab1d73ac4393475654ca7131d45014d9fc119026e61efe380ee451b3c4a308f8a1eb12dfdc274cedb4bbe05e0d208175f3bffe22ffc26fdb17ffe52ff339232ff5918f33e8d4b1ae25f690e9b1755950cb4b88b61eb90a2441ab3cf7d399f3c31d70484f51277b0a5d3da4ac2598619566c80453b09faff68d71e31f12058d0af090a2bf9be0e384e71d9a44c5ba8c6208e2ca9db6cfbdfa52a331bcf3bb33e9aa9a4de765482eec6f236ea0b9586eaa46cf1580cff46e45c7add917e2431f7c9a7456d2138f032eecd12af2e8af4e134d29f7436d55eee7b0ce09e6e4d470a0d921ff6abafe4d837700e2e7e4499c4b8b7b81666f799ff41a67b1987a7080962348afea4f5a2648365b8d7cb56f607b88c521613bf20bf530684e888ffd901f29b0063748b0b1fc743140dae332fbb2999e2aebd22d2ceeabb5f758a29a35fc4296ce99b71079e7fa458a6dc1a003287587cbcff12799aff1fd42f5983ea1a8ff8874bee6507a4d3071047691e1ecbbc47d2bc7119e038bf403e955e4291af12c72ed95dcbcba3e242142e301b0dc35f6332adaa95197687e0efb91488a3458dc55f9d280314eb774ce5165e22b71c8a3290d1dd5b1547356115ce856d3e3ebc7bfb1899c687d32cc78e80136d009581a18221f76bb61c61ef1a8faa1d187d4f516e3554f55f9a9b2f49c45dab6599fc71e39c72ed51b229b399819ba9bfc654b4f7e5f6a9d5d8eeac27fea97341e5a83c10b1dca0ff029ef1502c5d807936e561da03196ae72fe0295a3fef460a0a86b26c769c38e2346a68b808d89d5028ab52160118d003afff8aa085d225b48ab56c813fbf884515673260db6516cf383a7e1a56562aed3326a146d28addb4be1cb6701f4edac2d25684a91147d70face474986d7a883b0690a36d95e0ca3a8147a1071a565983f3c48cd18ea5b85b85b2dded22cd2eb42b0bc6d920387dd3aa4b55af0d62e92f988bb2aa2969635065de8f328503f462d3fc3d1e2a0e594b4af07f209fc5d6c0b232c48eb09f7a15508729848c56f5c68a4e37cfd5fd84ee911da045d995991121c5a168648249007c3d67b55b5d84206bef2673d725681b6a6cda251cb736b036b03f8568a8c8d51ab55e6b4d502f09c1f36c747edb4f20236531fb641f8ea81e61bc04a56bc6b01f56818fa5a2bf39bd66235ba2c55f20f3842219d22bea6214b545d29c4f786687e9782fe14e95f644ff46671880cea4a7beb85dc64592b02e87ca34c7c2f988d927ad7d001480d4a35cb48d8e4100bdde2a9c1aac7dcd0dafd2b5058210a02ba5752322c04dd1307ddc833bdbf10a64553b0a5d5d5f408571c85b15645068ebac93e2e0a42927483932d9f38f3ceebb8261b30d12e712da9057ce3921970e26fc631f67676f43bcaa4d949c885a2b64fb1da75de5b0682f7a492e0fc0980791896b3344bd3b0669ce27b318460444310efcca51d2db94f692717f7405828603147e56a8e62a2a87bfe35a5573cfa5d284e1df505152252ae874de437baff154fb15db44253656198bd9ee62ba4e0c4c9899f402b9d2f0db92c2cdc936bd66c271ff7d45215a711bc49caa26880909afc307eac32214e08e7bd4753c4e4625b80474134b8870fc8ffaa1ec72fa8a7a53699f7b10369d07577484e5028f13d1ecbba35bf3f999343e404961c63b1b8910ba448143a32d13d9601bf7f51fd049b9b65785327bd3780afe3f77f3509a13a59faa1d55b1da107714816ad21843e95b4776f5057abe2642ebba80079ccd45103b294d1eb6266fc233dd3481fa120d012202f8a69f86afd64d758907ffeaa1eba4c44e48f7cd160dde1b7b74a0432e7b724971d8f11aa1dd0843cbf2417b3840ac128c590ad41cf99cab276457bf0cec2b3e8eb661b37640a5a3a34283a9aaedc494307bfbafa016ee7d1ffd64e63be27be0c312fc868c53582a9b7b227735df9c3e57671c38a2af3bd7ac789a85d4d9b2a601b05b226c539978606dbbe60bae63d615ba680d1d65e7a7d2252cd9813b0a8e236737ff94d77be8dfdd3ae566be4e008c68e3c7306082609fa703b7358ca0c73cc92b0cf2e9180dd205b217d77f6df553ce366de16d4f9df352a27996c4735294;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h199ff099e53546f111bb81945fec910febe0cb14a324250e5bb548ef715b7df7bf79d6da1ded650ead05a0536f746f5293c2bce242bf6f4b8b862dfce929fedd7606d7322ca90b6e10c8698be72b0eb72ed53450f8bf64c200cd498037c7acb5545d9409b5630f7b5b4381eedfc1479c4ecdd08001861392f37f1fecb37477161a404e85d76cac477786b1da305cb197e5e7d0775074cd33c96b875c285b12776500fabf2506e81ea6ce26a7b56949f6f1bc94434c8ca688b0c3cc1b5ff08349ac3cf1be5da6360744aad792867630f7cc481001de3646a9035c154be7d0c1d22735b722464a34d5b3ca53b2c6e19931ee4a9f6b835a7c63a7ec12dff6e4bdbcb44b9a5ea371c0b4e6bead6d9b00f86912f7487eeca669a737bfc67f1badb1bd968a12d1a7cedd50f2fe2a464c3bb58b991712ff77747a44a9729f06894a8d74fff9ffcebc0761c5bb80593a48e2b0016d307c0fb46cd737f0135be1f06baa76b8ea17696a7421e8a10a0139d10749429037c1d7879302c8dcc712ff248c90cf000efeedd6ee7e068c19fefed122d45e68c0d67e15d35dcc516ad98b0af166e1fa36f2d7cf24a983b2879a2f049d843a22e187beb2b9fe86e9b34dc4b3aa31e2c250052073feeeca2e3ad706c6cb1ee728035d272b36fba5aac59201b028b3c63e228ce5f8ee261cddc36f037fc6db19eb6270b8689d3701c0f2e3e3b20fba04f1e19a6572da099c57577dba492af53dd7107b40a0ca9659e02b798b82afcfb11c044ecfaf09e98d69bd7101c3c15aff1d3d083a84eadda1555ef2ccdf602ce170dd59c4b00ab72f4338db7052e7568174f2336c4698ccd659dd31430d9f52b2fe273deecc9aeb103bef1401eba0104025d449c7deaf6640bf91f220ec41f75389da03656129a82bc0f7dff2afefdbe62c0103faaad9abcd858bd5886ae5d4bde147ec61ab9e58e904f06fbcecd63a3f5a8496f8e06a76d06fe1e57b8ebc8d44a4aa921f7bab96c37f8c9d3377ec03ee313aef900ad320423f3e487b7d18778f8b2b7b91da0d52a02392e64faccf4313235d7bc2f5fbf898f91252ed1e79a0531417b9a2ff8075528d618decce26a25dcd49926dd020d3449b4c04d1c600da2932dbad4b7fbbf43732ae4df550444c04f850d1c2f3a993b55bfee02365203a7f12ec6f264312d70870d75befa48266f996563fffd9e6b97b90e45d9b9b4401e8618a2b0aa0988f30eae359c3c6e69a3689ba757b72ec781c4296b4e882d015f56f29b3281fd7b0671f74f76720e823b6ff1efc84d758c3ae8481c33cd993ef3119674581e6bec51be150da5a407a249de3d89455d9a82978a8ab7541a6244436f2eb3d733204f53ef78008afdd124aeab9455e2c3403bc177990b2be702d82b80e7d6381d8b8ff5d03497c2dc71f4c354a3cbedc900b96077d6a3a17c3e469ca19e96b896074277e7d6adc9a2cd141eeb3018e4b0b08067dbe103871c0834a475937f935de845eec45a83022366752bc7b1f127b6519864adf702f7ce89687a3e0f7807738a3cceecb7d9af38933209854343b6f27134cecb3d14c41ca2aae7504c566297670c18caea0b5f35bb3af1c2e82ca70f1ff26ecd11d32b8265949bf92de709d69c9d8f56484018a02530b66fd07959a64840fdb58df8bfa5c537100c30e5526feac316644a5d05e7fc7096bc1f952b0c31886cebeb2f009d8d2bfdedde179ddea5f1200fccaab8fd56ec6deea93bb01629d2dd465c5adebb54bf07f4c4a429424f6762176b7b9246a549736f425bbe780028f975bbd965befbc544422b65d0e15006f93c7596deee579c2123532b05c2a43bca849bba4f3b677ad023e4c2e9996b5eaf8e22433d0850c8baa37d389089f83618b9390ae18de5cf1485805d283b35fd3688254e428e3ed9b0b6716eccf1e40710377cfb718337459f4c1dc41a59e61053aaf5da63c4c196158941f5a3f03a2cee5a548f8268af93656912d56ed57c918b224a64779d9e98b1d66c24e598ea2ad35bd1db9c2a8cdfb8d4841a2c1b2bf3d10e917940eb891f72cbb1c1d3b7a11666acb6967c509540406cf2ebbdb781e4aad67ebe9be264db7bf57677bd3f7a3d8a3193fc71a51e9bc0eb2aeb3d945d6c68d2b3ec57cbe7a76148b6d6346ae2380da459df7ebfcb20ed8d6f95c7e31c21cf205e324aa7c298f559e9e76191b0c0679f2ba58c2da1b47916978d53d4401cf3816cefb85b61e87389f338b279c69467b1bab80102a62a38a0853c430692aafa305ecfc22fb5d7372eb01da315ecd65b547490d38d076377eaa2054f2098cf9f96e7a9906ca4a4c89718e4e4fb9da6a54c731db14425302df1db1064ad96a34fc61a384d4c614910f5e6f82376f09d7c5fd15d9bea0c6a3546b9d5afd83073b9f9de199fb8aff7af63b59f08dc5f382c8022a7fd2343c67b9b5022f409fb8bec32056c71fc0e3304e948f9e91ab63f62052eff4a1030d149862af05ab05d67629fcc4a0bc4d9e782715a8e0c022a2e73ac7f9f1a61df689e670cb4d95d426f23c62baba3ff6546077b0f6dfa3cf6a8e5737aa4ea132026da2ffcf1357ca6eb5ecd4fd503e62d92290b2524ce3c9ef455e752059a42cd4838d5b36ca50f422c465e33c73900245bc3e05d314e74f71fd6543f2ccb0d0749dad13dc3a68741455276427575397030773c327eafe04fb082187e18dc463ac6800589b2b5fb8f0ba0b5161054d1b07c69b12c4f4b7420a89b2a2e2af2c64f4ec01a37f98afaa6669ee91cf1e1ef089958240684d93d7bb5da1861efb097ad666068716eda00b047dca3286d912a993da444d68198520223fe92214c3c7e672493aee552df8261fdefa8333a14b286a7d3987b22e14c1e41376f5713f053d3cfaf5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1c21cd022bb6aa8202abb9502472137c2ba06ce969931ab6e70f3e5d2f3af05284b904e9261c16d37b57ad78b28a1e668be16bc296b1abc7e0bfcc0047ec65e17b75996ffada9454ba2e9571afc70dbc62f48d85e2e04b00d24743053a7f8215f6f4032f3b48d280e09caab9d864a479e684f57f6b39d51e970b2593183493a9818fa855af7f5d219d23f3ab82a6193bdea72a2460dd82945e654609d605c4bf26ff06834e43d3ce23e35372f412f5191ecb6bdba3c9cc0e7dafc53d9b470754f022c4822c0ae81ff14111ebca1af7088507bc1bce4f186c4ab120589dda57d00f23be1c17909a27c3cbe0e5656a95e57df3d1742a974f91c8b3ff27538c3fb1d9f87e511d9666dce273a4caa77784dc6219cda8b0c22356c96f21de54fa30c08b7b25a9742ed0b42c06dea5f0436c5432920006b9a55fd3959b35438a4e215354a9706454d9e868eee098bf5f3a89a07b624faa0ebf137ef35a9b2b23dd1aa3e9f8b6e05ac3820e507692471eee5f8314bd18257db477d4e08df4ccceef86a40646d560959c3c161d859dbd33b671631a58ee3a72b2904029ab359cd950938c0d946686c3af101d42e0cc7434a0b879c426a5b3b2d1d9dd1f80e7d7c96dbb28bf310d5d8afb45c5944342f6801b91ee37dc7365058e2214e2e15dbfc58049a5b086fe267940f820ef574b59a8791e8a7e6f7eccf99d7d42614ce79fa7d815e1efcf69c3a50c61f0dca62e5f046387caa52aee059d69cd0bbfc1f640033396c42253e6ed221b0bf102d213d53cef5387b94ca92f240ad419d0e55abd7acd107b82f59fbe9ca3a49b8fc1ee96f03c620dc22389fc176ffaf5319bcd0b34623afb0af1c37cf9ecdbd9b780dd4d377d8f076af5548335c5ff85b785a101c6a5c88665c466cfb606a85f1b270dd0d15c51c2c7bfbee1a8eaf2a2fc3525ed48421693d11a3ab97a7f668e475a1b73cd07e26bbc0d5c3e36a049abde13b5507be5bad0adc9d90f045a86fab0964de392421c7ae2ead05c11c5faf6c88b55f5ae4344047c298f82bfe8cecc7da1f85f35a57e62986b2c04ab69340858bcde59575da63572372f1f074ad9684550a3e4bd3953ad86409ad517465017476526297e78c9cbba2fe08275f0be03dcae3614d2d8c47e456fcf22b86e5d73d3553838e4bc5880f2a58f902bd7990a79cafe980da926e6def4d5e3e86a78065ed5a6259e67a0b924a74fd369d8c27d80cda2ef514d66b2c3b0ac8ca95743b967750ae4aa135012ec2ce5c16af92613c87dbee6bae1c49183e5bf9ffc35d93d4310b445b2e51fa9e26d9056e0adc7ae6f448209ae6fab38c26d0e49c564a03ccece3ac1037f1ea613b2d13922bd149d720992c7740ff54e7c7e6bf8d02bd0f8fba71500320df2821cb20f58991c95e45bf083d391889ad0be2faf49099ae77be3c14e497c1de98d79b7132bc38da077c63f3c863929f65997c8300dc2914bc7a7444056cc413e857776c4f31e9c6cef1bdbc510bc1682335d3b5137e7152785150c6762fc379447f3596361ec0ddc2efdfd958b00f0fec8eccf7eda59b0208191a0d44df03b36d3b427515d4c91b8aabc1e9b8e8c7ece6638a3fe6161af3d5f47961214be66a6b8d6459119a7b96bbb003cd81dce994cd75be58797febd00553075f82fbcc2d570294343635fddc052f3f01b1aabda06ec6afc5733b390c7e96a09855be7214a20de3c3c8b6be58db838551347dfde99a5716eabc55b9eb4211682259b4c513a226f4df2fe602e0b2f8ddcfaf800a4beb39db6e8e3ef4e5b2fdd5e072d50fe4d510635e8c8ca07cfc65302ae2052d0fdb6e04bcac0a62fdac2d5bef6ba3d974a640f39cd7560b4f33cfb92edf6020d5641496ab2f9e2a6fdcc63f1efae418bf5e9276a990a2a35bbc7ff59ae060dfbb1bf6c491fe997318cfce6440f6e9b8f5263a172e4c5ead4e37af252e9b32e496118b9f33d09363e659f0a22ddd8efefc290bbb191681bebd2115aa5d9d87040b04fbab9dbd7f1ac558cd0da568350488e5fb62840952e46fc8bbb70e7dbeac71a3e5a35f6dd90c9b653c2a9cc4a8c273726cb77e554f5a9935fe59ecef029cd024d5299a513e12905cde494b91515edde28f5ac2cfd29edd469555a15e7ba299847a19dca96588443bf87ec6f5e9bbea25cd629d50e869e982a419ba9140ed06c7aeab07ab6e66c2f104065b47ce4c6da5dc71547cf092dbb49868c24fd58e6799b18cc86899dd95ed492c01bcc816e5e31848f1656c9702a5cf9152547dd70645f0456c12939d80fc5ed86326be30b0335f0494905282bec85d2e6f4d03533b224ff8a59b31e27160777b3d4c1db48983e457b6dd667675092a2ff78e07e785eb2f2f73c4c5fce0264762201223d90fe84ae2b8f69e610bc014966a244f554f8035917ad79e8c6f24df1625e0e7f091f12eefb1f1c3f5e5baa9ab5360013f6b571f9937c2a22934ef91cc4635489fb8290e76501ee52c7247ca96de84195cf36bf725977b9d6abdce3d4cdb271beff5cace18a04b5ef66c293fd7cda6ba771345c4f8de137ea69059827753a580a93597083ba2b658221d3017dd7739017859118b4f7e726ab3b4349df23e01e1a941ec64371a4b25cfa19e1ff25d2895e20c92b3df9aae2af3b270436428c4c5b2875b26a575ccb7440af7f515f4836d87ed744934a40680fff21889fe51f749f4231732b19dfab459b34674e84011918e5a04918dd4aaa7ed46385bb337c3373f787e9167d182cb15e184a8640b26bc3ee620bff5979345197ca6ba2f186ed29408caefc089e2ab8a9edaabc5adb874539393eda90f144f8f89cbf71d2fe5cc57b3477cb5402b430f7ab711dd531bb6898428139488252b24c2c8b2478faaed79ea6a5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb0ec4116900196270a5555c781d2f498ac6c1d224a0fc45c0f866dbdd9d533630181a359b96b10abb18d319fc4d5464fc5b93b9d474fa797a7b7e40d5e21880ab25fd8b1388016a5be4e21146063177f11b469026579a0bce757dc6ee67c46b746dacc6f3fe29783efd1a3915adb7e8ff93456a9e8616aaa82c47c223211601c8dc738c25b1c3dea6044121ed5fb2b8de5bc6abc41a2331d5beaf3bef985d8152d460a67d765f823ca092ff29724f05a289a44a38f7f80f6d0d4467df1bf8a75a272f4fc817916522c15262a283903bf0531d3966f036b283071d3a3b76dce6eab65109ce7e796a8a59329a81958f43f766fc8abe1758560dbbe487f881124dae9368126d5c2caaf32d6d5f051a9448713cbbfce7775fbbce2543633afa33844dcc6340e24db727615afd8bc3c9a995de9571791f1de6d62c4c89c9b7c42cf411674348682872ec312965e187c35ad8260e05380aa7c8cdc26b410eab4c7e635613f7f7535a51fcbe3d0702455c037df2e2a8b5cb87fe386a1109f78144324a2e2de99a50d1d3c54b21bc63e95126b633b588539cada36030c6df1938f69d25f3dafb3d9d458193cf8120305931649e3e85b1747cb0f1e732a0bf723c9fa82ea4aa153995a2c003c2fad99bcb3cf8de17b123a1ecb53b9423ce4b13b57c22a877291738023cfdf0a020d3adae78c325327d062d0e8c029464ccbdf9c526bd7c58d6a84ddfe49ec474a192af6c8f4f06711f282b6eb36dee357e1f92dcc47f1e30d83e3da662600ea0e53e90170c63c60503cb389465487a016a58f3e30b8add4d3c271edc94b221b577cc8078f3a294120e6429cf1392315a6fbb83c69d1e21ab3377665284739f602cb560d2dd8ea520e6dd8a87791b25d11bd79d2da5667df111ee20e1b76e96193854bcb444a41023ee53e99b91e180add28e00777480a5e2793e53a11d9c70107baad40a5877bdb3fe8664127a72933c6161ff0fb11ca663477484bc0aa0e4ba081ffa731b994c7e03ee06fea5e144e0c1301317f7c04ff24bcd71c2fc3edf2a9dd43ffa908a93264dabde5785df3df0c8d36a7a6ca374c7ee2d8c55b75302642af67160f3e4c545836783a9fdbdd99192774c7c8cf371a4e423d7f22cdeeb8a005695ba36a3065dc0d3a785a39f6336b779831c3c495986204eb09cdcbe71476757c4327d4f60c7678ffe5e734af9357b74a360326f35d94c54ab61d3df11997faf53061d412c0ec0b745dab040a60573ae17bc8a39b10be6288b1be400415889e43e77bbd2297297ce8cf3958eccfaf3c6645a8afa3118ebf161c6443c87da2bd79b6a1499b57cb189e5e948a42c303389c1dd2cdbe8afa1bdd36eb0496407614174cbe7ebfa11ecb5e6736b820b283d725d94fdb7d8a23668e8e255020dc89a3602e96db610f3761510d857643bdb4d073cd8ca2ddb163c73fb669a61fa626e4dcdaf8a65721c64f9c762764d605e9c72c0440872c651b680e1b2f3b4bb89bedb0322bc50ce4d4d213cfbbaafecaaca43eb57d9d66368c9f6641b3a6ea10bbabe92dd03ee4110b3ebcc73e950d50812f990f227d33cc652b1e1b2c3d5fac59904e78adc47200a100a9251bf0241d4ee24729a5ef3c4134eb99ba9b226e30af9318777a982668a8be6893c458b20d420a111b6bddf1c849ddd05b423f9404df20b5d2796f5bb5a7a82d854bc71e7332d41d91a05a75e6fac492fea618b027ecba2211eb1dd8b4f7ba8fe65f6f46a0165830196830fd14492b2b2554b0f82537b401d935fa8e7236742f5e979c6b8b1b52d437cf51d9584530e7236122c45405d18fd5568bdf7b621abd1289b5b2836ad790bb46a608b7382b475020e8c929f8038d6932041477246d68bc1575f692fb19c5f4ed712357f2b1f677daba332d7e29b84712e0f0fca0c8c2e0ab9a6d5f289186445656cdd8502166e725422ba0888a6585ed12bf198f3714bf6e84035861c9eb55e1f9476876ffa791498e70d16786877772cbb7c5a276adbda4f5b296a14572a98034d557f759b482514b2f96047774a9c4644136fabbc6306111295fd3a66489bd248b7bc4cba88bca1f44da462e040b932596bea6882edfc014279d453e431134ee5642ed67478d2764a570880f34cef5142d68db6332cbca6f29d8d51cc07b765b5a9189fbd5478c90b81770c117cd3c40fdcf8bcf33ff61c07c9bd312bca20b9c07493d6487f9aaab5351ce065e85fc7364df5f527498fd34021355d3238a4639bb4482e5bdbcebc98131ccbff5b4920ed86b2beeb940143b7167198ea66b2fac111c681ff450dee2fe6fddae4cafa4a90c914d70720bd6c876f2d5d0424538c0058745ba9d18bfa28061fffdaae3d70b13f5aa10dca55733214e774d2a9907107e52146cd24de3450a8033f2cbdaad10239782e50b367c9fb91bfc0f60ad5644863c2b7754715c8b7e213b5270c9423bf4a4c127b94284923cf4fd8133274d37912270f20b54ce1adfa3c663d09883cf1f4871246cf046fb1b06fa58e06c77695f4636b821eca085bbd78f657d3c877e5d1ef55df687959f3e8ebcd261d456b9708afe9ebbbcde9cb64f7728599cdf82d819b57a01708af94a96720e534feada485aa939b65b36624e523b251bdae1025b529e721c1e3392f1757184c864c85fbd50bc51ce6b4cacb2b8dbb3cb2322771260b1c620bd37bcb9987828f931c89cef209b8d59190e09c1be863eaf56648c52ab7b1925fffdf112ed44302fe696e75a3d8d01a196dac851183771687ab3a628d34264ea53f2ec7976c7b6285de3a6cdd488ca4079e32a6df1f44b8b83505a422e4a3479f15378a88abdd47972a02bd8ed36ce493bd542edcfe64b206060d3cae314b28bb8b023f215357d1fa7aa08d60a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h127a3cf40b72539836b6126a3acc750a619820a35c77c7897518b643b46b33b2a0b780386d4bbe3528bc719d54be1c14de4db866dd03b06779cfc4fadf32cbe0df5c5a3c6a190198614e92f7883de24a778f7cd0066bcc4133ef39483dd0a240b425769ec93af4ad93945984b8e070b8e1c7d015846675a30b8bbd85209f293c0f81ca333b82c5677bb394bef1505beb7c4c769a1a4e9c61909bdc8790f6d4b0de9da44146d352cd7181f5e021420df27b19d2028c3f1d9946675864800d90c6141a36e503e1ae9ad3b3c18025ff274867db74945bc22e6fd6b0c86da97c72ee14956ef7d92e6c4cde78f35e26c24d096e45480789f98347d5167c511e023a96fd3d4ecba65aa7df5c29760ae1e27c656878d9d1c3a36c4d21c91b83d5d8fe422fe2f5846077dc8f31290e0c532c834ed238896f440255e7115ad0ca73aaacdabd5d7af37116448f2f67019d662c18bf79f61f10025630d840e8389355798766f0328c5853ac5df6e4aa9ee5bed033c585a0207628fac7f9a11719147932e39e6b0f1581e389385520fdd853feacbc22a5cd5b0e996eaf74bd899ab22c039dd7c963e0477343c2d22faf98ef893f2498c81921f80725a24888627d882d1212665d8b71a2dd98133ec0e9c67b61513232f56d075ed880aba0c3af6c58886ce4eaf84028d535591939476a3fe834c8383801695a14c8ef055a8af7006a2a9d3161f1e9049e64ca1081cce01d0c958d0d1d76a44945b19eff6de80336fb1bde208b6331430f142f78f2ec900da0b9be5cd6beb323df093fe9b3ae972d43d953b7e17a1b67e7b2e21ddfe59955c57897dbe49e61f5c36eecd553992b80dc584a78c143053077589e20234bca29fd63719cd98fa4b4782181244ab1e17a3cf398d6fc6ce4361fce930385a7d9d115467a6fe75dc7c2529f537d99b3702a0467fbaad12fd2162093b0c05dfb4785064609906890d2048abb5c8c4deee72854f56c26774340a76d16b1261cf760e0c9bd18f6e996f82daee10aea7bbfa1db6a359e861307885385bf9bc59d61d83b4e0093e0b3f55d584a74123107db91186e819e84c9efeb09324c1c4505d89b14546211e37b8ed01abeac2a3e5794e2d0e4cd9232f8e86e361c95211b3b2a7920517b5096e83536a0837790ffbb6cbc2d2bbefd17cd7c5749135f7d68ad62beac7142a622ae0d2c2c533fdc9da8bb8e8c5a647ab72884227ce4c7f383c0a2da384812d8af657a29a339b0f5fba5f496122fc2210084d1ab3bdfedeedf7d8c68a20416725e2f611a34481d7d010982bf5d8dc3ac218cc2eba16e25fa51dfc88a598820a7ffbdcbea20af14705575475a7a18585d308e18f3e8c3053ca754eb8047bed76542aceec1b4c137ad40057793b4426d122f0692fa498136ce4be552bac20d48c2aa8d76d506afe60e4d76a329023b797906302b917a36e65b61fbd0887363ac0bf713ea15083671d7d1e9486dcdc0d26392b431a747559253f02706340a6ded3000ebf6409b5e29b066b8ae1f3b5fd11e8b55c87de0521fa81a07795ce0478b6437edbe852caf330b6f83eb5cdb77abdc6dc945e4d0a78a5dda8fcff59463b9bf8a1247b3212d8f7e24f08443f9d231432011e349c97f349c3c2ea5b265de9ea17c56690d9392135047b6c22553e41a696f5673ea510235fbbff66551d14c93e9a395adc3aa72b3196d5936aabce7036bbcb63ea256f79d6c60274611f2193cb57402d41b8a7a7db30bd6f56566997014ebf61aa880a3f4340f7f26e08a3e08dfffed435bb31fc1689922e5def6c3eff6cecebda8e3326047d33d5f3b1702942dd23fb05b065505601db9ec279e7aec9a8c34f99294f705d1f95997fced87f5d9c10d25ca1ef35db6726ad4dcdd4b1e2d4d92f3e8976142a89d55e3b039de3a8b1f78abf043712060c58d53526a30ac1d84ab5ec7dd44ce1d3a7c734b7a6688b472ad787f5724fdd9c75d6f40bf2c58ac55e0247a86bdf36d6c404460416e55a4a26d60052da761f67ed8029aab916a1b8e0784d362e85cd1e265161aa53daacc6faf7155cb92a2de68d879b3cd58a6bb957e6b718a756818a7ca4c409bd5ba4d64ce02ba9f8ce5a3b7a8f0adaacda073e83615b26a499a8f0f870860a36cec7badd204c16d5fc9541d7aaa39133034c594cda37ea2bf20f3848cfcf5b537b414baa48253d85d5c4714c1d33d358a6ecb7cb2e5b90eac81d2ace165943670b57168638e47fb001bd99f80936f07a0d29ae85f39272962aac9d5e4c423f65d0e1a4f7a8e151361e98d0d32fc2ffed8b9ddfb6ec835cdd353cc396662ceb68a132112231b8da18e7f900183b7440fc35da137f8f04ccb67fb83fed4da18e1a0391fa8549f00f673ce1da35b7888340498527e41b05f21fae29f947fcee1e659f4bcbf661e0d0e7c6837d5b5e922a4b0547c6682e4530e840c71e1f092bff7a2d3b9c6109e4959efebd819965c179b4588c6c239a6909f9e4c89531842669a1160aa8141bbf00086b88e1bb922c8a728190fcf4db388ca81e54e3a03c4557c77abc641143793906e85f98484cdc72ac3ed0795e96caba3177d02f6c235dd738ce31ea26a3feddf7565e3d265b2b2f6406b5e629113d3f6baa30584360eaee04782765e315a974ab54b1cbb0e86d19e51cdd5d6cf07a031346b976c9a1e22b6df67e130f282a048d354395207bf4baec48f4bef124875773f54bbe6109a3217e61bda461431ad0a9f566bd247651e9e71c625bcb381afdc450ea377c4bcca339b09ed75e89f3d77c95ebf426cb18849d16ae626516db483a6517aa24f36649aa3dac6d362024cdf3d14056ccdee520ff96ecac00206e9db1da0add544f6db85741d194e62817d665969c204f776838ca9a2b4baa7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h58fb46ccbebb1efa792d8facee6d6bc4899583e2231c8cfea6129b152c25a2f03185800c3010684e3301a5247ef273b8057870ed9f6d30a5eb5e29f858d9b9088d39e839791e68331de9858b2b3a7fc0c3009503f7001931c007ff144af2259b5af147dcd3a7d7aaec68ce0d802d9dff371d9e59c14bc8c4b7b8c25b94ce4c5bfe07ab5d7270b38bcc0efbfaf3d17a80218c9d97b190a43c7283be0dcb151b7952cda4321d7b23d432d3881266717db96d3eca1e4122514a6a6a28551ef966385a6e15dec229ffc0d8b6a0038a13d92ebe3aefaf57c0c22f2e919ea396341c46c98ee3eac21b21bc886578a3000bae78a29d60f32d1694c32414e81638b66d39cf294c8a9e8e8b938dfbe57f01e8f4c5a0076846b9371188300e8bfc84a6b4a6f3cde7d6e37e81b02cd8a115c117ebec2dfdae4755a3aa8750e562b3e3d89cf7daada1af8a139bbaa0790eceeaaf6ea4e0375b7071c4ddbcbaf3e01a535489a0df4b8eea019f687eb21d5b3b4cb975723d48cbae3c33bf3c7484f43eb0eb2bddb428658c1cc222a7419d8e96e0c11fd8a4b54c0bb9aa2909460937a822a6ef1fbe64e08e318baf09f410ee425f6f2ed2435d204ef8342c4c1ed91e9f3896723383601aea30d196c26bc13120fe175cd87140386cdc35a7c44f026ae3fdc3de5a1ba890caae9e6534cd7922fd33cd90a08034a696ceba4d5baffe7e2b5fcff9a6d320e7b1621d948cef79d94a58dd358e3764a6c01ffd45f17943793988f7b88c1989ac6030682a05653df36cc4668fa2bd18029010560f0d8eb0e8bc7ab917a129d3d2578ecede986f47c8b84a7f89c7d740998374637e84ac55fda9d1e0413fe552ec8835d7356faff4c1b854aa803b9c06a067e32117e74e8301f3653de1b45c4b885096b68c69a03495dccef1b0422efa6b52413f32ee4e4001d149a4f1ada8be1609016edd35f0ad08bd6ee3f2bee73da55b027ab1658712ca0702bd7933741e03b04ae518b9aaafa2e5ede1d346ac4402fb498f12816c149c89bd36cb39b2086ec9566ca4db72a05b251c25f4dd97798091b4fca6177042ffd6521f0a2519ac0f14cae1213ea18c51f3c878e91023ab8eeae4f0aad7f86b7000752d15386ec3c2498e51a7ffb9e439fa9e3116413f7a13884af3a5e295319ee9dfd57f5ef416ed6701a9cc733bd136cc338e137a4f873ce3823214aaa3c22ab669c975e95108db0a0523073158957f0e36760ead273ab29898c370b35a450a4c46719d38ea817fe38a42ea4b8b187fb397f3eb8ff3679cd5ebd7fd3b05a5571a6dc1719780f728b7fa28e510b77faae62a33f13111adca50bb97486a7b0fc130bd0b4568c2d6a88723b9a7664f3e5f01f538a7db18239c1f58b9e4e4feb902b9fc7780c4801658028deb2a50a6c53793c8892cb6725a24a2cc1dee78551b9f47e1f344e91520c8c225375c01b7decc61082af96cc0c3c7f4c2813ca91e79209924a5f705a04312e8f4d742751bfea57e78128d0764a81e09f0bbd01ac7bf4fc84a9f6af8e0ab9a6a58b42b6a7aec34e1b61841a8dd0c5ccd908fed1e5f5589667e843b314aec1351619a0f30e9814a849b02c0254e1fb2ea4ca4e73005cfd1113bf9ce814dd5e1cf6180c4aced442d88ee6441265733fd6af9c93ba4081bde28000e9fc5bf7fe044ae7cac689b18235c5ccac39f6d896ffe8fca4c6b8c3c315b98820bcd1b3f4cab464eb0d7d403a7c0af1f0b06ac9a3c869634aa3959f969f04ebefd6b980492ba47d18357504323c260bfaef9ae7cf301ee66beafc57ff4fa6e175bde51b4ed439fc4e98962d18ef58b7f705bd7f290d206f8e085af29ef1b3da8d0eae9bfd086530eb42c23359394f927ac42dc59cee65eaa931a19a43e379fc522971016176de014667c90e8d7e02e76b3e35ec014404a24268abd8eeaf43886fa5ba4f2d8ec0fdbb81b10a7a6e15abaa3d65a86fc080699adeff28a84e10c93d8ea8dfb160814966c9b58f7e81cbcf16d6b7888d06c37df05dc68a09b150c6c16649342a0248d822ab87a4a5b54dd9b203740213cb6fc185b332c4b564b12954ae23ab854a800940238480b3c3755f6912f6839729244749bd44946c936ff9b151c71c0b5a4423b53abe41b1ac67e3a717ffdd808337c27c89b35c0abb12526f3dfd24d9ae6f0f24c8836c2f621eb6fccbc6a407d144c2b76bd81912165dc622cfc0917b2373143de16dc3ec06220182cf04c427528681a3bffe4fb28346a9a307d668f926fb6634e7b71d30fbf136a13c5f94147791a85ea3065285cf9bf730cef28b8dab3de03f5ede459711a1b845915d7e494160b64cae1cf403940a3ef6db84471204368d4acbb2ae6f1145dd7e2a59dfff3cf061a2179524464682bbe386147e15644885e3bfae69f424094ccf4635107b7134d1fb2c9a3671cad0c5b3f03c3c5d88b2983e5288d476346cee93c4b9db6fd2d43a48fb4641eaa08453c5a62f519bffad2aa4644a65b503dbc709b641d8a1e12450dfca8022a03a5e7fafa94d8d67702d697b7b12bfc005147d03d89105a4d815aa25ad0f27f3c9a66fbf5ab37f9e314686639ec4aee5bd64262cb29913d4103448b6e2148c4e4f836a55dc84672aa1a1a69c47d371266723463fa542197d6c83cc94ceda06dcb4a0ad178515d4aff1a4d550858e9aa6ae82aac4af72c6ec8319f09ed0e46cd81cf62937c0d87f94e46ac7fce743c5d6a751f4c6ec3e1fc875bfdf9cbb54c3dc78f6be8b81c683753230259f5c94bee1bb77ddb0234d98174fcaeacd6f8234193086a22c5580b1f14957d033bd9ebf1e9bd8dc0706f53564d2577f16a9659684565b61c838c7b8dd44e4ce661aebf1bfebeb2fc09fe46f82021d5b27ba05c64b2f652c2c717;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h76e46cec926af46a0f817edf72ca56175f21706de2557eab2ecb4058e566c669f77108d905709e66166274a6ba022ce08b20765ca11f676fe1c0c63b39e8ff8f0a824110280f4b17544b749a34aebb2581b1006f369514f173cdaa0636c68904226db07eeb5168d04a837aea6e5602c5e6b0fc7626be05aef1f09b0bb32808dd0ce1929d78aebcabce4a9f0f1846799ace4efb409e0185622692ed923eb5654c65d3f5e294a7d3f51d6fe9dfb1def8205ad6f8f535e156de3bd5c3d0935cae572f80b8d638608063bed7e35212f00b0d3b9d4be02dfd18c5dfd76c648e577a1a6204dfe3f0c1d7c9e96fcec6269d8437a0a63f439a8d1f0b90d84bc79f2fe3de6c865308a5f54e4e063a11ea2ac80242e9f8799b5966283bd2581cf7d199456329d6e7bbd047ed02c7ef08935a9cdc4765f3659256603acb29c80e7a7b315bf4c5d36f21d31a6894b21cec37468b6ed939a7b85d2da6230c20e99b40446f8827d6243b24a85b4c2006f431882938e14e95bc703e08965109908617fd2f132deb2670b2f28b75a92e20b48a98acc9f19652709ae4c64cc6fec47a1ba537e8f62f62b649fb8f2f161c0153104af220d009e862527b56c5a6506064d2ad5792e6561b2b8e31de3f610d6cc3dbe4efa3fbc771c8b1c75e4be2dadfcb9bc45a9ed628e11e7c82f7e4f8e6150736412afc9f146c02c7adc40f2cb8a29552fec3402b1a79036a0fbea898d2b43487f4b3c4734f928cab4d4acea03bd8aaa17a5669c82aea8e478841fa30d0f45bb1fa64cabe7f88b4c8e456de995af4f4c23c781be091ee24957156545f415e3efc377d9c4b6bb6866f1f66ed8074ebf4beb0a14572b72f1fc6db1f0698279fcc8a00f9a3c849a512c27366d217e810cd862b3783d93ce1933fd86b592cf333f666245df732b8798c8ad900297dcdcaf62836baffaea750c12c2ae2017614dbf6507eafeec7a498ddfe9c9635ba11a011c2bc794a7d48f0428d944c241b3e1e42b80dc1338896b5f771e0de82dbd6422065ca32bd0f42f837836cd17ef49b89963e64184576476153bde1daf51d6c32de880d01827aaa8c3a131fd0ead4ea2dcf41a216387f4c80fa2318daf9ee9054881e5025da15e0faac03ffc329c60995373c2f452107bab04bd362228de6b592af85066d054c444bd36ad37d88793076768c6418cc03855b93a11ac084f696c76d4bcd9c63106c5229a8b7ffb8ff817b254a8fd35c88739895e16f3828359cb1c80383b8a33cf7cad88dc056eec631f14f2d9575055d89ac61152ad17f58f91b6269cf37685eded54c62caf5f1bcc1917c034bed3a5a1a2afef8d9599e2449932cd06b31634d941c18678e739ea521e59d3fe162d004eef9d068437c68be2706d2517fea08cecb8a4033112dd6590585fed00479446d406da48875f7b2556e2b372552c8442a1a4b434d4cda0bf29e088567ba461874e263a95f2de5de84724e5caf00d1456d76c4900a6ae0db6ba07f29a1e561f432b59a169b3ad24bc5f876f35166f798428dc79f91c0de3fe0990c9777f2ba8af534f53f86c0a9107982e930101f611682a367d0b6315d0345a73768cd459f34d9cfcb8d0cb1cd6c051cc9d988d17d1a62ae400f9ca8355989ed41410531b04294518b8c9c1e524dd325dfb8ba1ec9db717de7e1fe055d978638d2312831d15a2e175b61a0f1bb3cd30b3e15188cb99a300e43e06608d10d932c10654cb58d3b7d7828eff1b8119dbda8018a975a4747ff2dade12f1af39c6c9da5c07430aac78791dc9be9e94f03934935681caf94b9ee3734a797a390f40c4ac1184d0f6f74e16877e53a9f874fd3d77c3b07e6d59e2b0396b24c04b1ec04887a38f6c8550181fc47bdd7356d72e9af07ba875abf6a9bec86ed0a8b2e811c76f794b09fff2e2c1ec4835db9df54f029b45c9d958943dc1f26c3f248c44e996a53bc4607c61737f052777d312e114908f1a6a08f8501523185165929792dafcd96728cd112cd168c8668fe3ec7b1db8c9802ce7abaf8b6b71dc228bb954c5ac881e2e1643a8588c15a47bd93ea93ab8bd2f55fe5cb9c5fbf21ad2ecc145eeb0c277a643643135b7cff12ce1af0e4d1c495968acf50ac43deeb9452503d1401ea841fdda59a7a19c1aaf09605b7c4f437e55a20d779fa318042b4e2f97c5623152ef6f132d88fa74c99d199be85038ab913f64e5bd1bca17879e989634f1b5d0a811729833d25f4ca38e8a3af52f00a4a35e6bf0dd2abb83add2dc2e59938b0497dabf77583c2b48c5ebdc26762ec72fbbff8c842b5e6bb81f2c7e058a672810d2224fc0f945eaaa829aaf4cd27ffb6f35aa1ad8ca33c3e7ed99eabe9b5a8e3d7fad137f241213c73d4974f0a065c223d7821b0218efc0cb0dad66ebbcae28f539edf11fb14a43373a6fd991e47795e211c1e052dfc9e2f3e3f98da522c493639d144b90666621f64eed01c42594867f51e10790e30cb40ac149a4bd32deabf32747b363709a1487d0466ceb634f761062e12fe97203976a83cd4082f50756e5dfbfd9731b9d24de458dacbc655c45503da0965369759168915a328719c3e35e0e7b585612e567b07fb46d9d17781361c4c5cf6f54ca2d563d56701cb0b6a5e27741dbaaf24a705405b1c3366ed322fb8017c455a639e4cc9a8551fc39a7ad5bb1aa28b7da5b2c07a13bd21e0c4c2bf31c13b33b32e68cbe54974507e5758819616d2d7ac8d7f73660f0a513dfa1da2d63ad09ad78833df912a563470f6671040fe75339e764fe7e78de0d9131a414c1c4aff25eca434a01b947f2a043c0e293b52d031dfa3e01eb6c463bec5491159a09856e8d9d7c0b7f7db4ea7e62031709de9fe5f82fd97a529e41eca5bb40f292537fbde16e9a4d384;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h40db417ca9156153cbd0b743cfba5c5e3211f4c028f73f06614606e597db380b7e81d08fafbb0b37e0e0d0c4ce84418bade086fc27ad0d282e439a3c508d850e9c3e613f1e5c3e5cc27f986497f73314c7e62b822f9ff61eae0f3432d4c43ac9f4c2e3939316ee030baf698422370004f0e6e3d8360bfbdff60020d1b5ea2a7b4fd40c8eaa24d2ad68029e3c2ddf3a33734acb7451818492fa874a4d94fd273268f6cd7760ac848c6bde8d3257c22f4e72b580fc42691ac4950eb6d5837f8231953fa0d73d6e1536fdf1c1ca8b3824b752c0c1b90223e7e0d449caeaaa03b3aac1f7d025ae7506055c18c5156ec1f33eab035df8dbcd6b987faedd90afcb918c19964252b0ff8f1f8bf8d0a14c1b91eb5e9473ec94b2c1403599eb5d8e38b3c231e44c32f014425c6459caa5227db6647fb1ab3a70de5c3f2e557a79f5c56b9be3ac44e9297506d2d585921dfddc476044a8978c24caefe7ddeb73644ca6f307e75216f251a4bc3b8f0cbb5637bec063df5cb720471859f5858df31738d01b94f237ba2340816fef262d70d4d4837277fdfae3d24586cfb817236b2caf8cedf99add292e2e9bb2fa16438dab4180d4918701223f318c74e14fa89c500f8a9be16e88455c78ba600ddd6ce401fee2c7491eeaa4d6db2bb3b8a481a646e295effafdfe0777a119d6c10061a74d69a70b9f4405d9335a3d61d0e768a5f786f85873dbafe5203f244fd55b8c6d88bb49dfcb58c6aef0bf5f444896fe6520995610285d4f62ef3e1481759b411e8fd43a955f08de739fe66a677c2bbb5e5ee4d582d4ec070b3e8b01ba4b38381a12f2aded143582173aa3caffe92f94a16ff6bbf587336c2ef074c715118729f6a204678eac0f0c89fc0c63da3b5db398496f101ea424af6e76c1be7854cf8dda0b07703ace72235456ae658844b5f2d62970c4d9e2fd1dfbe44a5ddea33d4a2817406c4df1233d4c70616744966c9b10c11a0b59cc6dad520dab8512972bb611a851d08e0499c5f8cb9c95af30f9a4f17929b6fa989b8bb7cb59daa2094a2190958e589a24091fb60ecd2c9133bfc3074121e0b154107d143c6ec14f96a8382531702789e813ef3f5eaad1e925154dca61ada189607b0f00aec59283cdbc577bd298ee96760fe05301751e64b3c288ee80fb6acf56fa9de13d38197c74553f6d2dcaf0303c58effeb546f94f023ebb46efdf94cc3861880e6e93227f9cae56b837cb3bc2917287452a43aafbf4ce4e9a272aa249ca6fda670ea340af169d0dc250ba52db3d1190d8f6ae2b1c2c7429387bbc8998113df40e445278fa5663d57dd9e5f996e21e9ee8a9a116b2f7cc055fdc1a123e4cfa706c8445885200c458d2248fa944c038c958adfae9b76a5be85a5762949ae03e09476ccf1cf7ea9dbe3954bed26fc17aba3785e9fb016730455bfb6a1082b591ebc3fb6255f9571dd9845d3e1b5231c2bcd419185e17c7eabebb3b10529e4800c0bb4c3cf02f702bcac1c4e10a78b301daed6c2d160c0cb690aebddc7078302a9c623cd453985714d1b5628d9e3bee2af236515d956b79182d9a263ddd566eeaa4b7f86aa232de399a8671e0e02eaf77a654f88debfe8d948d63f5fda30bafe94cd4cb7f0debdaf2bad66d066caffd42081b39eeb18eab1509cc1b949c2917b86d43c17c671354c02ef5d93ed49514caa0fef913e496103443b3f6a3a9f652fb2813b7fd3fd35cfadc210efdbdfd3af42a184cc49081e77b253a95c64e07605dda5ce3a91777130f4ad8ffb7773a7169b53a0cdba90c72d9b9f1240c4d5df61db74b08d62e9dc6aa336b7913e3660e7dc3163826000d92a763ca475bdcd2f0fb5e582088fecc0a84abea76fee7d9c614f2cb3105a27fea9eec73196e0aa819e4f7eb1dca6e965f3228cc67fb1849f6dc2fd3ec633e4847643e64ed6f2b50ed3ed925fb3fb047ff758bd35abade283774d9206d756e5ceb17663b23eeb52ec2cf23a9bc949b557f89fd6acda7c033d9276a66039768d707a032d18d728108888ad568fd26d963092d71d4b27186cba4698ecf360363b6d87dce99a633309f56417e031904fcdda7a810f56a82b87e5b048147171076dcc8797b7688dba5c54592d981cbfaf4be13929dc2e66de1573d645be001eb9b18a185f2aced986360075a6b4ddb72deb92c648fa5a92a55d7fad497b980fa7738c68fca3698fd5e6597c2b7e7d4150b012a84326eb6de8838cf4362fdfa50ae3d20800c78ceba1c64a0fc7fb3977ff1cacdb408f15fcc9bdeefc6ab97b473a5608abe4cad9c788ac9ccb80d37ccb678d395392331de16f581c037293571f2ca715fefe4a88cb0eb6123ac611bb9bc792f8f4ba2aeb1120cfc1522bd028940206e978144a8bbc92d0a057cc52f61bd57a40c583c667aebbfbe1b01035301e362e2107bfbe61cfbcf2f64bc080ba52c61f87f1a0b8e5388175fa8b9d4fd98df55dd334ab3a7a20cfe23d889d041b7d349acd0bef97bec2af991cd1a39d5194defdd701ecdf78d3a1d6e1c0a631b23f7bc0a87b211da03ad43a4310eab681235be324faaec9e6a24f91b843c04162326b4f4c301578085edbbfbb7579cda6b3d5b0c3462250f6346af65f6a06796ad4040b956727aa8716cef2653b499adabe67e27aea7f11cf8dab202ece5d0e30ab1a1febb510558b5e947a9d972688d272967d4fe91f46d7385e500d07d237bd109d9ac2939389a42a7db93d3560f62e5b69b7443dbcb5b070d956161062582dfec3042c76f7ad73276a4bf5c0ba6f90a731dc79322d3db66a61b40a44b106804c0aed351ba0372af794b42e9c4bb995a087971a6e7749fa73e45a70b8ccf421eaae1a772a4e64efde83b7feab6cb1816f99893a9f7c5288e9fa40464;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7d1695bed0e0c032a4042391e0d1f518725b666dbe9d97adb95b9329539ebfe3f2424b4ff8227b485306607ccf22d22389cdfb48f6451e3f23ce797d92686938fcf790572e492fd8c51cd8a43fa5ce397b174c3741c89dcf9237feba635ddb947841deee3cc5e77731714e0773994137fe617dedb4fb584b93ee0d892c352168804d078ec1144017fc4a3c8fab5cdf0f8c28f3b299bdfc04843d84d2687e65cc755841791aa286cdc2463cd15ec50a386f654b08e8b42dfec83bde502e3457ea86c78cc053ad5eb3903b78f1a31f3e64d8dc0b71ae9130ef2325b35e3db54697f7459ef86b5e4c4330c507f269819e2182ac7d1addb1d9885514d9b95e636376c4128b9dea24543d5d81510abd2b62183963d4929a79ff9d82ac832b3e674b39be17570bd86b38c757280e04184b6209c73046b69a555f84ef3b058f47db03e8dd5f03f7a7bb49a5ccebc5d812eef51873ad53b4fb536eb7da29b27f78f4e87c855918b7ea7426fb53238f8cf4037fc644cd0fd0e06cc4f92f11c3b72f07860e6f71b98590a74c62d9da9de97eca88bea100dca5c0261d8b27e0ef32f5764273da7824a18afb272fa02fe4d3f0efb84bd4171cb5089ac4e0fe64b42156aae5f868da52796891666e20532cb215f50e9a29c2e631aad3841bf0473b8bfca7fe53a1e4bcddfc366b0e7e643d1710f2d4e0cd61b2df987195f84d7d28dbfcfa1dbdda5ba1beee416731c9769ce0a63dd1f35fe577e14dbb35033822c115e9db9bbedd95a5d2cc1c7cba74997fff083a30c4e614f044efc0e4f17e16161a01711c736a8c18a5366062d8b29d8b5b3bee438f245928ea513b5133b8e9d92610b06c18d7b0343040aa104fa0c071145c4fb5aa4fbd29d8b5b9f5602cd05736dbd44194d5c6361016ca8217e578b81da0f448ff731968a4e2f0f33e3ab9e8ed60a5ac47f91cc2bf2b05da1c32cda8e3555d6489d198f9e0d251cb738444c9aeeadca1de2bc64957dcf59085a6facf302766de51b45c47d8fc939be8ed0fa5e9ad2ee3d19dc9d1ae5e7ac995cc693d9da07677350129207351e11d1be2a0aae77e450427ae269a84928e50569761c256e9f651af82b8451df6ef8493f943595d155033cd0334a638adc2ca90f392c823880dcef6b5570222aee739491974f2c4df661f22278cfabfb8ae2a9f9a4be256a8f7dc062180f523df2b4d75924ef4ed604affd7a63326f1f59297617de4f2a215ee70fe662cd9957a02f1686b75711c0cc893edd6d2597ee6ef59443b74ad356c94ba83d6d7ad7e1f271fa6874efb2e8c06b19ed27aecacf9185ec690ef110671f620d88b922c82b47345a52862c039ffc8402307fc0263eb2d7695f3ac6a6fa3ef358e59065fad841371c23222e856a5933ee3f7402ca138d69822c105030d5d5c276fa2fbe686a773bc59748d3b8a5d092991a4c5ed652d2172eeba7cc740efa34f64937cd13d3e0b6c89c209dc96d331eb7a84be5e5beca55210da7f4601bfc0061a7155506447a8247fb224bd1013c1e7954a088fcbccc2b7b1777810a10fad00484e2d0363c87e7d4754060b7f1e18b634506f5659d4db1f4ef2152498368c732952f7a149cf13d2968a984dfd2e9034f7f87a53c686f742deb523e601712bafa9256d4c816d9b757610311dac862b87a2adb7a356e3978df1b21a896c8e64add6cf25582e87c24fa3e15b3bb21f82419d8eb0bfad159b040a636947f88f108f7c4f686607978d73d05b4091a945ee347bfac8fc617d754f3a211f8ec76d818998f184f103253f247d4b4201023b887eebbca2baac09422b56352fc17ea7d03975509365a983da002472922e11a7daaceb2166049beecbddf6f8b21615bea7e9763eb1f7dad1eaf2a4fe7e160ca6ec215a0475df7d5a42a464751f08531bfda223431015bf7d87ecf2e80c038724b7a66cb0fd654d39c943212bdcec97c37b9fcbb0991a35148a4b70955367a5ac0584597c05cb628356f81f3eaf4cf101f1e133f5fa4dbb8bcd740bb8a9af67ad22a300733fc1b78dac97b0c32ef4a26452a4b50af0e82a63f6e7d3410abc97a915c0593c2ccd702f917e2e358d3dc98ecef2c0c0563f0d7e67deacbb8ce3f61fc58f58d15e4778ac655697f72b2916ededca24542c4d4052874d3b29a17cbeb9a73c450f80e7d640cb7e3d1f50d618d725c62d1ae9ef89c3d7547201b81384138368608f02310f6f63faadedefe152b2393720ec72f64429a19cd05f5cbafb8ca28f6518db2213c9199a3115f62d2fd27a349a70cd3028f1cd5cf8f853e2997444c7362fc6e18ec4fa33c08a908434ab634ce828ad0b719bae3f48bd491255b265cf808a896ed1d8def61005209e838f4ba1658354977c08e28e488f879afadef81191af8393eb219f2c496550676cbcab0ef1f1960f75a8c0be7d9ecee524eac6c459d1edc45d9421aca8288c9b94b4286d73e4b38baa0e1b5830045392499c2427f04237e6c9502510d3710efd0fb0c842091f15ee03ad293d6325a1f3fea2598d6f419c31705f38ef0045f39e62cacc5ca8ea26477b76208a390a3ac04a82d2c1491abf69586c802a6e07a64e7b868fbfe07b4eb200630f5cd1f96002345d7e276c6aac51521acff3b636d33ebd3526f861cab958cea1057bb6c4b9757eb509393ebd768f869521a23a43adbe0bf65cc52f049615264d7d953714478db6369780a37029b32d0170ec5678872ebbed307c7b7b7a9f7c5d9573d0c444da98059017f80cf787456e93ac22c39d967b53733f0a13e9285c2026d769c0e3700595a47f7186cc560d1179d9c55e4a815d2b77951c433612838d5826806491d9c325b0e741cea03ece565911b3bdff292012d5c18b8c41c14197757f753189e8dc3408f3ab;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8604afa3c5ee48418db60b499b26d17a57238fc8e22d57f89be2dd0b05a9242deb9899a31a0e54e3a9bfcb0c0709ebf6ad195711e67472dc8592f1b81e6b24a536a18365b22e1448d00a86096d8014a7bfe29b85b017655b34717417a5cf5a5fc4720fcf5341755e7525dd8191f3b40d474274ad451b2969b8370a290f0fe9d9f14edd4e35054439d3796780f03d861006afa1267c042b92f4a67dba1b99e8be41c8852197bd2fdd5068f5cf920bd65d640e2b4fbe68394c1939dd93eb9e5318492373189b3844c2c9515da190224d34efd7cacdd663bd218bb7213a0f4566351cb18e8ca7fb4694bd37364f38064b781f66d2a7ea4ae2fb29bca7667ad4792fc21318ea11ad5900b0bf1b336b83b5672c9f796c5c8f875c02a9547cb0195ea4fa98c62251548717ac33c29191adc5a0cebc003e29ddae0a79ac23628820c33be8f853fe33b029a51b9f30f9a78e08fad7eb15c327ce67c5aa9433bae38f12c7bdd51351524bc4b91313a4b6b56b5fbfb15d4cc060e19414e1c960a589ff63658a86ff5f0f63aba3b202b6c8963aae38afecb8a7e34d5fa0ef593402003adf2b9f00f341fa26049a3d0f674e9e7c7bcfb112322c467d3b600cc32be9705b8ea640cea33f808d915daa1e76553bad974dd9e04e80364a6f60434bb0c1d5dbe2429280f35de6effa81b91dc5d1f5400069fa95014685627716fedd8dc6df1bf9e597bbff36aa8f1b4f7b870c1be2905eb521fc2d927e9794f00ceaade917a7afdddce243b63adf15859ed0c447afcd8e106139bede0836f829441259f1ed65949ed5ff888d837c934e637e57ef27cfcd10e5e2bb2b8af4c272679fa2573adf1f2d51cfa1d8a282418f13810bfe1a3d1690b5433a2dbf2bb037d9a20230c7f2ccccd3dabff59452c4c20779dfb4ef5cae069f5efb1baa88d6d8bfa590f2ef3aeba8a8fc805d3181d0271852e8f890352016348b883b9b61172d319a022680159bf6a8fbea909a137f35759191e9092c0446aea9d226da9e6345f6abcc083fe73b812c78d27dc5b155d031375a247927277e3d7f4e49e51ea6f5ebf35a2c55b5d74a0c24f28e7ab556a2cf4834e7c3153db918484a0a67c176807f1281387bca2b1690e7a35558b6cc98eaca4a0a6759db6ecf095d3bd3e1a81611dfd893cefa7ed2fa45a0b1750c8709b343f571772355fc83fee9930394a538d8c23b30d6c38b28b2410ee8d202dd969bf37dde4504c0ddd369714b8d85c422918189520347caab35b5e5631a5e1ddb358549ada6bf5b18f84f2b800987eaebc3a3bcb78dfb02ad06b4b2ed343665d75a03ed50f547795998a9c877b854ac24d44500ad9a526a04f7882bcdbdf4abebf64abe5f42bbb7e8fc24c302f410d9d24b9abb3156d6fbd60ca97e036b00028ef81c32146ecc27aec03cf165ccaa37796a5535333c32cf5d6a61de1b9db8e2a3e15208c7c73d44949b711d3aa1767b80ce1fee385363cfe24b6c5df201b7ad003216e86a8c1edd93bc6dc97aba1a6ff440580ef295757283a45c379472b877a8dfa666d8981169d597d20408182a100f4559a7b1a313e99dd379bc86e463987e71e8a996ad12b44cd3c0982d40bf4b512591b133e9bbfc71728909a4263ba3c4a6a7e8005d6e46aa6566a48f56b56ae2aded3b2060233884bdbcb4d48ff4538ce5567dd8dbcd29a28605f20ef5d21a87c0e54b7eefe38eea187cc5f6c8b36630651dd14c6c4edf7dd472254718a2dcb9eb743cfe211aba381b44fcc7c5b4566ba35a966668fdf4dd6b5000bac784dfa9110a7e57ce4538a5d8678446f12a5baf9530d12ea0b75e96653eb989d3f98218e7474874f8487e2cfdd28fda48fb138b59cfac80a4455d66c60dfc7b02819253ed0e13517cbe236a4ba496dd2ba847bcafd8b6b2c54e67fff7330454ef0ab4bc20b0e97c264a589e01ce8e9b27ea754c5393762708b8a5edf029b3bf95d6ae7a3d73f76c4a77daa071325d104a406b1b1d94715abeb76d6ce65563d15c446125f0c63cc62394f203ad6086be0bc2f1d5a1d8cee838a9e802daf7e78c5f6c80d06253d3bce3b256dac00b0b73d7d1961d66c2e8bc77993b00c001dd7184be4c7cd83c27bf8d8b801e0c13adc41d61be99e0852db7176396306855f1615bd6ae185161dc9b42919a16f82618c8db995daf1a03a43a7ec4983efb9b57c20a4fe21d372a0f52a02a5af0183e3364f814e423a2938b6ef7a7507d384e3344012a8a4e28de87100c962f72c94d1c637b74b767d5602a82d9f1b5bfa80d18db87953acd2997c51948927e4c14c3d1e31c7920d1ea2b68b3555a28e50b0cbd6ba61297302549afef2b35b4e7c5c80d6e50854d8b2b0d1e4450381d7bd26eb7a3cf2a5abfe051ecde4aa6b9a07c570a39150c2158dbdf51838073988cbf5e72abf565ed0190aa77613689555240aaacf12df03ce00c3c4133b710ce8d4f574492a1140f6f4e410ea74fce11c528c372a4db32c24a97d2bf8511ad3209f05af2ce392db6c1ca47d46627a67424dc0b26ee6339810eb67fb10a666ca19c8102273cbf859c1d090b148f654dc34a84642efd35e02a135ae48a63ce81fd2242dfdf8d2c2b08e3fe727cb476e84d9e5ac9f300fcca600e335ea6a79f02599ef64fefe0abbfae9ae645177bdba73fcf118961d39f49726e4b1c6bd8455b08d04ba48bcac6aa5a4cbe5e5d27c39c7eb0d70127038af58899643aef4865fc4b9fec9adbac1bbfbec84d0a79352158562ccffd745b9db2b95fc9f5649de28574428d5f422e7470a9a45fd0e36e26d285f26e81d7bd730c1ec2ddd0a8e70e7646bc2aeae1aa441b3fac8c282f55e77301c6e82679b719d4fd82219eaff4564a39f664082e24e980972b3a061c73d80a8ac2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hfc4030ad3bda6768f717e1d5e0730cb67f2b973113120d1edbf25f0c0a36cb9b6740cc0c581a2a14080b7562703966fae137237371a89240a62acc1dfa8c2b2ec4ac5655ad224b1f30466b3c59ae4348f3ec745a2b34024bd0a01cda5cd2e3a4e73e0dfe1a337222e00fd2645664f244489ad4cddd741891411e16c468dbac80fb81ec5aac9949103a37e64e15435aeb91eb28126572df6b71cb2e720a70559514d9e3c45d3bccfa3531b1fd865a44b6ee59e2e4672ed55d147993dc62dff2f7f4810b5fe09ea80f06260bac0591beadd221217ca367d0a14d12f72c75230596c8bbdbc6ff89d9e950fe4922d5c8da9158726552e76498639ad4816838811fcb6186586f6f601a7ffe3a97768315ce74920574734644680ab412a18b7d03cfcf9ab43f9a2874d9a1dee187a69d5fd45904340da96570515b0a1a3fdfc150bc7eda623ffbf7b2d2fecb8701344d67709852ea5214ac573fcf112883f3618980785848bfc7138678c4747295f8572d323b95d551343cdb1d18f9726a4e919739b22b3a42a86b4b09e962a6e54c80d1e7e84144e5e66e19b01234fa1b85609861c77a4cc04fee996a4f16bbb795bf7e2ce8f6df466f3f208348f9cade600dc180df01dc7b7e9e5a16f6e7a9d44a05198afe9cc77fc3beb11813164547ad44f1bb3c28cc4ac0eb89292fbca486d29d7fa4c1f29f31909225d805b40ab4b036a98ce0c26235a72db0c18353d26e2ed1f47ecbdb9a4a78614009520152a700aa9e750cbdc198b17073e2e28db72c80e80cbf7c0d5e48a40ffacebf06610a5fb21576bd5d518e6a3652ff0915a609f59b0aaccc97bdc9d7cd1c80eabbcd5e91b51b2ee4d581acc357547f6ff67b8de18dc59d85e19d8df748268cc643a6078c6952367f76c46df05620cf3a36c597c55f5b539526191dd12eed76b81f57aef66d60632d26ba1490f17a422bbb676377e6cc84d60bdab61bd8ca509da9d59e9dafba94fdfc2f38e601731c050cea3e456bbb7269fefff5acfc3a7ca5cb7687f01f7737927f8b4e27696bbe84692237215704e3546d1d89f0c3b3f4e06acd8de207a7256c4fa00ea2c79b83992555b6e4236f92fad7cbaab5987a608d83dc792288a7a999cfb13fe68f6bca33bb446c706211f89492edad41832db2b9311d942af98ca22f0f62f89a41644fdae7065573aa41fb65c5edabf01e9a6ad0f3f71fe61c2799ae49d67bcde13358f94d63899f23d555a128624316db203070ed210283cf0b2d44a7146fce0b3ef6d331b8f5e47c8790b08763ad1e514e058c0050b181a4cabb207c9fb3ae1fbbbb2b43f7d4121a1127912cdd44f6aa566b4b9f25256911fe8f0a4f893a5d519de388cd7bc93d6efe99b9174daa557515a30444c770ad6e4c3386fee7f53e1ae0b0b5892e6631a48d5ebb63d8610b1597f4c53bc5283549312cd7114d74e7170921408ae435546ea02561fe68db8fce89ac510166972346c2764051dafdb9d9ce719ae1c4db965b8841c866a82e53cd89c88f2dd83301fb49f0e6d6f281acf14d5c6fbb52836399dc1e2468d1b884a6a6d3847d75a5ff9be7c4b8415a23cfe1a1562f8e868c8bbe177d2056e5820114e21594d66b059a384fe662d3bde6d11fb2d3b4e9833b78cc5eb170e3bb6d39fb8e5fcc573dceaf4659532bfe54b101cf452298453346fb71be40401b94862c1928776c0c3dba16beb86537373cb4938be72fe2c7099eb1bd37a246b096dead62c41267217eee59c35b18a29e4d3dbed91293f1337f7f7d3d5ed4fc48da0de13c37c816877eb37cf9145e58dc7be86c665f33f08aa31dc147c95baf20a564a40fae391e4da25c582d775a7a7e88c86598b60d20d35f4a9867af81b7b7f952126400f34e9317c3b09afcb876073855c95ad5c56640f4c5ba1eed33e29607ed5c9a9febc9f1b5eb7370b302f120138b20f71164b8c9f84cbb47e2a2e4b7072f6c5cd6b76e448a9251ba18aa5916818e61e87161c07bbff2fd8275d27c4da80e8455d89832c8531f69b5a9941b66fc8a9ea022d1992844c718d35c5774676d7d9d71e1c5416d5056c5f106557b1d1424031e073473260bb01a3897bc010c7870a2ce5108c0fec78619916f01a32259a01f6d995a3e678ab3a769cef5861813cda3085828f46aa50babfe4fe1b480aee4ae9cb0fb394a8b42b0e344abab20f70ce0a489bcd7e7c3dcf980d9a5f0334c5731f50bf99f1b7b81a0bcc825f621c837a24ef58e3f5c83f63f14379216567ea9fd0632f64a48ad884e2b90e4e21adc096891e7d20584db595d8f34414ad5a6d733e78d72ec8766dff17329f1e2be54ef44b825d734d7f2c7113190689c6ad4f0180b9e3db1e7358738730e18a3b219d5b9efe468b5d6a30087b627760bdc3bdf6330316934bfff180ee9531d8fde039ad6ba91148e79928c77f04913f9d986beab58f69ae731eb225b1c68e4125649828bdbc8b6af3265b7de5b0deef90435dbe66c268cb8b38250b47d535237a4d5b1563a5be5869b9263638443a9a78a47a3d2a1218b7f5407de3ee3c2bb3bb5faf600914f92c36a9b335569ac890fe1402bd9077f488647374ca95efb9f9f179005eef01552d7ee94dc2201e4ee19184a44ed6aa947d994715f67de8eee040f96e81dca7fbd52b5acd368fd55534523fe079e3dfed2c1f5ecf63d75f61f084f61e126425aaed60dc5643b6a7935ac90f32e887512bf5812ff116106d6dc95c190fb344f7fe5ca5cd7750198272ed3dfabd7a3d4482890305b298fb26f74c5fcaef47cb25f2810723ac704dd003abbefa071f1bdcdbfbe57219ecaa7106975415b99b392e18a2f0212fd33c293ba80831a0da503b4929404093284f5ecfee7cacf8c401ad61ea3ecf1d8438cebc0ae;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc88c4a6aa03894ba5ec9b4e1e1c3e0a06fac905a99bdebc36e894aa83be9f62c6c9fcadf943f200258b48a5811900a9794ed01fcf9236962e733e660676168b6104d3b62faf971298b56742c181164ba13b119c5dfd74d9edb50d6dab987d2bb6ea598e4585c98310fb8a190ecb2be95b286249c44c94eb682101a9176a68b1ca646600de212a1a86f5132e3d13e40895a7d3dda585be3259facbefab340b8b796082aef9eb44096a630f1cad8c4eba18e50951c1c668622ac394dba379af3c018b6ab3fd50adb0592b2b906cbc64bb8f4d8356aed9c57fad117ed8612ff044f9eeac5af264da0b7b32c2a83f6a05b8750aa1ca223ee6656ccf0ebed89fd03eb58af22af89bc84a4feac8fc161f9f0a860f6a16e36824bb6bbdc700082f5373b2c2772b2f5410634d2c9b3400b6d232b581c897a962689d199166cc8adfdfccef8f91632d1d898f55bd07338dafaa26601eb4aa3e182c400c71c7071d47acc4347a1b912b11791ef5804e11f3ad726d9f709e371d7a191a391bad9d4ec0096342ffd9f1a0549d324f5a0a38dde0911bdd68781a2354da83beb81b791dd8b709e2196362682ff5bc4eaf156513c22a5d5bd77d25ed6eba73676950ef068c145b01b708eda2088cad66ac0108ee1939ebdc82c370d5a900008facae34949b075896170748041550db36383335f0bcf581354b9b99efda38510e9814c419484c94a6863cde3ca240701e93416cef26e8e6779084be0425c6a8272893eaeaf7e62a22c1940d90b31efb50d9657b678dea9ed597e88d0d5573a6902c6d9d7f867403d41a8f2dc70c32a2257d33e2416422f2c6c583e8672fe276577d1dda3b7a20af489da4924a5a131475d49960dc34ac622b63e950425e59acceed034a0dadab3b23b4d5d9afa0c926aba66f0213f4e24ea1cc09f4962d5b17c9f77c0e99c7066e3c6263da4f5733124b2a4230dc1ee0e2815c8f7c5ae06ea4c328fb40dc835739a886cc235fd72104ccb95b4211cee0efdee60f49080223a79bc787292531ca3c4107c6dc16c13cad12aa361d9fdfceff7ec1f9c18d961cbfcb5edbfce99bfd7bd31a4a6c8d3cdbe0a73d23334404f13bc3cc53dc86f95962b0abd02d10e3d88014df4725fa08a7b9898b208265f106518162969b8908db87d87126af3a133b2b463f62a463ade93274ea68a547b8b06346b49469ac461dac9d794cdd72b1f5c413f6611ae47db9b10d8f9d0d5d9dcde5fb25da5ade56391a0500f2e18525a0d597e59dd8e49a6d46811bd482a860af80bbf0ece2989ba09b062f955977172093dad274f394493059e9fd4093cd9379ee2ef6debd6e9394fcb1d75d108456ee8e89749d6b7fca30bdfa1708674fb9621cd4acdcd01dfb20e4a3e0dc4c3d029f5879ddd808eb87ad5df41f871ec663e4921107e38650dc7ffe6fcd3ad3bb5692e98e4258cbb3e414cbc60664d058c15beba9299c9dff79e95cfed1de6c6831928cd69aa7e9731d3ba306fcf9f02f221461dce5e68b4032d89d59097352124985a51e20c8e8bd97c3b6a72d5697dea63303101ee05a06ed08e7e27903174f19de4010cf9fd42b2d19fd5d3543f2d15248e446965674e3e299f94f5058c5dc065228f1c2c9b1d340b43ac82feeef58c55f5e5719781e77c1a75dac349b7212ccb045736332b507eda55c11d1079d7352547242823988b05bd7f3ffe05f99e0e1ff20e30b1de7e3ed581a3d99d02d0b6abba4ecfaa0c6bacddc597865584fbf947e7105810da7d2f952179762416147870cf4c05da1504c50195920df087a4c30c1229389d5e64890db2cd64fa61b3b8404f838e3b7b97d5e386bc08c14b0e29eaa4a0a4e7eca2883562f95f86ee6f66b9d2a0a6b8410fc92bd332000617c6900505a12b1e63e1067f77cdeef29e29a515b82f12f6688ad79de955beb1f67bb8ba376da8c26a5d0e3ffcdef565d2da77c2b9ef3b4b8bf4f8d116c6ab0e6a48d504b70f642183f341d591f43f42b6d44e56b87746f3c9874a003255f8f12ef726c84ca81c5de8c829eb4b7c17cea3ee34d793249a9f2fdde63e89dfaa9fe73b033da0fdd7a23051431da81fe5bb02d3d97b768a32a2747e86509f1efd21727c7b9cbc88ad1bcaf184c0b62d533775a14d12ba6276644a4e4377b4a52d8a536fcf1276357b79ee7ea8a86282e09accdd0261a763049747d6f724683037624eb62ca6884b82f274d5e70323ac568000090a512e21f928f3528732a6ade07580ad03f6381670b47df27fe9008883fd403e014ead349d641578b2364ed68a83554a392505cdfff45d7fe3589a71688d213e7b4717f6a69d81252909d630604e307f68735b18367df7ec242fcb9a6f7a9b1f588c044eb2305230b5f4de5a48fd2694783f878f54f43eb662e194cbcbbf5cc36c2ddde352a0ce283e105091cf145e833476b07e79f0a7374898033a3753c528dd16912666c644260d6d299f62e879d68a82991c5115bab3706a866702f8834bd6be950934a1469d4feccf33fc1ca3e924aedbbfa78c8d7c474738750eb6ab8cfce8a6914dda8a537cf78df2e8ab8bc312b21b0cd0d8b1845cfa7e70bb5151cbe180f21f5afa4d63e97c9c04623f94d7daaac8858df29f3e945f7b54fdf1a222e56f220e78ea7d62ada5c5a88d1631ca117bfc2cf10f319c26aab59dc1e6e656f7f4a4b387907addc1be702d2126b5261fe1e80f2786592ef6a3d94d5120421f21bbdf54058bef1a8fa536d60e75ae12fb026b75a67c51a5560c9cdc9136e4ecc1cc35131bd05e4cb0e17ccdbdf9a1477e2020c9815583f141d2782a9b598d19741e630e1e2f1924f51b2b8cf51c7ca43277a5cf5f81425e43d96a019bd4692992b84816dce4373bce0fb843a63455aea5aa1f0b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4dfc34aacdc9e58eb97de25c53f813b29a983d541e2b00ad2eb38ea4533ee257ea65172529b007a0d56705a7459669a2ed69a772b30047e21e76b2f369d966f9e0f2a3121fbef5d45b146e4eaed83f726f84160c8fe8239a48912523de7d61c461625c04a1a6cb9d45bfc03c117b8f57bb2abad3793a6333af65a79f155443a249b8870610ab8b1bf845d52989db1b8b329228a273f71bf81a0243f27d772a5b5c546a36f0bd6e28517a40430327303efd5b1087a89060a7f99281d251308afbf1ba7beeef23c3c0d7424a34ca9a30e46d36a8a696d168a8474cb55dbf8e07f3a8df27bec7f8d43db62a0c1f1fb5fbda7034c35af42c2bdd973738582637fe3907ffe009000f2644bcd8b10876b5adc2c13ed52aa9df63ada2fc7c6c0b5b5ab110abb8009003569e7e9369622c838662508bd22affbf3c86a039c27843319e4434331ce1d63cd581d07bca65fecba153c7868d6eeeca3e1a276d681dfb451a68b3e8f18b05f3015955bbe4f7720e2dca634c170cecf7abcca39c0daf35799b7cd0f7b2bcc2f7567e2c38cf8de037cd3561807e7c8e9fac791886b481b9f987a7db227fb23b6b5d79076cb56aa0ca496e2b70babc513dc927aaa14bf334bdbc62854952c3088e8fd650556b062c54883fb545ddbaa23766fd2b703b84b723744d8c97980e532c1c5021942ca571da7144d308a4910334130b4742993017489d771fa69627a2d137d98179606bd1ce00d6035e76c7e855c8aaa03e3054d946e7d2e52e9043a991d502343e99fb4cc615a32db3cffc1a991dbfcd9d84a65423d3ddff7349d336ba0fffaa32f0b44aa8952d1200a68a14f68892aaa6bc0327790ac1dd07fc4767cbd0d302ab02c59493e69d72db97e8c366a97c36b88f12366d2fd1c7f6e19e547b368ef84b94ea85e433f91fc48b1416c8a3961a1201e1f634d621f2f1ec20b42a864a6377f10486853cb279dea7b0085e3e81e3dab83bc1c75f9d77f2c86f934d56453ee26a87b288b3af6aecb182ae3f2c49d367c9932a253d163e1cfcfe8f7d15ca22da02d8e5ecfc074ac7bfd00c335eff26915fefd4b9fbba03e77771531f6c665fcb65e816dc3078c1523fd02b6c283cd2629f55114ed367268b0328b42278f69d1bac14658a00975484f0dff2f0fa3430d2b242e665a6bc811860a9666849759f47d45ee5db374e86c97002734d032e65f8ec3ee51c2626b1cdb485812f7c90d6e42e91a3a34842dfc8562bfdcc56dd91e6cf4eca011f7e4f0ac0236962ca572835ec0f33c97f8506dd5fb8b742cff69663738e160f2c21d81227e9354aacc7745fed1e9ce5216d071ed79dcdfd7b0376a80b7797232689c6437da4fc5de9f8f371cbfbb057fd589214cc862422ade95bd9289241a8d52c6625a7dbadc4c673b3ee493d200d26fa197c038f1555867a386024ffd44184b1d16e771e433f95357785b94488b269a21bd650fe5d3bc6fc809d59204ecaa85537a88b47865ed7d11fea4d524264cfbf6c23533fff0485ea3b4ddf53a2a208094357f1db108a3a2ec7cc055d125dfe344d79c2ddb01984007dc14000e108323ef8560e47b516dfdb05da1582d9635e503fe589cbedbe2205ac70d866849cd501ae021b804ab5ffe1a93969ae7a8468a62009542c085e44be0ac485c581ae6af45015c030c3831a28b7f3ce07e32521226f07b558747330e0163dd560fc35fa7bbce018c1021e5d37ff618c045f5bbd8073b628c8fe82fe442a7739e94000db0e1910c883f72e4bf484b30600a087526cca9fb724c5dff84ebb2e15a3c0df1634a3f80d403a505fec09bfc902283abde0e87eb469be75d846f04f15135d2589fb1aee960c3d358523282270faaf92e6a420eb3f0f3b699402d6b710c41e292b22ac81f19063f0e9e51051ee07400abf1399819a277122b675d7dfaa88be896072ad212e6136809fb586bd8ebce56ad24b1526dc1be3ecf8567b347757dca0ddc8f46b442ef6695a05e384136f08bc6d1cc11b4a645a9b72a3d414b558c6a36abdc899d83ab50d2a2b5322b4a01c81a40831d56f036d2303f5db2dcb0e47484156e978c49cac5bac65b93df8ffca575b412aed01c8ba826b04f9382d5a81a9eabc90c5be8d52a6d59760f50dedafe0d26b194d7e4fc79ade93d16106852cf166c7730b724c6ac323e60e4d1fa5c6a28db83712aa72a134698ac56692bba233b73f88648252b3150ce4df2b6f0c72727fe289e893c5f5fb4cfe4f24029545cf54e3e4a9ea6b4eaf06371bb98104dcb5447886988e3f71a0ffbfd35129e2b8e657cf0f885b67c653e62fd392ee445511eb2033c94d3a0b2d7dc1e25624b1d0aa9701108e5de1f0fff40cbffa4d99e2d213ade5924c36d0413a2da8d5dcc99bcb69fa6bafda343edeef092f4a0954402de38101e172b5025cc4ddf607cc88a1467a7a2b522c0f27f49ae7e8e8495b23b4aa2575bc08ba11f34f1dee320bcb3cdd0ff378d0859e979b53b5febef528ee5a88d3f0f86fed51aee4165a4a845698c8d5123de72098c165a844eafe465616be5b27781df1742efef89ad070a7cec0869507e89e7b824f43868645d576ac0de16f1bc226f3f941361e3ac8b63c0fbef7fecfa6b8d1defd3917b8b9dfbc0ac6a3d309358827d7de562fbcdd5dcc135ba6799359be4c185af4be35f8851a7c2df60400c4d4b9f1d900e97ca325c39da2e4506d2bda7391f73bd2cdca2b16a931538ff982b663c6c7a9b8d27cf6d302487c7562b3417702d0990d2b5df113bbffd8a695e0c264a88ad4fc5175e9cd6e70e4aa997f5a7326ffd699693ea87a6451be7cd0f86d2d1c0522d99e4334ce08115a12b46bfab41241391e15dba93cca649fdafb03fd2d4a5f7f690ca8b43f166efbda0f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h9e07352b545e38942e666e3e3e091ec114ad2b83cc5cf5bb16dcf1c9dcf82592deb6cc8843ce778058f908f61e8d44953f10406b1d27dfd9d4c9831f0a928a61fa10f8c5bd74333e3bf700b67b8fc23aeb6f1467058c509a153b894408021d8931707d025747bf79ab21bc64ba824600e8f7231f8d75cbaf7c89c97cc55eac29239e72cf1d450b1b07d97a2cf54a659831bcc90a72a500d403e286e3e82bc6a918cb1ad140952d78ec4d8937a1558dc747361a8d96eab731e81691d33a508d1b37eeb72837dbeb110cef5d3c32d6d40f3b0ccf2cce597e92b23be2e26cbe3c44f24703e984cd828e80d4b4756c18672d88d9c166b64abc7af340c058cf92b288f75ef8083f891043815b1a16724dfe9c1b174deba065d5c6287ded5854a53b9a12097559a63fb439fa528159750a1afc9a599541a9b3e7060946125ec2b51fe14f5c3b1d473fabe6106e0f7bc542a702a20982af7c6d9937c7f3508fa303403411cca2d58ccf5df64a7b25c702bbebe02a3edf19292718b070b322fb4f6012b80cd309ce354f6a92ebb0b592a9cc13ce5635576ccf1fdda45e65f273c7a6a220bd2871307fd99fe3b07bc7f9e32b5527fcd97410d61d67ec5eb20d2efef394974a483fafa7d2aff90b6c3d011c69320f81eaa873bd8cf930b34ea246893ea74433bd08bb50fcbc1bca581f6e76b1aadb7e067513a14e3ab08c456ce6253a6f9acde271c6dd378c2ee52ce8081445d39f32fdb4c6e6cb471d95bdf8364c0a9a8a066053efa609df5504f1d036a20f79f0133211d70830d2a785beabf83e0442a873d9212261572af9552cd725eeb85dd6fd52b7a1374fd1bd9da3b09c4520a25dc49d141eae1f7e03ff01ae1fde8764b50a11f26847b5e68e96dd0b4d679af35134efaa36e12d280d08197483af1a38081fcecc06428f007dfba88d6394baff7d72cc28f3c19d3c0b47a9bdca365d56c564a5b0cd63d1c9f2c1d32a185f09e0c3a36172e6176b9b0ff3c166ccdce2e338d898206b90e1e53dc267c2cb1ef5639f3a18d1405e375b10a0b7bdf42eff0c11d144aab0e65e6db0391451040505fcd1b03626b0d5208b49548a0a92c7ce11261d9311ebca38703bb2adbe61832bc51c12fb63f5a7464f66852a9a12a743bd20c12ee48d4201639657b99a3997d3e6e4e8235dadc3a9c57d353b2a9f17983952aa95988226a0bb6c149659f4a666fefc223f7d5bd568297c98296227ab48fd11c5fbacc1678fc4db55f4260d12273bc27bb5ba68b995aab676aed58e89f8caba5767f6489f38b4ddfe6ad06e16ccea54b40966b364fb119f76ef8bc0e3a8488b98e2666dbcd296f03b3ebf508b6fce3aed98c4cacdef7699da0f5ae04c0c38a317c3b2074eff4845473baa73b46941408db02f570c6921c1568d03c87dde1ca39eccc4d954c8015b89fcf3e391b37129c0192cf96ac809c15506aba6212075a7f9cc3d7acc0d256de38162708a4d25199d3ad7fdd2d1667b3e9cded1ced43b73d654d947e7300034489c54cd348e6e81270328b38a7dfb1bb337e2662b286d2b1c518dd5d437d10421774f9e480a1b62857b3fc7300ea76a4a79ff7ffb34c263b46036d7f4fd03806b2bd948df4a6fd70630a23c75b8ad7633497617bda020abb398878d5c211d7469bafd2012ca239a58808f8199129625f03aaee1c2c02a0cb6d351f1eb5de74ef5b5ea2ae8fa2ac818fc3138a0015aafdd3ab73ac15cf7c0225e723966cbd644e3b02bc41511938cd798e431f4f90076ddd64a0c23360ebcd9b57f5e6921a60629baa125eb948e1f1d4eb468fee45bf10e97b699ee39757126fa6fbf398334dbaa517328150b6d16391f05a701e661b9a8c0d5b55b0c6d526238b9d16afd7d618b01e32b79b8041c3d53e0d112a063b50c007b232ce3e949a46518b6303389c05dddc95cf6c7d88719167733418e7a376735bea8e3d123c87523cf791e8a7f23caeb846171fc5eb327b68319f2252397235a59c41a9b5ddfb84decc80dfa787c1420d5c13be5627416860e115ed0eee57c7fd0d4bd9fd754bcee7dff1e1e4e070decddc060aa5c8e5196ad6a613a52e9e4235485879264e1115230b8819233cc4b96f95e6e7ceb5ffe0cdcf431f37e82f71e45b1c776e077cce560185f1b6a2f93eb31b93f4b2df5abff2b4e0e875308bc7f3d26ab2659b4deae5fd48ab197b18a87bf90638276d91da8c87e46c9ef7c08e101e8d43dda5b368eabbdcb1a9c67a10b03bf803afa5c3abf1d8434daa3f51042d04dca82bd7c2fb90c253e0f1964a8a7d51d9b2aed62384c3807382806a5ab4cc55dca23953ecf55bba23c81c6b307d25e4afa47108e27e4a02421db744a09e1a0c61a91831dd567ebbb7378b680fab99dcd111f5dc9ec28b6cf5ed5fa0a0833c85f931c5b874788b24ca9b77fb02cf05e258a55927361f121f22d9659f1542b2ce9690e815b453df3845943f4e2f78b09ab2d821b33818819fbbbfc3b28a36216731ed4312478b5675fe6c1eacdf01d571093af67b3369a7e510f576f75279c75f10a6909d997c4b4dd33c493bc62dbba7803be7301eb40d60ceaa46fb10ca31ce158de745d8974a6357e4fa5a92c7a80669e9bcbea3b21c9b71f8775364d49ee99440d2beaf697cfa49d574af8135d2212b9627c41958ee56dcd29e76bd5e3fb4d899689df9f74b39d55a8b1705b5d3ba53dbf35ad4003bdd86fd110d6ba2286efe1e19b46f9bb98f6583adedc88bb9e885347ddf523fd1e9e5e472b2b00bd30dc87a43ebc7aace82e3531e67a5609ba99a4cd5517043e6a88a73eb563f5af4d1acbfab07a657232567bed0a7bfcb8386d25657fccd945441543e1744d482b93aef5fa0e5bd2d3b58a05e413c009c204410eccb226;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6387de0837f85911c3e8b6b68e689ccd93b551e59e9eaf416d45e8524e104e5a75565744edb7316a94d3da6c9da7f12ed373fa39159aa48f6ca8486f0de1dae1b225b7d88bddebb9762256679ec362679aa4f9f0e4a6cdbb05490faea7c1d67a15c06bbb81b84047dfae8e48374c2d162e70d95333baf7ffd5b4aa3644ef929638de4128d5e45fa0a72f37663c9eba3c38a77181054c2c91699cdf7c70414afb01b6fefc11821d33d4bec8053f17ee505cb34f7e8c4e8dab18aeb0a7eac92c18d643800dac6d1ad8ab718ecb2c21dda188601a392f0c0c65798dfffbab911331724597917d3c7cae9c4ca1ed4aa589c265d93d54b98077c3d27cea1f27e3b1e5a2d755a14fa58b583c33d4d2ab43fd1af50e0ab451d25f187be9f8ed5dfb6d93d54db373b04fbabbf96e265e4db10c97a81b861665618a042a9f17e377f6a221dadda8928bff3054ab1cfe70644f0ab160373a69d5f475fd74ca57e275fe03e311520f2805589b2f09fa2ee9f3be84d5188c32371e8a650d651ca226b0b57bcac1c146de11f6005087e6edf4faecd97dadd714182c2c4413193f05407075a5517adc370f2e0bdada20dde6d97c77c3489b9ef4a9b34de26e635714897c1eb375edce41079762d099fa3e9495508a4f19615731009d8249df7863c8043acc0fd9371fe42a74c6caa31e4b50ac2e937e4efd33967131a5e2821914c2fd8b293b58f59b1e97e959d412454ba9e74dea06c37d4e1f299829c41c525550ecd41d8ee632fd85666156a46b17cb1dc1198ddf3dc96b31687af2fc1f2763f8b14b4ff039ff35744c56ad26a4289976e1c28cb5dd7194d70cfdf3e85eefa7b3d05210451b540a597c7af63296e9807f25a75bcd5fb839b2ed2c604b116100f0bd9eec9751559742652ca9d84b0e87ce2619ccd11a07b965383775f6f0bcae65960ebfcf656687df5f016c8953ddf4b4500fea61057c3a39e086936c211ab10ae5fc4352ea51b8383386831524422db4d1490d02d9bc687bae2e89a3676598a2f96241da6f4b2a0ed75a8a00f7363a5da34106cf4fb4b678c7cc02da911247efda43e8eaf77c36dc6077463069dd051f7e7dd9a38c98d000eabe59fde871b3627862ab1057df4f9505321a6e4403c8af8f9597efd9e53ee769be7ca839bef907f8cf47be38ad94fcde0a1f9ae79620a974fb094e0b5a12eb02e8f6e6b7e5aa7f2351ecf33acfc5528b8f747e40e3c1f292386e91d6f2d89b169749e903c090af7279fd9632cd1dd3fec4d37916db9bf9d2218ca573f6c58088375ff74424186df75d4164af19c1112caffca2773b785b3a48febdf8c7de560cb37c1376ebfe7610486833ae79e069d865db441bc4826ddc2070fc21d791782d27d5f48c2056da55b1a5fd4639389cef8ec8e774dab2099caed515dc73696b76702ca2f43aab7381d0085e81fe6ec2ea9e61919528d3570b3d5123e658c4cbe4c08e44b819a57539ffd01a258af315543ca2d119f227e841c680a127724c5fa5f4393a18f6ae2299864f59441fd5b2ff86503257423a207923105c6aec8c1449649e64e005bb73e02ddcddaf7ed3b180460c10481442a92e77fd26945a66299ff0a2d04df6ab7a9290927bf4c1ee475b00f3dfae788e3e8d608b52e86967356ba3174f4b0921c4d197de9e22b4f0a12b848a7dfef6ff95db7a76f2485a9151bd47be9f8cdcd44e1047ed67793516b201341459480049823748e70f7fbc73d378989fbda82d71556633dae57d94ea96892d4afebd3294766db56e3bb865af37e6cc68506dd2e9449c23db13e56c82cfde28e4a1323274efa7e844318cefaf5e9ebdc30eea94e87ac12d0857db8077d1aa48995e987b9f5b7936ce1b8d3dafa8be753479bff29aa5787d289fde899ce68d053532185f67e5b60b9371bb0d3ea79d7381acc7a23814377df23b92bd68b5dfade30ec98da12fc717ec1b79079a3b424fd5f1caaa71a84555f78df4949a821d39c37eded09c4b134ca277e02a488ff0975e0e0cf5ded4c44c42df17148e9c4851337f8a028e168caadae434bb9dc4a56d77ae4c7ba7922b728c622617dbae33929715f59898b45a44fc5288bf44f342f983aee69b9ba3afc584b6272109c99a42d711388585a3575d7bc6392cf73690f268ca7ded64cf9afcad44700ef04694233174ace9dbd228e8a39b02e8929c366f15e8ff539f9b04c86840758868702f8aee31f85e0c2a137781a714c3532f4a7314b57d1507be35a2a3e4b6f023cc3a2c0f07865f33bbfeca2e1c0e5d6da959b13338aca4aafec45615ac96decd8f49ed70b9fe685a84f0d18997eaf55f419f499b6a86daf75b91a8b14d61bfa42985099395e2546ca06c0db3e4075f7e7d10121200733ca2592de4a73911c5119eafde1f38d79751e490ae07d4e4abc04eb31cdd341f67484ad0d077a05b553bb51597707c6444d54df7f5e7d51d49eb1ce4f07e23bfd375c96ecbff5f93354bb7a66c3bcfce7b7252281b74fd038bc87bb18f7d1a371242e7f07d750b285de36dff7e111279a12947f962e33fb2af2c707e641b0649082b6c0a576e5f7ea3a6d8aa1be5c811f7428d82e5883a3167c3bc0f56b758dc7996c401571fe2cbcc2cd80570b670de0bba4c05c7b8edbd9b83067282f135a8907708a4a76982898cb4e012a8b61dc30b6a0401b4157b9da4fa08a56d91bb4cc8a7fd74a949b82d5f3c15f0e9fd4fe4f7a5118abba356e022a9965d544beefc47a8622b815043b3afed3e43f9fc48e122a85745f65d26bb4b356816667facb1cfac1b74b6f011dfb243180287a050b82e8bca61bf3c1a063dd9f452d424ee9777de8b29b908a98d65aabfeb5ed7fbfad997050f82eb2c5650b8a6d29d09f6b55f568ebc7b4d756;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hec1a46ec6002976aefb2900af10432dc81a53a066ff80d8f044c2fc2542e0bd9bd20500c178aa238ceaf789008ccc097e3d09671123f90c178ef70b9fe4dd67eec6e9a8c185e32dc65988d013bfae6ba25a523ebde46f8afd48db66564e7ea9745dfc98a40bf5190d2c5f2b5a9c2c474fc0e9c07f42e3ea3de45d64677a51c66b2f1cf2af745bff0f4c77767a6c12bfba3ed290b290056c4b02d02515d0488fe153da40bf484ed33e94b5206db4ba6f5b197210eec9503bcb30603677248cdefe1c92e7e0125478bafab635e4a64782d4aeaf9f4f3e6f2fb37b6eb0b8b5f57f5677ec110f9c56b60eb7af455db1e0d14bc37441e996fbaf328515f763bf565c942ef0b33894afc6c61a351aa8a0028755729fa2ff378e799a547a5d8e962bbbea1476a0f450ff99eb7a753cc54f324d406f1c56e65e0039e6b565f9d4fca64b8fc2a5fec1802401d5e7dca0e53e2cbefa94a1a36bea5c1ed72d9894474a4dce0a9f9a1453aaf629a1c1d2a59ef630d1d37084d845c258ba763329a4e879766e062fa3d642f14dcd4baff0426ac5a66c13707838e23dd0c8e721a84d105c7e407bc1dee31621fe93b8bf14fc38ae0f887b31d624732b9fac3a51214f0fef5dd844f46abbe21849bcea922c928fc483a3753eb74ce5e9236daf119600c13715388dd600e9b053bde3b562bc5e2fcbdae5d1913a602a539fa970b6148e3907de20cd9f5658b5318edd4feffb7c78474bc1935ca55d7b634b6c9c4e6edb25efc1cc554d51bad7b8d250187fe16e3b0f682fcc6a08a3a0dcbf8398602f2d4ee42af50f1bde4e28d171f163e1ca9856bb062dc2d159bddcb18e07da81ad7fd3435cbc51152a01945eda095bf6f22c3e266601d00da80fb573289c52e1c6d413d48c1385a01ac82e67c736ed734fc16022abad6bb80aa6793c291cd5a034c804a1f1c799df9012aa9e31d50bc0cd8dbcea50557142b0cb0044e8ca201665ec62bdb0eb6c18fb2d91c23364d94f88892e60b974d130b413931e827a894687b3aa8ad9458bb0f14b166b5c1441f30e20a2972ce0eb6fa2fbf4fcba821e77e8f6c2ab34947967aa5e77d7549f479d6889a35918bfaa985e952fc74608a12d6d04726a74a6da7245f2467baf6ca6f0042538d7f634e9f90d4c8cf2296e2a16d775003bb76a03182374b6cc71675a46bba8bc78e4407388c9711901379adc05f7f680ed64c5ca93cb500e6ff4b0d73956004388742513899fc62c8efb0d84848c278f629104d14c8c6186be3117d2a40d22c29a417e8b6b9546701124ef846ad86d5f7711dea7d381d26ce73b3476f35dbe353ecc6066121d2196dcf4dce7166800137c3564570918b0cf77d039d7923e352db71d0e74b8330a777416d68e536fc32a350ce1a2d483b48b99b2faae59cbf998c9bad7160cf149a23c72bfb79b0194944f2bc39a162d7334f65499e4b2f4998c69843729ef30443a492f72e9057ce8fc72f57943a7b01f1d6ce8a32842d648dce276705af9fc8703aa8335d0febdf75f743fed8548de89e058158e8be3433b9403dd7cd802159cd3f8c76a690ee47944db2e44eba55d7ac49a7cfa08e95509745dc66645a3980f93e9a19935006a4d35b9b062545e9f705e8ce78aff8f5fb6528147fa65e5a184e9a3a7e27663e5cde6893a1a3f08f38e9d85c9afbd707c46101f810f54346cddb48eba7f60d14155f40a248fbe15bbb01fc24836ec6118e8b3a977e19cd1a9bc255d6a83678bb31dd834dfe7f5195af4f6a99fa6bd827449314d45dbee87b1fa828c67d398bdac42531cec9c78b6ec3a9e946f1eb4f9abe5e2694d63d4e9e081063422d7dc2dc296a3ec04f11a12c2eb4ed6983a80ebff174149b8122232d854d2957a8e8252533da627071cf396020825ae8feb33cd96b602f676c0c0d5d8cf37c2a37aff68b4b0ff7739351c38264b62b4cfcf923d1f8346731dae834116f6708fab9ac78d3824373b0f0cc0364da37073295086dbd8d48ab69b6cb2d3842d8d2612a946807386e818d2de131e5785c056760bc43b5fbbc7b5b2295dd49b9f0d7df82fee23e0a2114997b8d5dd4244d0175dc34341aa9f19a2b0c276a109aca8330a6e57054f0dcf13768fc91987978f4e1bf6d1d8e1f061385233f9e06300175f5de5a646907af4b4f3af1af0cf14ec3e816e58e5d1385ddf7640fe6c88e8cdfdc0f84451f78856b6a201a3f9a7afea0b7ef9f7c36851d18e366b1bb3953597005a521f137baf418e31a2373a1dc4b3a8ec08d3238e564b0ced27084170eb7c303ba5542a86ad94a22efbfb562ba95d8d75dac913cfe49d849f95d511c7630bba88e459f55f621528cd661d8a13ddddb29f34821da49274bf04dcceb658a8d33ce95afeab798d85f725537669c05da82cc04220665c281fd305ed9f6a7f888ccce9cb4ff726fe223b2fe5f74e75e6dfdc0310f59b0d7b0b4fd0715fed5be6901c32bcf01fab58b024cc33156f0bf40abcf336750b1afc01a5492e5b800995f61c57c94401647999afedfdea831b29e959d7a3a79dc681e9c516bb0ce2799010f7530c6ad00e81b50910bfe1e51b3f2d76570c14930b032047c491ba05f266b1846eeeb0dca372b6cb4fb99d06da11b9802110de2fde0db13c4f7c618ef3bf4b66ee43154f7b20322c65c863faf7b75149c44ba8560eec159b0cdfbe754c330e775a068e338c58eb736c81c5983c31edd67fe2e7788a6464c14f908f4f36a8fb58c8a6ee50b915c9544a1fd03c4d16fe09fb41939eb30a1ca82f8e55660586a448fe4a235b824a75e66359685395cfbfc683cf821a4001f9c75b6062bf361ee19105990e742d938cff35972c19095e1bd2530df1a8e3ed87513eecb8a05fd5bb9b1a84673ab9d2ad54253c2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hff307e33793730d3d8c9f94349ee1e4572cffb25333b5ae31b20dfd42cc83c11bf353b1c4fbd1c8830acfe30e16a156a1292cba2b7f9510f3af25463100d45fc90a6ab5aa58fccefb5de4159378902cb232ef4a7ded259a371664b8c0ba71d7b78c4050917f948a2ba43d80814820cf46ea2d36f51687f02e343d6eb8b7c27877c56b73b451b792a79db53b8607b371e11f4b679cc395b838c227e0dbc3d88f74d5b592b6e6deb291ac590f56bf537f5bee3d223b1dcb9b31a8338c9a3f56336bf92f6b9c0dfaa8b3bb2e1c418f99771a0c1026a3a2d32e304144f0f4dfc6054ee9427749a417170d3276ba733805995c820261e881d354bebdfa3b31a84fec7489f95078ce846f7feb8834055c2adc6c3eb68fca1e47155b44302d26f62ce920cc441e38ebd171ee54bc761e9ed63234d8da815f5ed9f066e86560d0a66acc16fe1011e12452a0a3688e1e88bca9431ec42e4ff2bbec65efc2565e14c1ae977945cb30781b9b4d734ab5b1930645bcd17802c82310f328b4b35578980ed1a3dbe4b86ac9d6b6300ae2b5cf5caaaf1a2d6ac656709552e49e99a7640f643be1190252f25d394c001e73455a60cb07bdf5b0e5c032fd0b7b6575b46f95c8c185c17ecb4ebbfb0d814b948fd37c9addb62fb9302af606e8d7d0ed1fae71dcf70c4a565100b50c6453e8c4c74111f2d8799cbd398e9bba6e830e07e6b916865d9628b620c3c725485b452850288672f1b132b9d5462bb7ac4705dd254ed0dd8197eff728a825f1933e58ba56125467831e5dbbb5adf2ff6df6e9a285121edc2b867a2303561175b467d014947e18885d2e0ab9678324716e17eb3db6813fc8bc8e7786898e6b0e476b0e004005849d6a71fbb2b5551b7bbc895a5a2e073f49703cb22b79a22b0960c4dc2471f7de6d0c54f603a650bda1155e7d6d996ecc41121e4924d95ebf3a212b0a73e3664d6dc7d58422abda9dd52eed493fb15a093b48fbf720a76a209f590f84ecb00625cc3eb4eb1e375402571a1ab2cc55d7e947ca7aa94addb43c1b1ab4d8b49809ec321a6b3f971ec691d379076c0ef92a0de72451ae0431a0add87dd4098e0b4f679ca833ee29ec8b8f5bfd8c99081b814772c328d13ed1aff8348e0515044dfc034f491d92812680c041d1618c5f784e5ab3dbd4e2bf15dd663f905809c1018c9b960dbe9e8003b069b04767b5d330af2678e54c6ecce0720cf7ae5cbddd262c88e15e832f724945e897d8c7a849a078df59a7bcae69a6cfecfab1f0d6d874e5b160e37a6ca61c15ad4064acee9653670d0e6fa1f390e33bc02dfb1f8e244428da5745660508730a5797ea0651a58b95c663726bfe4c3d1f8769286d82d8df730efc7e8162cd529702641b1c51bece49247ff35afaac34b253c307dcbc001e6790d6d76e683c93493e980bafd9f3ecb6ae94779514d913f1c794dc92193e4798dc7e2a57cf8aa2c267e816a2162269d604592f0e19c60aac47023780818edc45e831f9dce06e8f725c3d5c5d7ab52a6ab14da3a21e8d377fbeff881f80ade2738d5623baf5209f18b234fef33b5f1850b9a92e99a0700a0cf8d9d2eee3fa84b1f6a987e3ea4b1c433334100dda0667bb18abdec1c87a54513533465d43a2dfc759dd38adbfd121de0b63ca9f5c3d5b4e85f13a55d7ebd556d563ac471a87f4b75c5ea54b81e95d0ed0295aa66ed3a436b1ccb6a6e513f15d2636374344e4d34e26b0d82f56ce4cc97660989b49bdfe669a2ff70ae9cb4d81a271c0b3f025790ef06fbc15785dcb065a3005cc5849d9d287be98ad8f634870d3dcc7aa10c9c2334f5208e7a8d6fcda65a3014a6004214bad88a3e2ff3ac864c6b2583bf246fb947a5522d4e6b4d9183dad964ba6223f5a2d8690fa3d59ae6559f269cc44bac116c86273565c958d7c428cb250b5dff3af44623b9d43c0101af0b20c276dde94a936e5eb4fac9a42bb4fbd870c0cd47b2e7ea38790430d26b9acbc8b01470a8ac06ee7f4f579a0a5f398fedb64648d39f4d956d149a9fa6129a425526a6e954b4018f9b5c8e9bf0403838da843edb9b32324dbfd4e8e4441f69efedc2443e7688c64266b2ef720ebda3cb85a76e1be3bf93b0cfa78dd8e01fa0e7d8646506af4ca2551a973e3d2906653b751dba8a3b886420c365a12c9eb0531fb87afea63381103199716e101850a37b8957d9863211b307b0aabaabd00fbfcf6da86aebdc67f51c5c1b31ed8b262befa561d7270a2ac0be3477b710f882f7cc0521ed36fb55ff7542ced078d014102b52d7fb7801e630993a1c939c03fde655c9e598254c7abbe4a944e334acdf401361c1381483296405e596d5e634737a06b68d331f96de85228525368ebf246ed0b8128b43a3ea576fe555a1dcc69280ad97c213d5a2e106e6c939c6eb7ae942ef7bb05342a16d6a327a26121d053cdb1f374d0e6b512398045fe4dd8c9b318244c4d78cc6921801355b368ce9486124700c94ef8119ebbce6875c1cb8bd056397296ec94368eeddf2a7789301916d43275f883f132b4b3156f90c26a34a91150ddea0e94fc7a0d92ecf8a934a975e89754f6ae149c7140c49fa9d9771ed7b32db507363403dc9ee9367c83d3cd7199da88fc951730bcff0b9cae008eee70b9c8feb5e170c507ed8e7e52c269a5ca1c3ac178827bccc85656286048a8e84b72791f26157c2f879f8103d9186ff68c4efce57e5a83e18f7421ce0cede43eca5557d95c2c4f4edaa82306251af11a838b41e4fd3ddb9a571f13550e6ac4b04d0d9d8e94a19275240b702b4c34082f5e6b9ed7e09a98d499416dfc0f825929d0230e2dca4776dcb234a34f4a1f45cf7d0adc1675b789bbd1c61876544b7430de5639bf91c87e19006ece49b4878;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3d838f9a278239e3b147fb852efa18173023b81469dffc91ea2f7f9fb36e7da871272fbf3863883265860a3a33ec125d235c3da65aafff23c1b5b5b6398075cf1b7605721a8a2a137e0b05bb3ce30b8a6db0d4e0ce22cac5e70bc99cf45be36c723ed97db8d04dd226f792521af451e6879f2f3f0e5b745482c757d90e0de7f8c9a131649e2820547c57fca2b1a12239a594ca9e5ccee5245f3f79b2af657b265b2f1af80c2543b27551e60cd331b5a6752ad3d8f4d6316b27291039ad8e798d2d7eebebbb3c59840bfb0a74ec11a27edd20174f336b8dcfb431c190e7d50f12fc3d2e3d0114a0da469505c6a0a74157fdcff667d3919723b3daeb4d2890b256733837baa26b6ccf7ae9c8002d320ec4cdb113fd01933491fba02e23c2afe2e5d676137e2dd0890c5f0f5fac6fedb5e43a25649a50f008cdebf7535870247f83d8723b000958acb94f6f4acf705a09dea4ad06822f9cc70f795b2c28be53629838330f757329122c817fe376d70d24eb8619fcc49717045184f3de37f8c44e7e7ba8a843ef1f20e446ed027a6a83f6f92439d9042083f56ef9706e73166959ae8ca728c47705f5076a2d415e9f40a128e54d2170f43824fe0a34f91d7950c0461ebf98a61c1bb867b2f81cbc92536f9cb464a8ab4cf2ed9438a88fe77300c9e792619f90b92167e1450460e563f7f55e9797c274890978c2fb00fa46fc6997d5d1be3a569a70aa17210db799cd5705227b5b07385b7a17384b9ee1bbbf916b5285d0536ca863747eabb482a39904aa8e78c778cabcb394926828943de78b6690b3ab8c5e8d8e00205fef7ac574b6da1a4213845e312663ede67e05565c5bef1b43d51a67b899912c8a6c228f2d7c756d459dced784e261bbc75761ad1a750642c9d694242ea5b766ae2e6d872a99cb82c166e9daee01dd4c7b7b6784a2de6e4f6e6e93f2c0df2089d796e0eaa886cf654d2cafbc914d0b77a00abf6b8cb55c80941ab7c15732183360ec184b1b5e61477e83ebee438eef8e078a6f83ea40f5d9df6dada7d6fd4919cdc8acb5d8c565b8c0cfc26c476e9e34ca5fc9630e37e0567709227c41786f85d3c04dccb8b9a46d058b7f780a0f7f82856c9354a668106789acc20935e4cacc8b3384cb484f91c9e7a56b349103f213e17861bdd13369976b1e81f08e4299fd293730635bda6f86ffa37819a35b0ad4bb39277ef62198d05bdd50fbe44ab9c65caf09353889390c3982c81aa8469b7c48200108a6d13c00341f5a77c1a6458734dd449df5e77dd4629b52dabf0a31d7ecb1fa30c6ae9545322b7ea8153ceebe8627b68029b664bb75eeb8030372dbae394e59b27abd95969c5d1a36c07490c1aec727321ba84d0206d4b079869ec0a54f6ce6f0fe75860c5b968f8d8869a90fcbba650a15fc7048ae3e456dd6347404c3bf082c10f30f4bba3b75b17094f11576b54216afc55be89e3404182ffb6ab675632f55a9dbf3dd5f9c0dd0c7096314c63a15eca0e44a71d6f1dfa5467094ba9c798b70403ef6f15e4accb0aadd1f00fb203712cd49d3ab5084c59dc861f21536da9cf8252f12f31255e73d79afad3582020a5fdca2767e81bbe5c8450854d4e56f8640a7257281a184b6117f35e6270b2c6330379f3ef5f340ace5a0e116db50560cd6c060ed61ed05ec0b41cfe02455580ea3ca558e911e7c1cb478fc642d6e0f104c96375af1848b1f671562a8a7e6dc2829ce5e3e4fbc88990e1e1d1e57c033f894638c4fadebdae9b86c6ea1e3d7d236e2c9c3255a106b9996588a5b09fe669b79d42dd9e17be19d574d6add55620053c931cf0416cf89a34188d207a9e73806a8e28573447cb801b16d310a606318956610c1ec827449ba06fc0b8b57be50e7267c0140fd2dfa6fdcb57e128d9f42d2d9411a94da59e876047e2951245efa064cb4734eb376fb060debd8325a40677e508b5ee2c253a933d052fbf36cd261705caba2f5770e23de9fb46d8f969d38dc1c425fe482f932b4977d71b1aba226db09bff3fcfb2bd76e6988e57107031978534806296da08f2524baffa632416db43739746a9378af874277dc21b044460b6d0a300863a2223f0207b633a61bf3a3bbe1fedf1f104600f79fa21327492310c58c463337b6c1a33850dcf28409fdce4d80c227f26cd7e572e5e1c2c6ac784c997a17166265880aaf62b4a986040e9ca4547f4ad20957fe22d3c80a2546f1dcb45f7ea30407f6ee1547f020fda7f5df74dccdb4fe17b2e9cd883d2629fb9133467089cf31aaad198499c57db5345fe302994fc3abe3ac5891992da531fb32af382cb2761ea0f8899438f4041b1a0560378ebfec8c537bd950bf256f9921a0fb5b1a172c69ab8ab6978bfa9e4c2134d83111b9958c8171498f875f918f9501d9261486208cd88aac96bf0e9b9f3b62653746fd42963179f7706a6d9a38e42daadb24236df81b41ab65cc3f7461f2580b8f4a2eb4fab3af1bf02e19e8081c79abd31e0c635ace949637c1adafafddeb4426c78feffe17bc674681a8a2c2343b65f505633d7481bc851d106b9da011cf7818702416761e3f7fa53459da4312c28ecb373ea9e84a15ed1334dbc1e193fcd2bfed207884bf710f115e24cc8f840e80a1db23a6b2ec970ff50d4f558776152e9ef1a9dcb0650172269000747fe311d382b9d6d8a85d6081a4992ac29e6b8ad80cc4bb0de6ddfc440b5e6e2d3ada3478fe71d42569b19263572e0c8e4de56cf85d7ff30b0425b2f1d665c433ec3a505c3898004d0b062e2e4b3aeb8f5da07e205e622c3456a359f0cc62b6599420d51eb80f8d3534850ae67d7757c1fc03144ffd990206b29228cf4a3cefbd67aaa5f94c20060b3fa3874edda6b261161f12c70ad00f9fa4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'haa7f14277c538f9e978e1c42a7d0acbfbcc2252ef86331683fd22dd00d4df3afd27ffc61832ecd3f7affc3ec39024801d3dce068059bc22589b91067c37f0a40f455d2332a64c48986719777cced9bd93109faee243d5ec2de3d3a4b68791dec79907871ab15f24d714e699a8593578801bc3f83b979d823575120cf19061f38bfa1e44a8a3cb40cd2bfeabfa1ef095f6d6fdad623a8833a45815ecca4b7056387d0a478ab58182598876d323efbcd3e811424acda67c8a26d801a6cddcbee5f71192f89cb3b9366988ea3bad0a816786104b1f4811bb30a7d36c1a07687b581abaff0fd149993d4b55d3e62bd72b3d50c0484f92ad881cbe1d806528cc6b6ddf769e0e6c5233fa766c53e0607772eca70996115602db9427fbbc6587624349d067de60385c819d5e4d3297904f5e94a0d03744a008c1c8ffdc792d26910e3160ebe9555d1f98017e10140857b2858724dc7541b9f8e4f35d41dd0aa57aa186395b29ee21fc1a417c195e71e684a389c501a1a4bf9ea37e36e9419953fd27dfe9947efd37cd31eb98aeba35b263050d7724337f483c091e41fd01f99eb2c1c0e71aeb7056e2009045ad8f95314d7f39e872b30818c84c66a08094c487580d707ff63d5a8e6f3608cf41b13900087c51968f632746d7650c748dde62a27d3be2770074bf9f0df74c7e28c2b800fb4c303a8af5457e85901d6080e557d034c184382266c02219065832b45427aef75a11d4449f2903ddea6c6dbe7157ee7605427def9c516ff1f9822b2d3d2ff20a8480634cfea86911e896d10b45b3f65459a2f4d56fb0ddd7f297af7422385ad6a5dc311b553daaff9f6ed5deefa2b455ab9f60c1fc61682a8bb2243fe09832d538a65075447195b1702826adff72db09fc7f923bce479cf472a1ad8b4257ab7760cd8a113c8557de63130c50254d37df2b308a45f34069003c46356bcb7fe0db5b3f5b437e532c8214d334dce945ee81578bb572ff81d56866a1d25ac50ec7c39bbaf415bc783b4c668d8213ee061040f41a2e109a86ce94bf96564da349d4074adf76a3683f912b11d99e7c4540b861e2b6da3b92ac5fbb782dff52d3bae602e1bb09839faadfe094a723c7ee8b223d0fa2f06ff7d3a2a93beaf6adefdb9994ec4678fd1da343eee4fb52cbb2fc74604a4f36e8ce0964a6dd7bf9373cda603f9fec1725c4317367d7f41c81fab7f03830e1a5f64fd29743bfcc870301abd1f046338ffb80c264f4e19188461fdbc73c8c31118bca238c285a48aa3a847933ee65d4f23e83fc8baafd7afbcbdf8c4c84c07d80306eff62305f12a057ae046c2c31e8a61b8583e716165aea6581e7cf6421b27a5511b33b1b44fadac72ab325cbe72e41099c59edaa9927a6df16d71fe8cb670fef98f394768952732fc209d8fbac42a23ee0ec589f18242ea2a85b970a8248caf55c15e06cbc83776839a5ee08bd0784e937e123805125df9b8d3e27f3d17ec8c553c37323f13cd7e43136c7605557fbea9879270965cddf1e71fc71616200f9684b9670e0b8a80c8f4654ca7e731710fa8e24c728600d31f1e0c8d9a2b4cea41a55d023d72020210b6af448796363cd883641ca8a2c1c337a909317d881117b74806bf9bb49ba2687ee786e1df62590124b5dd9d1137dba475bab9b6509a52cea65a685f2c67b8dcc2ebbf92ff8d83aa543b5f535e920ea553f74e9b05c63526cad929e52ae523114b423f4333dfaf75e64ca7a75f0ad96aa9daea2ec96fce3505453c7171347e4c8c3636a37a8548d37133d331e0e22e4fbf3ab794c6212e7641576410fbeec8b4ee0197ab36182b49481df9d1e911d886eaf7e29a3157575bf562944013cffe4f78eb61bfe2e91fc89f8fb4bb56a6ec504fd8f932c486ea6a2d3664783b9713458a72bfc76f40b833fb0071d7ec37875d740dee5c64c39a0f9bc46fd0623e802d1d27c12340962ad87814363309d832765c9a32656f6febe5f860c3d7f1642a3b141d32961b6297087bed96eb98e0bf4b967c3524cdc3bdfaa6343f1dcb68f7eac3145c38bdf9f62fd6242c67d8aec4b77cb16825ec3cd1d037f9207cdb4c14071787cff0666d8a2cce7892b9b1700f1c0366f0871ab9636436d674f41ff2757fa46a3079cb291c5887ac6c86bd266bf31de4993d669f42b5cdb6d30d6b9deae20335169c775599c67f9dc1bd9287d4d3bc69038900630f1a70a9e780038c4aabbb6226eb04299f46f67eceaf89bff473c75a4b3e6507f588e4da0cd6c7703f6a3ebc94bce69906a06bcf31957409e6b51b3ed32aeaa26c3639a30d3942650a1679e2695998d6758af58870b8388edff6a632f1554c0d7b81822215a3585947ac18b4e2597ca6284a643e39240714ca067c3354bd4c1157e1bd6eacdcf729db37c4ebd0f279a177bb9321bd0a846ad81a6f7519610996849b704b3b47604d02df22697d6d50df73b8b74c2759ac994f0b4ed13140e02edfa60ab77f328a792ac2b5dcb574707812ac62a5359064b1c6c99b1eabc79e74738b660c4591a4bdb33ae4ed6a14b84dcd6e7f1df10a6303d43c9bf29043cd8aedb1c65db74ece27d9be03bcc3803d12e242cc39574d560113ce4910f869c5325f87e8262286ec3ece5537b8447c6160d90331e635af5151a4ec83d942b75a9b4261477e549cf2a9a82e4ec55538385ce0d88327fea8ca4f4e79acfa2c3bbce071325a93ae4a3cf761c2a39cfa8c988c1cdb86d2ec8cafa26c012422a933f9e5bf2992c8fe34ed5ea96f6f96aad860ada0fff15d1538dddc6e4a1e2c15598b5a2e27e4d71b4ec6494c2282fe813fe52e1a576f2d7622a4d4005ff9722e4b211ae582f80b2e0f6b6114b76ad81df25dc5f330e2b18674c66ba851d234d87ac03d3c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hebed378c005d5ab211f50307ee49347c4d58b60ace2b0e968ed1c7ed201eaf80a716d2505c84036dec93f785886b5f7d9979b8240428c0114f4f880942d56edbfbf6b509c02c8eb7fd94aa8aa3a087c1d2d59d55761d225395473b0137d2272eb0217f2f8dba821d540e0b9a3ddb047c8feba794d5ed60fc238a71084507e1be750c6311eddb98e2ba3c83e442075067a7e84d2f0bbc67667f0ffc186308ce4a521d0562e2210a2e86ad219a6ad95feed9bc985be45d86d7a48a71e68cf5468459df45055856a9096016a35eeb8e7a40b7e5b18a427b69f7389097dddff172c42d58899a575b65c8dbc07a7bb32391f8f90fd163dad8a9cfec15eaa7165e58c731b7ea8c725ec5a1829325ecaf462aa40cc04c13b0c3e7f9739885e6b759547c0c1f09b70df8e215f2ad5623e2649fc27cfbcb13d3c4f7c3d4625d1da98dd42689214370e9df3cb4fba1207de5a5b3b51bd44f238e74c7a5b6e7768f5dad8097f957444d79b0c8c355fc25b028d81df4ff79466f1fe5a9fb804dae7df49d6757e51cf70793569a139f17508239cb44a0707d5d0ad1e4698dac7b75a43d5a0027a3231c8b704c81a73516ee17e94fe6a9bdef4baddfc9ce38582e1a77f9d26563593baf746b3903727082ff7aa5638b2c3164d5b8c649a5071cdcd1613c75a94dd1e6dbcd146fc87b2395076402e4144217402710b3998cb0c416b7ad2f19152b558f70ecb5c189d079d77832c194ac6cea313fcd0cc598e8c012ffac73feca960e043268332be7a389501272b3b31847d9a22667abea133e1214cb24c74e7df378a59b986f1adc588be714a1aab1b2af70fbb0c57684030766adb1d7d212e42ac62fe29de2cef9e3790b5fccc05a8f81a3909a32437f330845142724891c42ae2f1a76b325c230087c305b520fc26cc00f89f5cbefd66bf5e25eaf709ce455038202c5403fe2c7a1b5059ce1172c5a82d152aad5282442656b020b20d50cfff8f185d139a8b5e27ec0dc5bf1ca383aa06204d5ff5c23bd24ef1ebe296b1c6c01ac5681841714ca650dad12ccfc2f61a0da9a6e730a31c61bb4d85bad14332dfbe1120a1fd23c1965628ecb95afa68f146c4dd6fadeb55ee53a840aeab6e1ec23cf606b01b50fbf80ac4de906c74f001c065ec56ffc4451f020bf49726ba1df1538fd373bf61a10831988cece47e750be92317ac0812ccd170834a03e1c728cd4912f7e65bd057ba271c944274444355ac2a21dd0d2d1cdcecc047bad11220f6533eee6905fbd1ae34f0557ed8f244c52e5fe3f292bfae4bcfaa6d1dfaaa23d3ffed4ac3595a7301d5fdc2474c955168e153e4b6304a3cf3c943d1559f1f8161cb72c606e3010e0a9a9546c920324fd02b9236df583e246db6a840ff21005017475220ab5cd2bbc5b87b313aecea465c44a75d8d1a072e7d177dd9c4feef7a57f54a069b97cef0d02def50c1e379fcdf5dd8bdd801f29ca8d00b433d07f419426f822b1c454a810eaed0db2cb5c542458b381b75f0f9150549f974f7905c4fefb464002883b09446014380e1d2fe11f8e25de3604f987d6f1e3c7a477c875074ce05930bd482a8af24e0fa4966525ed8cbc0d142705ee7271d35d945fa9f2757d7a89a8dee7e12185c808bc0fa3e1e4cf7ca69f898dc3a553afa2784304faf65712d7156c533fe62c2915dc12fbe49c97ca4f7be80548aa4df42c160b667493a5a8331a02b14980a4c7c22e6f3532f340f32a07fcd1ba5667ac0fa60f786bcdfe0887ab04833e4821bc1aab4ba16ebd9c439b7ead0a308d414cf62b735e788961a2682fcb8e30f44b97ac8b55a6e96dce97389d31947e4282075b35df1d3aee66a6e873d81be0c2cb34098e9c901555b3ad7b0d173435726e0f0c8b1351d37fba9477f2eb685daac695976bd7f4979604298724ec8f3e62177ace8b5b56be87b242d790dbcff367fa6306d65a61e844fb6abe48a31ef9126408ab67ad42d6d3b00a3e3944acde99b71a590c4961db1e8c38926156ff26f97d46f1191c557e8cc04062e9e455c5834cf021d94037fda6500abc2ca604fa3dd2e19586b9989e28b97421f367ebb12e9ba4446de7a04e9efbcc3dc142011fc39a5e4f2a128cf0e4f128a82168280379273d8891abd4f0f1ec5d0a7ac3cb63b4478f10963b2a99d647351ab76e2ef13088c76c98073f1c8eed6cae855fed2100f595b21b1484f780ec4100394d735c472a95f690b75cd0729899fa965e2e9d6472b75a21b07eb3acd9d743221050d6a1cb9d181581f73d463a9d6ed57255fcc70624992e6f69aded992b1f047c2806656cb4f1d6751f750d9eaa6dcf58b0db8c78f862b10362202fdab8e973334b821c1e0b8fa871b745f407202c3dd2dca85dd8c391c26dad617cc744c6e7083c9a5602e518fd93240ca1fadfe9df4e6fc0409be4b59473f39a5a9d7eb9974db8568d0f302eab5dc03b1cef2eac01618510a4dba2ca7447bb6a9a89fbd12612ccfade1898fe57a6e371c8975161ac965c33cd2d0e83b496bd4973b56d664dd92c120ce8e3a08ed0fc94def22736a06515e71babd786fbb4e6865b596f8535d2a1b8409f61c6c691d608a79bd6529f28ff89afe5dd45e78f5dc3ee9fe5c251d05b9eeaec5aef3fe8d794a79b1b037d352b972dbc14b1258c9fc43077c2f4441faaa47d77ffef63e292473004f691a33b6c1f098e7bfabe11c33081bf1a3866efc790f3f05be84a688b591ddcc46951764545a52415bdf1251ee02edf68796e1957fc82dbbedb33b1ec18ad7b3e319a17e2b0aad8a23275b1ec6fce083e224b46f06fb8e1033cd8eeda2e0975b54e0b3c965b5e1c925506f22320d4f0a81d5ad5d51f6a6e0b224fc126a456f44b7c0e09c9de7b56df51d0fde372979c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7aa029d7a4643b483234dd0f6cef459c403d235f3ee751907458a3f1201430d98d8d55179377a29e9a35416f6694912f73810eccdc8d0e66a6a9c618984706427a56545be46df7325e333f7c65cd82a308bbc7c84827570d93b06942be8ef329e3ccff909112037bf06414da98fca663cf0335ac5e4da494c96f0a25dd6ff8f79fd23d53afd1a6a0b8840033652f5d3b6644a06f9de1479f48cc23466d202a3a1f9817483a820b30a5455b12a84524660187b529bcf58e5db6a8018d9f6570d74b033620cf27770b6f7fc0a64d2810f1337011fe6dcd969aeba1d8b7cf2a9eda3b2275bb19fdecee0def1c0468e7173290b62cf2250f4e6ee21109d9f9df88b4f3338316c77b61f0b443c8812d3d716712c4d4ab3c982df4d584f4407fa2d6195661744b83fa3c23f70f720d0a8ff1efc4885a638ebe3298ea9136c71779503874a4f2c66d37a826a16ab6064e7f6061243a859fbd8087c36fbd951783f3c223ad2929ba0ba87d6e451644e33c2fa4eb5fedf0196c4ffc70cf3af7e0177147c1c5a194025a384cc0085552668aa7716b1b2b7e35004de27b880c62dd9c861f48982a0e49f0ea2d96dbfeea7d9e51fef9ae991dc9bbc0215595194da31de03076f475e69d686eb828e06cc0b47313b0131e52b23c38dfb6922ff6ad1a1494367d809ebd5d1f5f1a47988beab789c8be3ecf655a2d682d9148d0ef6b26306dbd628db53bcabd108ed5d7cca23df032a910f77409f98405ddfc73db3d708fd0fed976edfe8f4d040ef2dea0c510df92ead24e6115febcce6a67f4d7b2ffd4fd9776267b257071d4b26b7db2b8d40a0ea1b88b37c609c1690eb94163725137fb78efcfd20e93d80cafd5f5b1f2cde1bbdf8aadb7655520b25453b108ad8f8369b7f0276b3b9d3cf8dfd84d09e689b1b3bf099656d164584f1f40c8d8efa9e257d5ab0f63074c381baa5663c1959cf0e61bdde7eed25d458182cc2beaaef540db9b4907e1033c28c9ae280fe6e24e2c06b2e73af6a5140c2ac9a12e4f6f2a95fa291189d7ef80c6dbbf10dd476f79815e6240479d0423ee69840b86b1dc9c402568c1b61f88843502e8fc90c17d2277db2b15d937903489c243bf0c53450f0a2029f3388ba62ac628a29d5f3659d2c526ee3077dc1ab0919f1a2b0b42e37b90623bf0bba6b0b9d1888520fe4ca694f88fdbcd88feed7fb23f369a61f5fdcac282735f7fbba5bb62fb17f2ebbfaefe2f7bf932eeae69e1398a4cba9d26aa9b17086405f9a3d627a259c3c215d9e7bb63afe1e307dd8ea44cd087e2294cb52acb80249dc26477c310f88e693baa2c757601c016e4fead1df4d695444419273ce8f63ad82d0cf1f22d31c59e85eec483b452d9c7d355b983da05ed76f1355dcdf1917b61ebdf11b7302f660c95e2605ea547e1e622457cda434e78a4b1cb21daad7de9e99a7c070d18f8c2ced3be43e80e5de3e948e4b17d75dabdfcc9f8a50849a4f1f24bcb9ed4367ff657c2112725d17e388628dd9b3971afc2234e01fc16a074895b3717b6ae0da296eda5a86f061206d6588b994e1049758adead4f6854563d3f0287b2d79d0ddae73401ce502adb5b8adfe744339452f1dc6ac72fb9e50db36e2a179b1d2f8d325d1188417cac409d0a44543cf9f58520b33c2709a3037a5e5fa7a758d3daa36e078ce18ff8cde7a0b605898ae1156fa2052e630fe45f3137a61f4dc4709ab6f4cdbdd03486604f2b16e1c85edd8eaaa04c50121b190da48081aafad6d928a081186ca324fbfb46acf4f71d1b0986be98422cfb604c99cce610911196ff6856998ff4fb6153f513eca13686f5c44da828a7fb9e39038e93ec1152ca7f0194e19813d713b8ca606bd39a27a8d6db343e25a2d50da368b4a7e553b509ba2f2eee51cc84d2f6a38e5554c3830264ce7c42e670aa0159be4eafc1354eaaa434483a5b6b93869b755f77a57fe13aeb5d2140f9f56b689651d3f37cd9637474c5bab174881f5b1490ff04e69435d0a69809d6fe18aa1cbe386c4030c3c25c5210850affcfa700e9c6c6946c6d0fd68402a11f9ca3e1d8b148d24f709c1bb90aac299cd65cd97c578bfafb81bed272ea980c644351e9a0ed2e5c082733dccb52e8beea6c9563c704d3b379a567b0746ce9ff7133e50bcb40729dec2bd1f6f8890abb6018cc9ddc12b0bfe7079ac83fcf151961ba7560295514e1fd1caaff2f6d407a14766eb25012297286cc1faded3d71f7538715184c6d448311cb84573002748e6178bd8a5463322be05fca97a52d17d8f3871b68fb7ee30e18c9cbdd6222ccb1391bd7e6c1e3d7c6bbf6821de30eb591421f414aef199860f4e5235f7f6d3db472c7ecb500619dd61c9c22ed97168965cf11f35192bf2cfede39dbf8b37fe65f6296dbec47e2fe8e33b8f629c09433c031c6ffbc055ad3d818ffa757d67ec5b9f845585fd3eee8fc8e16b07272f3ff419364ca3651cecbbe587fa380d1c9441484b9506fca9fd29fa18628702e4bed033391ad4466efa58ebb680d96607a5ad4dc0b19b4bd5089e2263391ab44cceb49a0275cbfaa1acaef4df817f4dc291e0c5ab3ea9a5a2c8153119371ca078532b17ab730ccadbe8833e83c18e915108335a1d73649ccfecdb783a0295aa9f3e46c0b847f756ba5977a9216397ca51c4d4d623dc77f7510c152b1027e193d5f6c5f7dcb8ee3d990188deb6dec3471f3e81cbb87140d93241440ffa1f414c148d66dbbcd97030b47801d03abbc55676dda258550ab0d25b65e58c84e60b5b78131c70f90842d4721180b14841e42c5dbb956b5a961357c9fada7c7d28da0e96b8ca68f18e5f73a710cdf37a795b8b29bbc30a928ee3e641d365d317a2c5a16b2b00fcd5d16c89fc2eb478f6703f9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hebff0440d2a11f5f5fa18d5b18d5e7cfd64784bc966f0bbffcb4b6a6984a9c83d6483cbf32dc39e4d4d74447464bfaa9ec535bbc130a22049d266186c9363c7465cb2112dc8ac8fd1bd7656c1fc503fe320c84bf89e9545c88cfdc03fbc977c8c684e000cafb18b5c23dd91480c71a0907b6ba603cd0e6ca00de591d7acf64d4bd3f84ba3f01ff6ffe5a6cfb60af1a1d88cd146abce1fa9ff9f866c34eef22b9423c9a4f1485f78aa60ae8db5ea456e97c16438ea67edf3e5d5aff606da9ca4c14f284e2684e89d4253dd783b980bb57824fd40376a932726da520cc339580bb0daebb8844ce50e1e9cd3c5757b96de53ec05eeb3de47bc545186fa93f9954ee604a121686b00d24c67a60608c75186d52ada93e3bcc76ca605a323f17f33c191486d3e1132c9f9805cd21a3c1818654c2eaa321ae136aa567943a2d7f6ee942869b2f38247ca2fbf647313f3f467c75d9b11c50b637e3de4cb097b7f1269e42acdcdb502e2f70b3170f72c8ff4f84c4476063acf2d5499ca3d0431a0fce45b89febddaf41531916be0c84ab2547682955a9864712281651fae54d288a254b71c306e65a45e7bd7d4acf5cd635dbdd71de9c25fd7a1c239bf2859350f753f136a8722f47d0a9c98d31f281586821a06c5bfe8b93412ffbc448645bf7c14b472cb631bac65bce2e3c5391065d3e61d848f882d5f118766c69adcd3b393aadc9b114b4327cd1abb33d2f0b0e3b98f8770c1e644e72ba6e8df59178c3ccb59411d33c838866c9a797432b86528278d041d5197e52afa36b85600865dcfcff13589eb3301b8439f4545a7466137110980671a64eacac33e891ccf46e45c6e723329068409a249a7d442f10b98973cf1069d071d8960c4d29507db2275674379e9365ce91d068ca808a1d94b9f3189d52e2eb1418b48d5b09068d0b9fa819b966ec35840791dd766c2255caa153dcbd6e51225259a88ff1da844f00990083750aa5c8550a9b0bf4760d82f74d4d923740b1fa5ad98ed6459a66c524d419e8ec1e14ca13b772045488e8c8e4b6cf0b0f23be77e35356662d67866cc66301927f67b3a9d1f6fe7d2a304db4675e6bb161da61df2a5fdba22b432d9ed40e409143023837a970615ea07b2a21aea2b4631d15678837b988174fc1adac2c165b2b9a4f71ad689ed344d7d89ae17cff589d811a5d7bc87e53358b3749078c9eef163229134e3389132ffbbf5d65e45b2e6830f9914d6f0902b0a418a784119e92a0d425bcca0795e8280db5685aaa627d229ed76171598fb2daed06f97bb31eb0e4792adaf046b6296b1e05bcdecea65c2a7ce589ee1c927fdb43e1a6fe51cdc0c99b1e702c0bc57b11302c5677d35a8f8e10ac23ccb488760137f93ebd3b411e57f5b38f3750556dbd90eb1c51444b6e5f51983484d7a7cd7d28e18a70eabc97c7597d2dc79e7138304738071e37a2d56c5419dcdf0747101a170b2c11032a50737117c0892d8536d247755f4ba9319cffef0d2047e1fc141c4aaf61c8c8f54a165f4b3180c8b59b37e488af41a73feb16b37fbca7a405ec9aa6515fbb3db5cba945934fd1fc5675760f858b3519f3af021b959509181afccbacc98a5c4f10ade7f50bf3afe62627c730bbbbdb52d73a226a4e635026bd4811c9b3d3f0ffea074e121c514019145b0f52ab23176ba39bd1238ab5773f9d7e0abdb1b4065da09ac66dd32cfbef797e3403fc0d9c275c64c64062795707442651b82745af72d5a586b087ee14f1ada4c0de08892c7ea109cda9315de68b69309f7b7f689904b143397b3c6e74abe84c2f27671054381d13231f0d10ca9f4f8c2cd5ee10322deb6223a46b423d703950eb9428613b11adc5d9743ea1c68d5bf36db2a58aa67e25192892680dc1fa28c3e09d02b114dca53bee983f113dbd5cb3d359c05eb318321cc23894a626b7d5afb78d6b0c94eb7e324ae93e5bb00f8cd81ba660994551fd660d7cbae070c231d1b376c59a236aef6090bffc8f3310ee4f178f0c826b052683922e174c924e0c0b0d42b564144c5e4ad3d3a6b6263ff9bd5f68eb87f93a0cc5a10fc1e95aa51f6d661b0f52c3a2e4935175f811abb80fb8ffd42c4f2ac6e86d954cc719048c2c86cb9fa28ade56166e188e4e60d594f3728124b74be31b32047564f050d668384b15a8bf0c9cec648ff606d6703295444986aec058f32d0ac57f1bdd8d4a5a9e7bc4c93c134adf9e390ab5695dc5fcc641b0a143db1547ecd86ad83a967bfa5aada2d5bfd4e1bdaa934249e184efb9eb2c8f1ab53f81a55e9f13f649f2e52b86c8b38984784124a372df6dae7debb4ac6910bb29a4ea90dc2eaa6dca695e1a2b404006dcf88f53458642abfe3bb10ed2506ccd5bfd4c4d0fcfa338eb6a3057910db6cdb77573ade9d9b8ea006aceae695d6013cb78fe8e5cca7cd15f94b7d8a2afda3d21e806ef693aa19726e5ca5b1bc0054f9f48839fa75634e55252e1de5f8ab2bee06d7163a4c8dc769d906a22f6eceafdb4d156818c31c1a496769021aa8708ae5da5909287fb8523eb21d95954d14437aac9b97f5433d08700a220dae1aa696837f81c1395d496dc34d4c7350dc18a7d49b2a84b4157c5926bea59e02b3f08c5d3dd8a9f47f6d053693541f79f7845793bc08567e9a9f59d6633e779bcf3e3a727b2171ccc13eb7ed0097de525cc0cb651c018f159be388cde05dda2c089f2eaf6cc55ddda5f6db04eb140cdcb338158406228d5466d374b3a05fbeaa7dfe33c8a30409f80431024aa8e6a36c38e8c806ae31c47baf4df530a5518addc65f1e1c203295031bf3da4149179901a7a1b40574cc0442feffeffc8f57407f5135fd73f91b7350af1b9505c29673f8074a1ba776a732a5de56c2d4367ef;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h42d6f9c386920dc73b576a2c64fdcb0a9425b01d4a965b4864753c0d2369913859f46ef6e413f839f04aae19c74e26d093d3900e58718518f96f7335e67fecf07d52afa9cd2cb6dc2abbd5b126aebfdfb6be9cb956b0e1bccced8f81e41cd62fb880c3a8882f566e01827d8ce8e43b36e03f5a7939d14adf8302a059f188b8e1df8afecad5c5fe8db4d4180717a86850860f6533a975267a6a42f774d4bc5918891a72fa0acb800eb066730d2956aea134d02a67c4102dc7a6779ee72de74d5d457e1bbf728b82e484ec21f27a8f5ce3b1561415d7684e4e227da874d50d41b5434ece1066e7f9c830ca38b8249453685a485ec2f6a64bee76199cbe6f17d92ce124781a24f7224b786867e8efae75e1fca7ef4e00344e7273202be1bbe39ffe1e71c13c7e752538cd84ea7b4d5ecda5bdb1d030863f8c0b6d97f1f2a32181c7fdcd9a946334a4f1fa6436b5c4bd21681b5ebb951652496d6d170387c5cc7fb26f31ef2bfce3ba60eed80f1f4106c2bdcb632eed8d9315052b95507ea54f6e0ab4b542a4ac17ddd6da227b2b93076f2c2d7fe44b36a077a76d9f0f9999c7e3071bd78309c727106f6e9ccc37368c32330f86ef685a10d248204305f4c9d81eb7d75b074d6e009fa30153bd5d179f0d57c5712a4f1aca4e6ea875caf6c16db6a37b51176626d5a9b6e528cf2876f36e762abc895193e5631fee35cb67eee4e0ae43b240819215e204b5decdd1152e0cbd2259cbd442da177353f3e64321144786096992038ede5549a706159a2f098f3f53699ab21292c50d421fa0bd2d26c2b55ccdeb764a811f95d0792773fbc0a007e717d2945eeabe34eaacfcd2817f855302df4a8a23007a6dd84d27d4bfc54553b26bcc500a7e4b3cf99be2b073ca380e6e459dfb0118f71bdfa698d7dc795c18e2849e52054a85d57f186d562a7f66e15cf0188bae999727d7020e0e11a55652306f25aab96c2f8a83784d52acdd977a580b78ff8591736af701993a2dd92ea1d5c0b2588f3aa44c94b8cbd49cf6aedc5ea4ff73cfdf1cb7b5e70a3fbf9573e31a466afd326e0afba996586e0df166295b2f5afc20bd56c40bd09fd1643a98fc21a1297214bed2c325c993cb3d33c9d68d9cb173f9172bdca966a3929046d78d07a789692b2584d154bee2b965c167e1a22c641bac543304585f354dd83a0a9345c0e31535397c8e16bc760b72060fccb05a9ecab95b0283425e490966f019dcbbaca2406d6c8d45bc0cf521177ca50db73bdcee86375595bed31a716452f10911cd7e58bfb29f84024318772c0d23216376e686d2ba99b2493bc74dce96ae43c156b19fb26d4ef4d5cf8ae8de2efdc58a435d486a03d10890756e34048dcbf1a262e712c8830c0a1010fa32af49af2a20ed6368e9b12bedf5bf1e8828bbfde36b8b5dfde880404c3343ca73d400d89c3b3cc8a0a1eb45821b9d35b74cf02e2cc472caec39528cfd2ffc2dd2af623bf161b6d174902caa5d2db319ebff9492e34cd9f1e1e4416b3883e32e76cc63b5c8da41c4150509ed7d25a8afd83564eb5544cce1ef1b22292b91bcb42d32637ba2276be856e7939def1453e00949d662183ef0bc8931102b0cb660dfe9e0321dcabea84aba8d7414f5a8d83107d73a63bdc31c104dc9cee19d7bc0c76d60869808d2441d7192632f47bba948f268947565d3afbcfa1f04780a0b66db008ed047cfe1c677ec8ec32a3d8eef7d103ea274f5c873e5853fa0fc463dfad947314dc26ef580c641c9ef3c004ff9bdb92652c1ae5c44edf7468c0f896d87890a2b5663c26d6776e5069e0928a98667f9ca80ca010e7a61c07360e19c07d81b597ca669713325265e6264a81c712f5ce660e66788d4164af3a35f5073e3a9380199087372961ab13e8b0aa777fdec249f9166cb102edb41ac2dc51b9e0381cd32d687f644f290948aac2786c4870f3909455a8fddc87b2aedcc61662800d53258b71fd64075961f39978e6d1ae3460421f0d61d635094bc86ac5bb45becb5727037de019d6fb46ae24c0a6bb5854a4c6ae1b527ee179117ef7d005694ddd81edb1197e2fdfb95a0f4b75579e8747aeac8f8ff998b6d7a9de4bd0a7a3c8d29c99644ea1b927b3f5c4de4db1abd4b51689f195dd346aa5809dd9d1e48d12397e6c057b7c5eefea1c85932aa292de2dbefa2c823c542ffc5ffcc627b945f11f38ac5bcbbf1144fa0e50925f6e47d9aa479ced4fb161470991f7fac60bee7b9a837fe3da1bf674fa43d55b06d8a146f4eda4daee4588da7ace8871657ef7123ee9635353502f860dac4d520961d178a93ded25734537882a0518afbc6bac7979f8f68b1fd3784d4be3330ff73405b798461362ccc1c13eb438bbae2a8e57cb94403e10bfdf42dfa9e8fe861836efd6287381428882cf28c25c045b422d9668a0a31064fe9abb9a01f70ae338d728b561b4bdf6e051a26f7c8fc179a6191522568e3f17cc5ca87626afbaf659473bac07694989f7abafd05e5272d7b557fc8bc89b621748d008d2a2572a6036b007a8f90375347007a96aa53314d7a7ce51b4d688eb3a1770212e532472093fe03e9e138ee4fd15a7863007494021e55a54e9206d28a301ccb7b66cd7bf36564606116fc8dbe805d1f6400e0f3a01f66a0461583cc2b98e2a93f9abc8c3c9a81e08cf5a76c088f3cc42868736c2b859774544c27e5e6740eddace4f6bf3c8089fbd1c311ee8911d20b512dee7fbcdccffeea997da3bf46e634c32c1f19d37be0fdfc01da5614241d123434b5b51604766bcd3cc4bc048060396349ed72a4a41a9f1932356035ba5d08fba478dcde68445883bb97195f488a21789278dea708962a15e1ee0eae242cf6f479b44ca95c8654cb47287a36892a00c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h42093a14a448a4df3bff5e9386b5edd97db089ff5a6a80eb12d2ce5e966175c5433ac92987417fe4697e92356f20ab5c8a8970c82b6ba1eccd551ae9bb1b5ff644d5188d06da9855dd840e026828dd6be5f9954357ac4775284f5ef3f325cbb3cdfc28a97e868cca7c7ea7a37662bcb23ea8ded298355f72724258c216f4e9396cbf8afa75dedbe3846903903016d6b40f566ea58e5db05d71de46507bb72f019315e4a892bafcce8ca23cb43a7d3ae06b19dd4aa5faef9341cd4f57389b5412b2f9f7758a1d0cd1bd18cb983b9f1842d62e9bf0405b8030c2f015a85922e64a6f0bf98baf4f137f3ae0042be367c5b99fcfc1cd4f2ef810d17ff17147a106429e8a3e297ee37a0e6299639f6673db0f8c7bb73d0f56bc240656b5a86dbf4f7be236c42ac43c697c46c58d5d9fea4ccfd5eb36b1135e43db278957796f047f1322e5fcdd50cd3528075083bef7c40f1cf432158daeef3f4e2e740f7a41b0fbfe80ef61903e827d515db69eca5e5d86ba93d215262db5337ea09441316ac3408ebcdc21330286073078e48a53b685c4ec758adae469bcb7ef9d5a6967bdaed849051d1b80a4e441b962d5b12189aff5d872fabc9eb64a56d5325fa23b176527ec382dcd660d19c36b88186c5a05f2f6ee215ff46bb8b21f0b0eb03442b9d775c9603acb55e3e853986b916ed9b51f93c30459555f9582f369f19755395738b1009c66134be87db87fe903349cb11049ae4bf9eaf9847614d0519c16c509a89ffaf58ad773003d990349bb4d1207113d2e59017b754c617e5a006e0aab07aadb1465f62c18cee943a1df84b6472078a41069ccedf25e12a2c93bb3527e8d7535ddd09a08a0746f9b803d93df006e992024c523f7ee994d1bf12081fdc389c6359ebdd791515c4a7a8e3a782ea741ce706ab772df2e584a0b261d8123cc56100feb2c3cfe099bed49aac3f6db0276820576c27841629bf4a9b112bb6c68cbec8a7dc43c77c0deac14762f8309aaef7cba62af9cd344d2f714e780c373291952c15fcf9d97e5d7ea3168163c5fdd57177154fd6cf737843ea46a27360fbedb057c4a31332678c096f7faeac81c48ec5ea6d15ae9bf4e5fa6306ad014fd35cfa7097a22b21f1442e2c631ca47f245fb646f949cd3f59af3ed8be21b1701e55072f223aa7d9b4e419e29e871b333e56dbf6308c9494868e1d41f42384000d076d3dafc26b1e3eff7451ed9bfb4e3b735c15e5d2f1c73c7414f7a8ecf5a554b08b2922c04e9fb1599a5d0cbcb92b468e1e1fa48e48099c244e82bcbba87ec742e19a7b45b19b77b0c5703678123e85a2aa861ca513cc6c5dd55e0fb2799cd3b7bde8be7e6c6815097721cf6eb517e5b2cea27ccf6861593f0cd1f1a82358691c92d61f37a4feecbb7ed7548151e3703c72c0e012ba900ffd71b79f131e8f46e713e6adc9a3436152197f28d8b2458c0f7cd2b678c40cc0bee13d8a5e5b3263dc430d36769ead287ac4c1867284197f9efabac74170d308b20713658bfb091cf7beeeef99464e821d6f7329f8c937a94d5a9ac4e716587a177a405cd393d615928b04ea700b1ac1bd5a71c8ae3bf5d80b5cb6eef64581250c074717adf0b614631df4dde0269b51033bd6505c9c574959d07dda6168cf8f7928ddc64275517d6889a9ee2f798bf30d6be9b2bb168a07200583a0601ab149fbc8b8dc82f0477c7aad30345631f4e62bb3874b61f6e10ba742cd1b60eaa55928351da1f09976eb6ee1aeb6e41a6221afd7adbb8487f83fb411686b23ef3cd390bf20b8b759346a5333634517bacac6d649ca33e18b7af6aae407921151f962b786dfa55d3dd2b3a30fac2ab38f5381988aaf141d93590a81956af8fb4f4fb6e626415db79f1c0a0f969fbbf5c2b2a875748f79b843bca821e1815f37a96cd87d24ffbc6a6d6dc8e0233ef573fb2abcbd3e9c70c0be19d4746c666e43155f5bf78a653ef510667ed32b4d64c3b0ed6ecf188e2300ecf0ea78dd63e9b8798399d35744f3fa07e6fa9b80d919cf04166cb093128922c9ef3c6576a34fa0b3ee224eebcc3806fd8fb908bc67412db1c1c72da045c49ec0844e6b5b9d3f761f2a8021531b61033b2ee4dc83f45544ed37d51ba77b0109362638484822b5e5dd6c5efc5bf844af91ca5bee351e1af92959e6fe8de2f82cd33b1fbd9ef6d6238b84ac42f37a92920a43d91f23a7cc0df7b05da2c1bf625b03e049fce007504613ddf2eb4f64c876d2157f7a1ceece726e366f7d30570174669272663c3fd259e20927b555fa13c5ac17e30f396425f232a58aa71ebb4677cfc2c62e5f210bb1723fa92205c93c3852952c58d03965c5c55080afca69a13454dc46fc3dd7d4ddfb142d0e667fa16cc148a8fca5e83168e698fca5fc1363c929c5f29a4a59ce0b4388336d59f82ea72f22e422ea8f83f3abd3d37159c50102b932fe3424ac650e86d75d5b72e29efdc839503c1397c58d5fa670c6f8aed704fffa65d2cdf512110217ff2739df3a97c4a35bb996d3cde6d29c7e34e105e6ffee232fda1884883458606e3ea521c7d625a7302503f62fbc951c9960e66c615dbb93e927a28b819ad21c9ec73cd7920e2644f97c805f14dc6fa8dadf91b799ce661c8e119994e945e53782be4f4e4e00d909b5c327085c09cd9471ca14ed8c39952d816fa9d77f5e112a114ee60211d3d06278eb858bce3e4b8b5e53c5e2b9302f96f23fa86c3f4dc8489f43b5d4f27bb37ea3848cb929ef4320fd02420ecac51a5d9698700b72baf26b92159b5a8d96c3696c678f106efd5005aa5365aa6e6f685edd61e1a4f4ffdd0c6d688b315e35598db6ef44d1e1387687f442b8b6f35d230856120d63eb7dd8892b07b092d9a1ad50109d6ffaecb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hbf69920286629e6d46b7b272bb0821340cd3d80cbb13d9a9245ce044575b35ceb82f3389f893f5be7cf8299878d612fc592a36e19ecd2e0f27067175833b6ec252cbb471cc7095d1c4aa8b79edd1d86be717cd8db501cb9cbe6f4df7d819a27000fc614d02aa855afd11127fb9cc08e323ebdb9c1b81b5158d85302797b3be8b40ea322eb307490bf53fd31842864341aec8b8037f5217c335b5c4f6564cc2b2c41e9fbe6470053aa3bdb4f8f3a4b25af3c7846caa4e867cdfff8bf6869351b2b90673fd5badf94c70a5b2048e1a3f8c9cfc3db461e76044929ec04978021b05c1e3f9bfadac5e33a2358b20885e0f3329afe700f4322f5f9bf5a47407b7ded8d0203577b37c0fd95ffd7b18e375dd2ba985741d6c5caa5b27629118ff5748a1bc64dd248cd7ce5fb6d9bc2cd4bb3e6a29a6ebc4cc9b9cb8818b034474699cecd9fcefd5f3c19744eaf2b5514d231460cda7e234f81dc27ae558f006ca037bbe84a8bc876705fa2973354c1d5aac743aec59ea69fe749729fa0e5103ff14ef3470b760a816e9c6cd67d6e70f24eaf0543c425a5c400daf63f12b0c884ea469287238e4aa1d3b6a687a1d2e4572b9231c3bc7ca4911aec521c74345383fff89a8737b31815529fe1d0413a03382b6ef8405efb3eccc54724cb74ef1f7ad4f1bec676b2f0aefb11e3d4c81eb1c1c82a16ba3e40f0a18d63d980ca8a9dc8711c61c993e072cf689b90ba9bb9edf5700bb4108a7e65c582f1fe9649049744981565f0036725facae11c77096a701e7fbe9ee9b80658d879a98259336da56832f2ef65d59c09f4dc1fc0b8ade001bbd9ed01acbb87452b4c5a236b784c69c009cfa74e1d947579072ed27f3db3e476d6bc52056066ceaa84faa35d9f8f540430b5a061ca3933001c891962e0aad9f21c79ce6b5285c29a86015a6adce57859e50d24ac120838af211bd37f3cd4038f7ad61ac806f39c1521132409cfef5c2ed32b49e239fc1f3440d9986bc2c4f877db4a5364e1955184824c665299199abf7882a0cf3067f13d928e18077ee64cb1d4691042e10749c8dcb186cacd6232694c1af3bd246e5a8e1f9646dcf3cac86b587ce6c3bcd715ffb43ec4933aab95d67c32308946886b46fcd364979d9c4eb4327ad99faed9e4f18c8963c9f21a397c9b938384a0e383e1c1b00f37afc956cd83550e1c9d521167983234c99f78e32eca9ade5a68298fe7f4730d1533cd4dc415bc85efc3a4574fed76626c138cde87c3afcbdca4e646fb4e5fac179abaf540597a98363e4acc16d0c71d2f26519705c641cbe16ef1eb386e140cd0d2fddfad9b62f93ac08f68fe09df81373a6866d510d17767a2d6187285c06a8a48e70e87442938672299bbd63ec1b153ebf0c7906e2a4de77f55b3729a753055636cff76af3d0ab0f719d0d7c46040fe4c513fff74092540dcc3908c5315c57a03c75d822900313d40aed13dd4e2e53f039a6571cb6b02b0c48be928d5f1763572a3b405a4a0f9d3cad1d72038dc244a48109aa1851deda59d102b71e8277d64f9820b951b11139379dfbe691733bc54d470e3e434cd5b8a9bc7151a69194fc95b645697c385ceee5df4691d95354a7b62a03a182261535e3635351389cc8b10d5930c803d6f8cf5d75634ac66a75430b084af168c53342c370734266fba382fcaee3f6fd331f7f71ff27e3d963a68d0160cea7daaae054bf9fd980d25bf6300d61b608b6525487b969866f2ad3da1d146dc16ce482ec848010361fe8480cd87512097246f407b949396affaa3a0add0a975363c07d6130b2b100d7b3015514c0037664efeb645b7d1b58973c3c64e76878b53cdbda3402c09238b7456bf056576785328a555a78d8b19c5a9baedc2d00c113f83ebd14bc58126db82ad2d2ff33be99e17eb00af6a08bca8dc2728849a260d98efd2b1723c220568d1f236d4f539eb85d413c923f7e62245591ff8bf010fa80e18626e9a61b42bd07a9c8c9e40ceba42259ca607cbfb5864b51edb1e4068d0f561086f25049e59752aef40220b7a2dc55a92bb116a36127174566d09c7431c865b04213631fa41171f64d444ff1f4fd0a7fca1465c06100bb23f2e69658dc829a52aed233085fcf92992cc93e2c4a95be0d8895741be458548ae86c3135ba5ba36c88dc3992c7d47ac515a61fefac66ed962e928c711e352363f3ec9319f10a0e95cd9179772aef13cb4f99f9bdeaf707690ac31f9cbbbcf548cb5a8e2013aa759eb4df6cea29432f409fc09d733eeae9fad5393f52ea10f73811d555cbb800aa4052d914c5f19bb934c0d8ece72bc7b2696596ade8be768c3dd1ea35eb63d82038825495b3a63c2fb79953dcb40ecc886e6ad1041d48a42822a6fb1b25e10a8b40a31f9006aba0fb85522a38243e8b09d255a4562495fecd57ce915256f4865c023cfdd3d0b8ec2cd816ce596b7e2b99f8b17b51861ad9b3bc931a8dd47e8c2eaa39c657f11ff597944fcf43ff946825da0116bf006d1a223373944ddefe43a9a5689d9e9c71b4b09cf1042941fe0753f2faca99e0fbd8137dae2230534a2dee578ff381cd82c5951f6eac2d9a714da26a329fe439c65d659d7f7a664cfebc61022d52c441f48107db051ca9c431bae80dc0877df3c22ea4285d84276367821519f0545abc24f204e9a5e4d664649600aa31431ae3a15063e3d97f5929fb79e4ec896271ce73f420b7fb8664a17a9ecaa749ce2b5057de8bc45d31cb65f02e8425e07d9fb4043f53d595b901e23336ffe7545b314d6d502b7ec30f3491d4bd8726c6e2d2430bdc684b5baa722c21c28a9ddc9fa1cfe03ce29b9c7fbb28461bff6341edaf9d44e6d4bd4015bed44d1fd6a16c9e033ee13f3a6655f57459c360ad45eb38cf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h747a9362b1701f2267340bd792725fdcb25cb8c62af3df88a4cbb8119161973286186361002d4ea3f401353f387277ecaf99e30f205fcfe3fddc67075312d686fd49acd66bf10b6228547e1efa0ae6236b9abb710904e0f78544f592e1266a5852f5c53178497e832ff2471c5ff700e943b1a9bceebc7c1e7d9fc03177eb35949a0a0ee42311cf87b7157cbbd0fffd0e787d0c1070f73cd6756866c7a065c2308675ee1f435218769e960261c3099f507d5c40f95d90abde6ab1df7dcc8ed121c5efb3e02494f9c364685fc295da4beaad77d128ec459aee7ef9da3a2b544389a64a0bea6f838d2642055b11bbbfdbdad0658362e1caa0180f977fd5018756c9256095f04eb6e162a624aeea5769965ab5f0646e468555d40038a8dcb6a44924295611cef64796948c0bd43142d76cf74bc15c469a77850eb3e3f358f981f1b1152f4d1bd7be8fc4362a63ba788a432cad53ce0b4fd32ba5f1f4cb74a4262bd5b7fb4c8b4a50c4ff1b26c6f67574e2a79e43f1a182ad3bcb1ef72f6d49606e42257d29bcb4609ae682a817fb69247374d82f9b8aeee80b0715c3b6389cabd840f630fa9269150731fdb8d6e061b65c7a4e9e2d705189106b373067ea062fc14943a17d5b6ac1b7d6cc920439fa3514cf1269d8f23fff2f5f4661087e9aaa6dbbf10e948cc09b12c18bd2ca9dac4172ed44cd6f967bbc691421f94bb68acd031beda363d2e9c7fe34fe2f858e232af59479ea0e19ec66b4aa463f61d32ac7d863823b83a2bd76a777e42677d412a6147940cb12bd22b0c4c7fedda67e38b45e533defad6c25f32d1ab25d588b4cb0692532b32257ff1843c4892d8b8ba952ed4567b7ba4e88fa4d903fe6c7a19e94d931a2cddea84e97ba992aee42e48e1c8ed0f7b1589733a116cd3aea30838c2ab6617f3e903e22aaee9ad568539fe1bd3945df9b9af91ab6b90a5f8ad1e3d66a58d8d43e51f8d6960a8e1b526e625a7be9c32489fc993fd214b6375b529ed086b50031f73e556757a953a4e8b4bc3cfbd85749ed98b60538672dca5bcc1557e1f782a6fb0bc7b04a30d1678ada10c53e8588f4943bfe560fe97f8ca6dbc28b6c15d8800ff50f88bcb2542cec2ae0085e994ae6fa8fa61aa366c9c3ef6a06db408aa07cc0ee7842f9d41ab891818a1033d755d081ed0951c426f75dcfbc506a37f2d414bd67b18e54f76ce325f85be65c6cfcca19ed6f24d08c0dc60d7401af47e69d670680d1d8e50766ea266b0f4362acbd6c5032017d3798c4dba408f717922f56f9d6e468f09e5fa6ce2cb296b5ed24b77dee70b90ff48a027854529f613bdd00c8d10f14e8246f78f1250af2d1648cbb2f54a7021d826ef1bddd2f2e3a223187cbc14bae57be0ad4d99a28570d2035284e542c4a71dd4abb797ea61552d966fc15e42be6fcdda2ab404903e36d4397acc12eeabf750e5f9a8f55b5e3cb4e7588abdb0773774e38cf32fa3ece018259595ab957bf7e08f4246c26399fba9327f71b2a5bc3ae63be045e4243bf108b028997cdeed347ab538aab463d78ba3d746d9181ad8389ad51412fa392225aecada24696db939cbf47182b4fb78403ce1da053a2a211eee41c853e3b576d0a38b847cce5f2ae0cafdc6913113411c7e0ba9da57bc59e57e8d6dff3e77cca945ec7b10bf0a39ef00f348da7ae609d9174488b927120ba59bb02dc3b2429f9c765090d6382a05e6e26852c6805222ab425141d094cffb6761e2bc9bd04a331e7263700dc9272054e98eaa322c759801e0bc5e8b9065d8b80cb005aa44ba1ddb84476af09bfd841d8744d21127ab92d6e3f0b64fd02268ad00c97611a8d7259fca0b3748ee9bd0e80c642140064801bd7b5b4da75cb6d9781b7a6b1a1c7548b6ee5d0f08b1a3b9a75ace1a9c3b013b24ba25cd03d8d5713114e7e91a9b47b011f6daf0b4eac33fbd68a5290eda4b4ceaa9e0b68b528469a8dcd0d23cd63f0bb5a60d8a622699664937ee039518d0e48186651c94e68897c1ddef5b291c5cb81a2ec215c2fa8d5ed79cd019ce3fd5512d74a807945891225fde2eee116a6034dfd99990661ef80431f258dae6c7bd8c11da16875211c5a6bd018e824752a71ded23fd7c1db8cd6d53be1c48afc0e094d45b7bdd7e4595cc15d4e7f9c428e7c6bc258088eda0798a050670509942eeb348dab1257efb9f03ba556f6baccedeea414a07a7371050dc624a89861f46eb529bcd298be455eb056465f9512255de446f8a15687243e9a672e7173f3131856b4a43a496bc396779f9c42cc2fe4bbb3c99614b29c354452ebf86b9e7c12fa4739f3accd1d56b2c676dafa767fe2c2abe77a101bb000d2035e69fa3be5a664d5c8243d13d05edd0554b8bbd1dbc0391d2b9424c4f4ca96e2da6c2ffeed63d8ff53d45fcb454bc1fd284621fc59edfde5e012c7355ac6ce7276708e9e66efca7765fe2e54b658e5dd36cb4a706fa454f60fae84350adcdff0bf21246b2a16505bb45f8a3a73225a46760e3b9b4f360869a55ee972997079da62f2c8892db0efe95741b930a66317c55b619d1dce6d55d2536d94fc5f990fcb309c9b73e3015c82b9b659ce5c51b57f4884ac6d31168df3aecd056ac0637f1717218f2613bc77b57fd63cbd4f1894a474d456676181c90a18b0b68fbe78a64c83447544fc1ea3375124cb2b8b1fed0bc7c8cedb63ced89b336449f8780ea497587d1d2ea788f18bde9f2d388c1e3fb7a3590401275470cda79f3b300321acdd0b8cb1db1859fc066312317c0103fd34d35cc032799ca589c62c6285facfafe6d0160e87d0a1011723ce91cfbe2934d077e75506506411d384769ec8812a814af7ba40b892c8d217b53aebf158718619bf27068c45b2ff7cca7c030d00;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6810eecc50fe91b33314e4a45d0b43c44fa2cb2a4a2eb22d62b288e8da9c2eb9a874a25e979573563d2477c73b8d12cdb8a8253a7ae671bed946ab4e08347ee97e0089cd88da3a63f920194390e68df54e95a3a3efe37d96a6367bcbc8e516ebb924a199022fbc7b6e37494ebc3278fdcc13819cc59d288b7d30085b4a5609fec566609ccdd0ee87f76cc041e4960810d048f10442e5e77671a577a5fa4a98f4d93307eb0da4308ed2a4b721a150e40fe88b0ee50ab3a1d93f7524471b667815869b928d8fccb13a56f2f481a8795e390f75f73ac18bdeb3de1a365f4cec0f1bdf1753c3797eeb8d273da6272662747e6cbba812ebcc0949772421ecc872c0acedce726b8016db38d272edd03b246e326b4366ca1064f845d73ff2e704b8a6107ba43fed8d125d8a5ae3d0ee69009f581a540de3f1db4ce223ee32bc7f6b2c90c91499879b9926a736e605e362e44eb3060aa71c5e1bdff5014e917fb43db55d0f708b338bfaffd4097c4bddd63d167521c808eeec3ac2c7a02c09abaf4957649f851c76585806a57c9f29045260b2d7275790380f77cd78431a2c0e861a5e998c9412273dedbfcf15f3024210ab62543a6de01c27aa360e3f5c66dbbcce135ea89edd94fe3526cdd18fac91b81d04b4f167afcdc6e3e6f2b2d27b9b3df343fe9a8af56d883206641b69433f9d047e0430fedab800b03b67742c71d2e0e3d03608a58fb05496d9fed24d67d5c35f3eac2b94f4ffaf6f2f1ae4ffb95bc3ecc98c96b9829c2d8e53cf1c9aca8da919736efe32e9aa0cee44e594d417c812e3c9584a651f8068e0ba3e6ff3b739c47eb45065cb8ef8ee23cc477906ec9f881044425233fbceacd49b7e971b201256526f7bb8611a8057b1c92a33478190832f71907c648cd3b9b4f1c1f2de41893006c6fbbf007aeb1dcebe4ce0151679c18abf028d5d05f3a9b12b061f2428e1d005b3062b832f2f5dce1a34b8e9ca4444905638f1f9a1ec1dda9b9cba3896b17eadacf90f6255ab074de19bf3671872279809358f8446cf0f970a3b1abf9b018364999a8ade33c88101a338c29685fe20db7d8a6bd2e69f0b63c1061d2909e47f58592c2352850307cdf884586a43dcd29c8f5163f419a0c9e172b9a964a88b8aee8a96e28fcf330f079fff9236df2a59a449a74707977bb1cfa7715f0c6b2c3712a6b3708262452c70cf9970b2d1833fad47c7ef20aaeb873e1f4545d1b81d685618f0708e8f1f0941c47adb4b004cd93005941a74bcccbc98ac710732e31f964c3881e6beb98b812de77a9f00fc757ae96dff09e9f23465b47f1d8cd3837a5ca8bf53af4e3ca8acf7c35d0f299757057c9372d2f1aa05a1130349559e0ebe11d443dc6184f8e04d1fb4912da471c7f939720a3616b58d401b72b19a10094f08a620d70e8862bbc283faf53163173ccf2866352fe5fb34e0237ad1456c54c55702d8a10fdfebbbb46e244a9a394941bdec802a3eb7e526468d249b6603542eabb7bfaa3ba93ac59eb73d34e7517e91b8c66adacdf6ca42247ffd482b1d38dce4bc4ea26cb5aa8fe2f9c2b7f4baed5b70090ef052f11d51a59ce64fc30553f95d05842c6de026bf200f14a4a96594e52b412fe5272b5c519ac6352f0ee3865d8717a44f751bb9dc6d6a740b1b073b1b987ca5a161001985eddbb803fcca61cff21ce789f8c7d30bb5163f3501435bf0a2abdc5de5c87112670f8ef82aa427422e8a685028cf41d1d2c02b470864976d3f1c18a566fdaa8db5f017d64688284483f539760af532305b32d50b7373621fdd8887c0d6b48e5c43e3ccb55a34a169b99eaba7537a4cc864f5abcaf5f3a3f00bddf3022dca05bb3fbe72a121b3d406c0d510b76083fae1a4724cdfb7f7655fc094c9aa5db29f2e96e6917420e1d93a80fb4b8774a8b651a62715f8f60694b6ef65678b90d4caa63109c66aaa0c1781633e3b87c368341dedebecb7b7b96d9463211dc3cbdcba9be9468018916a4fe5ee5b219286e95cd947a80107dcbf9c952d6e412d9cad5dade548501949ed8851bfe2ab92af1670599adfa133c9d6f13b53678e5a5e452ca3d5491520b5059e26f8f233d42849842303e3fc47364dbdf04f9b97be2748a9704740348c71a5f8e8a15517665e9be731b0dc3862001566b92b18dfdc252625e68e50e011f58bc3f7128c94bee0196c3f1d0ad7ec4f43601ab49ceed18eb20f626d087c46ff0c41b6a05eb2d6816ecdb45207867b7f00d055b24c777e5c60b57f46b4b2ef3570c1971b89fa88365b0911d188fc1fbe9ff69d52cfcfeae51930b508cf35b12c450310f3b3d51b5c79461353b0543ae89026a09d419a5d25435c8aa378c35fa26d2eb75b4cb520d2718b61f23743fce25fed361a0a3f800f4ff6672edf79c3ed528a050fc78ddd9d47a5fd0b321f87908191cfd060075059fa73f596c2423b76d61f061fe154e580157f91b2b7619cf437e6e4d079586201875451f0c98df876cb5caf5c95d5b24ddeab9a7925803367bc03589f4b2126b979906649805085fde92f85a3eec51e9c5fe4ed12a76a9d28d859c5a023ec03caf50bd9674fa7175c33bce1a52aa8b2548b46736e81bfc6cd39e42e1540c9714b51bb93309bd953979c34e2f00fcec24c5c5285726220f741a20c320a1847d27888e61cfb54e5c118d8f719346deba2390631c518af67235b23e2018e45ad3ebc71221543692e94feda938cc1982f905ecf9e5aa435ac8f16e3342abea0a68284b9fab15ca658f0bc053388cd8dcaa2dd6ba24514b8351b7f397330c16f0ed3a1b2c8281b9773c2c59a502a2f1bf49d9b55ca8ec8a4ff62c39c5eabb54dd62e3726d75714e6b0af9f71031947d0b3165f8293a50ceea90098b6586c85395410;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h225002defccea41db08495fa6add3ee674a21bc888f382850dacdedc239693d4a59d8c6cb5cbce25a3bcbde64bb40a30cb7773a71b79b4d48f8be728bbaaf0521a118d227cf1fb73b10a2018d38d59959ba038cda12b35d611d246db4018fc00f753f2498de9ae91daf768b6cefc6a44f4ed8f9341d758d078de9136c376e20ce15a0bc235adf446656b7a91773714ff79ea3c70a2efaae9432ac5f1f17929f0dc8f6cec99d9ba8f78d8365865c2524852b84d8f8853d4c9be2b541b7106fbf1f49d63b8a13573696099f07a4dce18b851dd12b644a86197a49247679382c18e84fa64182bde9ec1c14b42fee6e43a7347b13e09a6f041145f36f4da9940344b298a9113b105ac2e1a885240b18751547015621771389cbd4aa655db74dc2e3a1abddd35ea49c22d933e5f4e0909aca62b74757dd70cc4a2e3508ee80874f1ca7a659653745ec7d0b70442df8c6fba1ad355e50a72df2650180ccb912b2f7bbb7d2c2cb7a23c330b51f9b4ed4f03cf3a7975c822ec3eedbd2565ee00c321444415bcb5b6b204c1fad9776661131b7aaab21b274745ccda7d62b979b94762354c3392fdaa15cf9378db0e599c7d9ad6be2ce2e6b80ec9fa26b58be3a1b2a0358f4d227b64702fe5814a139d372752118dd768caf2c8d277a56bf2398474ef3124f067c15b88548f2de4f61ed660567694d828126a66bc1b2fe74ab54d11c6e471de8a4643d3f02f099651a89650f485b635990df3cc2e8464edc3b9c22935d6cf37ff413659f35f07afe8bba801dc69ecaea3490136d6167da652308cac516e6d8ad6b0d36a2ca60516f2d3fab6308cfb84f4cc50bada858d51c40bf16362c0a342b07ceec7ccbdbfbf140a560d8f4127756c22ac05d1d282e9e090a4c355945f5e430dcdae4a990094fa155aed15d208c590ff3147de9f20e0286edbe7f897bb5863968494bd7af85e259fa32812a14100bd4867f772cff1dc47bdae08a07d5e834b8ab14a0d2b003e4ca09119b7d44d594702aa9ff667c7a05ff2875e1503dfb7b8c47b5b73d90ed61525f655fdb1ad930df35b8b0d1631e03abc50cfe2a97b3a4eb209e1f2b2ec6278c71c3f556baa3c21d9d3e4fce536986ed8e367b545f1d215386e3a9d0e2a54aa53a34691e7e202be983bdd0138184b1db4a54bb538f332398c1a247a1870ca047509b7b89512662ff6bc4adfad367cb334c6564638e69ca392e961e71c531b05f615f025a6e4b85a41582f52b4f6db9bab949ee9b478f2e4ccdabc077d89373e142b52ed6b77cba55bf88d1fad8541523decc4bbc737300ce06a548a645f1580f03ddd3dd013004fb0cc0728ace40c2d11e284654e98eff8d416b8b2552c9da094b55fae6b28407301d4f8c965ad088fc8b161482b1da5cd5a5be3f1d4976298b3c92212cb6236e75460ffc7fee39f987b4b60e551cdd9d64f0d173ee85d3de48bc79782c70379c1ace48dd8773821b185944b90f7cc3e29bebf54176b7ba1b997e75a5ed4fecd888d381eac5dad21d02ba99f175c473389de882f2fce16d19d0c34ef1306f260f94a3e70f3cd05301f011a41656587d16d1d1b34cdf46c5a0517f90f68198b9c2679c6cadcfa499974fda299be835711141be77f163ff5b3e39cc9881c8380e450dff53bbd250d4f2fcd4261761790e90a3798c7db617d4bd514955779819821e1e46e2ead0b3db13d73c455f0cd8bde5b3fdf5ee2d4fb65d0771f414d63bd9d962a7cbc98d384761310ea89b25d64161f209d6262c621b63908ccadf043e3bb2515361e1ed2fa8d549ac62693aa328e6d5d360139ad967dd27d2e0ae3533bb1bd9f7394bf4f87fd16c428e471c023bfb2cc998f7344b9bbd4bc2a17870ef1a595c731b679b7d9e7ffcfe2c2afa4968bd4161ae969f0078bef05006f72cd3fd31c75e8698029f22ffcf284962dbf0ab1b223f4d9045c2b7dca69fc626f100a95294090dbe42dfcc790705d713f2cc14ed679490831f9ee81072c714a1bac69077f7a7cfd2771576cee7e765e6f9bebc86b3ba89419d7b440f0bf9ca84e720d84e30a2845d6086a6f2ccecb295efa92dce7d547a285b03c16b790beafe46d2da0cde382a986c0484d95073e96278fab2ef9be759590dfc23f54720f17485afed7934f095702109f02c59469608ee883c56c8c87c1f2fc3e2737f10281e2e8c7524e49fd2771fdae7cc73997a4d58fe41db9f33f15bd36a6a0398e46840421ae0e5a3cf15d7642c175714cc4dd23829ccb56a5478dd4e6e970d33198667194e8e3b0feb5ca257386f0298265ca28688ad63202ba7d99e672f7b9bf150bc50109f510dec95eb4567c1da51f4175d7f8d33de7c2c5b5af13285aed990031daa075b47a40355d8ef4d116b113c7e08e75846fca5fcbce7cc55fa1b2264b139dcaff0a53512820270ed0ee842d7b5681e8473b91cdb9fad9d49bcefd2982d87a192bea718e6aa9c7b908227dba4c44b309a0d3176ced96d927d759ee2afede56b95baf835f394742f62060b638ae0eee4f0902480f712f4a778042bf3405416ab9a1c98188a62a9a92aae580d8c3433a049737d47aab1d78039b5136402ce7f0ecce2f66c00dc3bcb63b2f1cd4c683941b72543ff9855d67c35af19e3c092f78588b52ed58b7a165c6b24228d464363964591a6fd1069226fd235dbd3516744cd766fb91ea34a4a51e85886370d205739d10c1417ebe69b40e0e4e1bf8b02f5397c27c4f3f00a8807f8755fdae6c7ca5d8876184e7921c34b4e450b6029ab2777d59fa7e96cd3a4dc9cb34645d973c42434a4ac76ea7c048ee44d86472f1c139a93349d7f9a5e272ca1122b5c0502b3c778c811f49796f8845eab2becdefc12cd06e3f513fb90da725f607fd692c73a7405c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h93a38b09375b857b04131a3eb4269b64c3929452458863450a26868f3d3d17ff7a4cdd118eae508b08aa0bca95c5aaa81ce0c0076b6ea183fc07fef6f2bec15e04632b1d88e441f6c126e6c02106e7029a907f31b780e06b25c91e75dcf9ed66f6ab34a6b5e8650e84235fb6cd2545a32e97eae406d6ff1c68f7fe9185b4bea7e1e363b09b3377a7f420df8149179c572fea24b6bd0435ad771e4960e2ad9b5c01ec23fa51fcc0cc612f9e855b39121cadaddf073420e0ea19faa20947b078114801911e16a4a7dca00141c9afa13748c49183236ea888857ee6972b763821d1078d7ea758b7ca619dd6dbbdb081539e4f8b9af1dd0d3575af369721478277b84c68339b07b1c13ccda686398bbe05b811b692d9aa9c81949d58f0f984f3af29280b92542de6ad7185ef0ddfe818ee4a24ee060add5e70a2a6efcd63076dd327fe967d7ab28d34a082e2dfd1352fae09f5b44701c2c2c86aa1aca95c96e107122f9528666752b85237ba48bb63bcfa25478edd5263cde19d1fb3ba7ac48d8fee496a51512d79b5d5a8a6db4ad55993ad8353d0ef707d8a3b92e283bf35cccb1456f4d3be0e34a53f9da7ece8083be46c41c1ebde6efc583852d097b09772383fdb8e8d8492efa584245fb6aedd5123cf9d5e70e5905309c16ad149d57c5cbd57296d102147b92f38f373e2b94fafc0672be38a44cefa1fbaa77fce5326a729f58315a7f0428cafc65bd53e4715a3852e3300dd08d63dccf045a7b7810f8306c87c693a3cb8ba48ed13b86f9fb6bbfc29fd7de1e46e215fca35270cc56b03d03451fc2bf3163a134836a61f108d6d505e28f534d353c75133d128eacf92c72f4826468fd87ed8f61e3aa6b733c34395095d8fd176c0e304af4503af98af96d7ef9545b1de23c7790edcd3e6fe221c8c9350c76d4a8b815f4e9643fa411f73ef657a93b15def2b6c4ee640eb91218ba476bfbca7c8bc8c5a1a0ffadea4a8519294b9da3f304d467d11940d11078b56435bbcea33bc6bf947a640374ee740fe48893d031a9eb3f81aa1d6d56ccef7372aaf660abf0af9c8ad89654c3bd1ab83e7f339686c071ee3778e5674241bf43b309a0bf20e19671419053b1cb65e0cd23696db910dab63d3133eb9f88e48cdce00970a943cf8190674ff39724dc08a009faadd6710dd588ceb1b078f135072f054fb06706690272d7030d69ced6a7d879c72e7da430d0e637643bae60600ec5f1c76989318a1f6e559dec60a6cc22f8e201949148929c21530899089e928dd1ddc98058db6fe6da3d7e0abbaed5c662ed625bf2ad7094a86bfeb92e5d0000040f641ba07e1d95dcd9ef17fe67abce43b912792e914d95f5fa75cccfe5108f81d640ac38c622827737356c661fb3940fa478606f04614d05f928b1a31ce7fec5ecee3a5770f1da53b858718afef3f9e5c478a75341a0f3ec7bf039e4820b13a6adf9edcddfb8c8068405a6cb07fc74687620e4f621e8a3acf01b0fea1d3076f2dbb549bcc8d70762304729e4c4e232c279192a0f932d6447aa3002808e278c6c472fded905dd19c381b2f33379eb548c9d2d3a20582ced2c469fc45eed319eed1c508d8045d010e247fc33ed5a18da0af39bfb12ab9c2673130bcb0229244cd1228375a67f938c13b25d61ccba7f452a44c0236430d4b1a7593b2d369eb7674d5350ec182c943843f6d1011d753a05b0de3eeb7368cc807eef4c5ba9c11e31136dc587d9990de0501bb66337ebdc154f32a41183549949245118407d4bd3b7d05d838dd8f5bedaaf0eb46b8862d7d3f1d435ce677b312e562871b1887497a49383604447911e6d14acbd4ec93374218780b980adcdb8493ecfc0973a6a414fa2ea9d7f2dc25a04a2cab8afc6bc70da274afa00836df86fb6d253d7e80e94814f11e87642de7158fad8750cf828ea7dcd0fe3d9dda19975c7789907a2ae91a8df200741be38a4b5ba7f308fba4f3a3e2b0e57e2b5c1a88bd5f67b65bd47b0b845f9dc0446b0f22d83eb028fd2109273125626df52c0511deb4508bdfd58e4cd341d91d40604cf210c28cc336f0a1727b08eb48d8e88ebbf8582f03b93375923777a13f022df41c9cf4f13966ccc0a21fa7272d64c033c20a2c4582fbfda0c299d350b446e14149309e8c91efbad3a084c6dcd093bd0fc8acd4816f7906c7bbff744896fa6edf2c05f2aa682fc0d8b5e8489c849fa31e0c333a0e6f3961fc44a9ad89cdaa79376bdc90629480450161362b01373ee96d3ff314bbc8457c12df367b492924223538c9578c53ce0094be8da2e37acc1d956d036838ed0156d86621ae92ebb4c841c8cbd9aff2c63726ec73589ce7de478e079f16f43c0b2f5a33ea1d98037d6dbedeca86192d1a5a0c1938338e3026a1b85fddbc52e674756ef820b491629c0607bfa1af99c698a2791538c5531694445244c9cc55864e12acade8e7e3d1bc8fc55bdb86cc6cdf204762dd8928f81a01cb9d51c840e0700d3a078d800a8199332655d21a70b1b1b265b22b94e817665e462fee5e051784f878025ca32d9488a3e80368146b68a3159df796e242dd00556497038e927e17279d47e39d458627431ee6acb3778beda2a08eed033e993472c33ffc7a41ccbefe07f3a09383aeed659e3d18a9d4456abd50102c2f186bea9ce9b4ae950a6f1237bd069e2cae2445cb7ceb56a6ca059464e9676a0e8730ef73f5c6b30b0292701daf21f16f222cc2bf7ff8c6e1046f37155612586f2fd08cfd8d59f19cb8ec7679af8c77bcbe67e7255a08758893449ee4ea9de9aea02f8c4410e8e5e5d0a8628ed846036c2b424ee103e9b17b6150fb084baee4a3973870f6b18ea8a47d20c8d2b5a9b26358a9473b002181875ede3ae52ad09f480cf0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7de7a68a762c168f58a4c8cdc081f735c6fc5196e00dacfc8ad60239641afd3b73a5ddd0e6e677c617ff5131e5f837c4ae397fbc2d42725669b6d254319e1bac81fa40ace0b6240f0f834f1de1bcd61aa6fd726e63a829217b332dd5dbf08577da392e7daa880df71d9eee23501087dd8d5467f02d8716653137769c1e747952a0f09276cf38fe617933a5e90d277ac34e2f8d74fc99fe2373daa73c92d7b8fa9cb78749bd7c2e47c7051b900eb4bfceeb243fbef9eb39f438b3e927ab0b57df76549443f3074d6f253320a6765f20c9d91426d11a4e8d39ea4ab47436d85e36a65cfb7d2acc351257ddff43821b4356f4a86f56a8572e9d1cae82c224954b4d8faf9c6eee05f74e50d1fa3cfb751d2e73e12a593b8d485b24f918e4e16cce7de0e3f0070ada82432b18b051f857e54b2298e1df67613ad99894033348c4e7d2eb49f324cbdf37c5d5c8ce4fa6b004b969535fa5c44fa8e0dacb92745fa796bafe2f3ee373f2bffa3506438bae0eb8f1cd637b774ba0d24d0ffcb599fc349f3d3b5ceb066b50bafb16c9153a1d65ff781f10ffa1f7e4be01d33d7c9f1efd4569126a4fde4d5d5522afdefa4e35c9c40dc32e50309580f636a8c5e56a00b4af4c0baad025b8b4ae5c31e84184f4350e9a268a321dd2762b2ae5b292aee09ae5b047c985da65aa4616e09e2167ada5cbd68375b18246a8dfe1deb9a0b040d96d1267a22f99ef0b151ff744a6704ef7d8dc69f6a510e054e521b8391257af9fb45a34d192fd7b78f496f3ff7d89447f5702c68c0286020d83afb3d50e8eba73a4102a29c0f275e019125bc400c866b21c9d65a4c9dcf9c3aa8c1351c0a6ed28cc2178638f46cfce76b263a310818eeab319a7dd26786a3411f3b0161694182d96b83b06b5dc5776d72c3985f9b72adff91a0cbfff6ee2de356fb5a6f350d472e2fb250e0175ed4846e814be6a733f0cef3cb2d466a438c51ceb8138c90d45070525a5fd30bf735ca9f9df9dfe154fb5073f23f02408b503a60a2fe4d2a001383af0b31e8c41f001c2b75b4f10d0d0a103e665f5d3addfd907c5ec95c54ac4ad0684a83a8cf9fe523cc98cbae24415578e13a82f8e4ad1009f1616ad55f506a696af25b20e4eca53631609106804c580fc9b5b1ee40e999776db50b3c3701d3766e28072db061ad264079acc173d0052225ffb351224384dfc991882328d651989ee6101a4993df138f63f40578757fbd05f9e5a59127f942f871242e60a2dd9b2946eaf1d9e4ace83a7ffe8e9f9de315bb490777928d790cf737b0b7488f95dcde2f55ef26cb19d4bb28f9c0470eec52b787577c74b5a07d3f2155ba10760bc4f26108b20abfdda1a1109600291acc4d9257168855611a3330666c1d137b9fe183e6590f90c7724e37d8189129614ed23f54ec1fe71e57cde414abda2d7338601bcd60b81859ed7bef9753cd121704d92d6773e081ac66121b2e454af3507d09a1753260d0e9c4cef6746dc5f994ba709c6d9b9eeca4c964a10374d782dcba10fd28159743d3d4efb5bbd00189f404372aa85a9fb08934713f52bde07df4cbd9bde8e6def3bdb70ad0edf73b30b10e36d7a39ebc9c76485ad602bb876b545a80a56cba230234703f9fa7c40deed22a48d014fa0f62ece6251fa9d4c238034e6a09ac2c7274e41e0fb28fa8e322989127d8ec0d5645232fb9c0f72f6e90c5c2bfb47b532dd7c8a96a1bea3fb1d69d297cc9269f09d070871fd4fd98b7ba56d1827f44bed68c290919fd04b8a7698c638bda31963d70f7e9dbd0a4d8aa03cf165fca44ef6b3ea8ba9bee200cd61955048b50db8a54d5ad1c3d63a728a03560d3b7eb23d404c02878bce7d16827202cea0d0836efd2dca88cdd2373d93fd7fd3f34c1b923f1c29c1b0b47cf8871ab32ba273ced88ddf2f06d68db4913696dc6623517be738531fd971031092c13f624e4f5dab337e5df44046b0b9d39307376e84a9abc2acb188c69bc05db6f2219039d87be515a4d7e06c602048d30ff26e4044b3a7495143261587009d5c53c025c4fb43e72aa9a73e87a72b4be4cd8960b85530c0c1afb4bd0a79768c40fb89dfa45e87ac72c30d94c81e771f360dfc6b5ed0ac50bad04683ae610577159b0764c94389bb0074b54bbbdc74b7dfc89559e8411f4145efcf8a13b22b7c19c266be34993baa2e34d5b8d95ca1bce990400fb45a6ca31332acfbcb5bd2f5517cf5e83639d0846fa34b2b44c79a8a07f26bace74cdf3a2f351e006bb75367afd8c47ee7b9fb32aa21a7250c07357e67b410ce47dda66c7854e426f84558d8e88e3b18fbaa7f8fa2b627c6f51d7aa06de28fe104d5987a067a5c3975b6f753537da0bfe7f3b4e8d762701a840704e084ca4822abfd1555893cc053da7fcd1d73d28a287c7fd07be8225c3d5ca34bad31b73e5c6130502be5a62362f59f7dfcb1035192b6b48219feb52ada6c3cee069b86be02ccb0cca8df99c7c9358a85b30ee858182214fea6e821bf8860df957078d45e24ca99d855682634c5e7ec6763a0f5ad1fa1ea22cdafc1943a66b634e2336341da50a0df20ff86046bacf56eb1a4cf041bb56ccd034548a70a86db0111037dde101c7917895fe956449d6c4993aeffd606aeb4ec48e1cc077d069b3c806ed95592177a02e4954bd997147a4e85aa8fa378e4c6aee7cf3aa62102ceefa3c4ee6de68a2d5fd63cc74f894c7060d8f621686cf3bf3a46348c5b63544a857cfe74dc924748dc68e19f13f56a17732ef00418a93cf1cb7af8b98271cf55814bc226bd2b8fe7cc4a52d7c6e0309618aa3aac8b03dae8d23f4fbfc157dc8dfcaf4547324652e4dea6ceb54fec53abf19031e39403f3ace8a9a709c4db6519786319d6662756f9fb44;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc4839f6a80ae3c6b60955a9a3e259308bedd737667efb1c9590a3dc8e5180075b5ffdd6ebc6c1d175cbcee07021f94811f44fdb4a42257bd9c4a1b8041c88e99a72b105cd75d80f7f3a25ac3c2bcce5cd63a8465e0fca641aef19c7a52084bdc17ec58f1b07641de5c0b9a5a8169bb9e8a00d71ca316dd9b297cc9717f58f059e08c781d37c708b3ae7cab93a4e4c7f7f07b36d25df678ee8ee85104dd3cefafe36bf22bb672a7c3b371753635f31cfe9c5091c61c21adc3f0c5f7f6a29e1379be23362c37ee2bd2e31e200a2bfe173676bca486606d0b92726922239b2f319e5e72619569f9c55c3e56cb4270939a62b0d619cb011892353c53a27d3f5109b6c7c2652bb2ad5d982007c4b2577148645927b3f9424e43ac3c95b5e86e1e8b493b84cc2f9d5966a47694225ff6bb05db4d36569d27d7e16330598e6c658b9179d93a6ca4e305ceb6597e68e58dd41d09248edcf3842d2ce4793398a0648ffcea93eecc5861f916c2b8e1a554e132815433404b5d64ea2dfacfeb3ea74f9ff04bd74eeef56ad79201d95da9cf59257ccfacca9ce0bd6aa51697c0dc2c2178d07251df858ead39694007e7e519f9433b4a6f7cc4f97ba74c9286c3eb15823616ced2ec34d938eeaebdab970aed012c704e47d802f1622f7b6b70cd99bd689998dd5bcca1514c6729b7675e34cebd4bec1861b5ce73cfe16e3af3f7af470108b08c02977258f4d900fd0ec25d20637ae5956bcc5d31fca782ef3626410514bec143fb91996b47e55aebb6828e1c068889394c60549124076bf506d341ef03c82a19b52438648531f0df6fb33f218db9848061db957050709cb30149139e09bdeed5f2534334b9fb6234794d10e3856e565fe29a4ad10108dacc099f840dab1a4f13d2857ba1f1e58ce09ce35150672eedd7aff5a7610b6dbaf4427a6c9f78cbf772efcc080c169ae2388db1edb51a79aabd134d8adbedeb634522675e6dcfc7af0a91206beb02d8f3b586f3f9dbe61c37449b8b3bfb7f593c919451500256a3d857b593218ed2cfcc2c482f10a98588a5172ea30def9f36eaa57402f8a9edc662bc391151aa4a135cd50db183cd89984aca281f56cec15e53b6eb4ea9f0f907aa6818e5b7b08dc40ae960e2447ec9130e7a5f8d689d261207ffec1c780bfb63091ecc27a37787afc8d22eaee82f5ff08b2f53b7ce59754314006115b345b6489acafb8fc3ae51195ef9c29727d825f4b6864ea7b476e2700d2716b43f8186074d7c5c099651bd54edecc93361958510c92a22c63b01a899103ed5d400c566d9cb41e0904c1d0c3fadd3eac4419972f4c9cd2bee33bcd6efdbce72ca2f43791e6dcb7ead9c81a18da99e7cf6d6336b12ad5ddc2275babc70bb061f09ae56099ab61d53bac229d126703044156dc1c9eec51d2ca9313eac6139e47ae7e059a6b5f44305a472799bb440581e7760846932f78f10f23071dfc19b89fbcb1fc08f850e7130a4d82b7f27086d2a40250e1c28e60b89197e2548320380f9947d07e71b3360a70b16d104400cd0005cb6bf8011f5e16ab4f81d132a24c9e74e8c6bf5a4df62750c6b15249cf9fefd618fa853072194458e293bd0892c2740c61163f189be7b18c3f9fc59a86f026b47a15ef4346db719a7e468a054cd0f6a29816c9ca71ae0c277080212cd404d22ead8183bc7019a05b270410a5599e57f73007bb341cac1c661e620e632bfd79233184eba1bb29bbf3a0baedbae06ea096848c8db2bdb2fb665b455d40384c511f734d686e574b5014b04edccf8f343b2f35de5d84581f550e3cf8ca2fc4cc6ff2e8cf106a264204ebd620c7592bbf1b627afdf89d5ece06893b18d07efa35a651618acc037b2e236327a9f5df6ecf808cbfc6dc30423455e553a372ada0b183cbc39ddc00165afb7cffc4d25c2526b2d71a39a7c4447d7efbe375a60e68b24b499021f8e0ce4cd774b46afc088c32fc0b015ccdf16b7d0883c32a08db3585d6b70e122188692b48e1880c05d2fdbdfad46bd69d8cbb49d996732dcfab97fa4fdae393099a264640e8a63d0d372ff54f315e604260e3f392c08cb1154a1f3d3a394e1481456d404b36d8ea6f2d836f179712414fca918d262554618057b4d38015ab930abcec30a53594dad10a282f2057f0f6100af5ccbc5000f99e2407ba8ffde1bf87d4e972c04ecb6f65707f15c8fa678b8c410f3b7f2a81958e14b64abf276d2060ba97f81945dcff8641accc6200048038caeafc14048ac0c779030c7802a83d8d6b270e27e947971fecaf67027f42aeae221cd66a68cf579a95789698dd5127288ceed39a676cf13fd363e998646844c80160087f555af581d2171120aa04a340161bc67f6adb49cc994c6dc10b09c84a9907cef36fabf8462c2b4eea6cee3ba61448bb2663602cc728504f236449155ed946aa6813d4162cc40ed779c2cc8dbc90fae129d9fe629de20b1e7e099bfb8eab0394ba41a1519b69c9e97e1c6bbc5fb75b16ab32ba58b08f4b520b079f4a317992421c0d7c992b4d7b163b1c76cc721b381bb455e765d1ed7e1bf63e4b69ffbee6ecbbe04b5c3bc3e7a700f9f621971873550c847f13da2f9a7f797daee69756f083c325649fc09bd71cb97a52e31678857e15ca7cf51464725876d8308c491d869d2e07f074553c3d4600aacff783eac337a5c596f34f07e61ab8507fc90602ca5c7a3374254d2a47983f79c4dd864be86d68bb1de7359e253c3dccdb1309b05863c8220d76cccb406c4df167cd937358c728bc3c4efc4f0d230cd735cea051cdca5c859a6af7654849532e73b3fff388c01c27cdbb73a354b1d7276bab037bceeb8aac065bc227bff7cc9dd1600158e76c0b69365ae7d0fd6683a42e31468f2ca36;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hcf99350a4d6687bcb2dd4cecaf7e27ba7eced162beb105a2adff0b14bba8c71fe24d466508440305889902dce4dfae668c4657def1cf941233e1a42740e2e854ec669d7418c81c52b99459edd7d36d436a494c756b2be0dd080649faade22b9ced0e780493ed86ed72d648dc1814a033421a0cc8db982b1e2e96f8418ee124dd557d67cd72339991f15ca1daccd5fe1b5abc55921604e2547841aff1dddda1e312808cb0a204f3bd0d5e5424c75ff38dcda6c01e70bf3a8705918504793fcc9d6205c9248c39f30c028b883c77c0a656ef05446577078938f201c8bd9423e4b827a56c073507fc0278500baa21d243ee00588c06b6bd0a93cefaae879743aec0b52e1a9b30092bae2dca40c0c8c55bf8ad8a2e29601f33a508f1c8e8d3f07711be4dbe8efe57430a1454d3a89fb21345188bdc7b38b7fad88f0121f6f4f44cbcd8d2bc75cbc1e000095a60b88d8b18447d9323fc907c9f2d945d1830bbe04d3d02abce8562d40712d63366c146a6dc4e40bd0ff2bc8a755ba218358bd77847ab68b6735a7f95d72a798ad7ef9ce9dd989bcb73fb4238aa03468e46d59fb5aa3b60834ec456cf7e6a56d62fd71e95bc5ddead5d255384473a5fd49a9f2662da44eda219970ce41779207be8cb7fe560e58764c97c290973d828a88bc0fe385e49f6686313c0c08f0b34f96e33f9d1e7f1c4f3368bbde22d9a8e32c45815334601e25fb807e6ac36581140d727f5e20dd0aea1904d8649ba65f8375e8128a904349b1b90e8cebf7e5bd9f12d0f7dcfef5b235a5c1d00032bb4c59adb44460e0686e4df8238c23482a79a9b4363277cca35da69fa6402ca895f7db6ee99970c11af3eae5dac44d37db1e7c1de85ff65236c7b4c862c348ee90d615395070b5d8eaa7a65740f231d2c372b5217eeaeb1d6470e1fe80d294e2813dd1eaff6274f1c11ceaeff72cfb3532ed2d8ba6550336ffde9aeb3afebe9dcf3c9637787452d9e3a204ac11360b4e03ff21747128ded32957b96664f811816811e4f69a0729affb6f6fc33a363802695a1c797aa7f5d2a541c6820cb0f0e39bb730aeaa606e0080463e1e0ffa4198be95acdf339059f8eb7af41d5941585362e572134e88d72fa11f887786d087cb5810d1af4cef9b81b2f833751e37f35296e808db11aa4cd606261c145459442eb2d95aaf7bc9a714de89960bacce1d0111b395c98986770e3dcb94e9f4a921021949c50471fc32a4fee69baf905497f57d15f8cef8320bd1e705e600da52ce52cbe5c35fe2af240865e55e61fab125d9d32d464efff3db77d77b7e562b681c8c7f1471290b51d70690df4d230494b6d842f84692014dec694696c160e51563f8ed55e944c66539ca1ba26ccde28ad810a8253f2069c9dcfaf503c3e695a840950225cef9120910a12f372e40d3a7a7214367bf023543d8851808a2ca91d99c043d719ffda4ad15a29a1e7c366d8c4e6de71e9f42bdc0d14c222b66b0bb0da216a328fdcfc882b3c7d7fd8315a71eac5ce196ddc3dcd964c0d34d48292319e49aec56f73d6061772f5b3d19ae860ed6c917b0dea6b33f4300789270c3e91b536dcdd8c1eb535a7f04a4663fb4fa9a9adb9be003ccffc1783e14c3e9246d9722cb86e3ff3b5b5dce121bea2976dd00fe7755706d16a5d3528535b110df00f164a0d78ef48212658de5d68695a1d664801c0e6af5364cded3f91c59f99ea112fdef189c80fdbdc5602e705d4d281e2fb3b2ebe17ddca9680c5db8a607bf0c46f37c94e704f6a7d6a54dd64edad73e361fa06b8db16df635d36d8071a39a1ef89c05a3e371c6f96dde46ae2e1271a29f2320872e1716a07bbba6e57aa128285c55fc1319f81fc24e366e8a84ac5eac1f522d428f83ce32c7a6a2a24af1e82c81c495bfe9dd276e442812a57a20dfd2bcbc6bb31212225d711d387ce549c65bea70437fd83328a2b8bb7d9ce30bf6ff22107affc59f38fd75eae7b01cdaf796fe57558b94ab021aa1554fd25375bde74995f73fa3025139c05fe2b65ce771a4b01fafc4360ce50b34630e2362020341eead6c8d305ea1d19a3617d78f956e7030f501bb261efde0d5f95e0e5113313b1ac6a74cb465f2b8734c2ac5116eae7284b79b3f17693445333580fc03e16e1fa1d33c0456f1545c91bf6705079e8da2e73db3ba6723ec9679a3cee576c58ade2c88c1e8eaa587ceed4be97107b679e991d85541cf972900c47adf781829e2ef84824d9ab0441cfc6381b4587016cadbeb58c663820f147072b9f2a917af2d71a8fcb7e3e2f0c7617b51407c8d3ced1c57e30a1a3e0de2e64a6bffaaab104f7efd6383424b49e20f1d7d66260f697c4ec65718cd9e80e4381ee1cd7218b901f43238ad347f1be178b4ebddd349e7958f8c3e5bfd498e766d99ac1ae94c3dc0a0fa10d6a4d60ecd51a0ca418a3cb7143476a491fb3a2237cab4830a4563be156d0160f3ecff280d02a588d3d5ebf6758e273e632543e5591985c1cbb3c15764afd450f0877cff12440c948f2f773332762486fa9fc01164af1e2d6f063acc94c4f7566891efb3c87bdb931fb4ae45b4c2206a08f3613b2e7e46392db80806a97a7735e41946b82aafaaab66992fed21022c5631f39c206c084cd76f38b41f8e76b9c01a79d11c6a3c05b2a3aba3b28f833e85730ece5654e74c40abd037308f133bcdbc114c82eec4d1804cdbc82d809f362c55f14c67dcd09cff326de6b7fa3432551a90c9442d4aa7cd05d96ca778a4ce13f96530066c8a96fbd67b71a80f8eeb6904fcd4c37d72e632ce464619ccaf5e9adb1555b1605fbd28dcd06a18b6b489bf656ab78fd4debbbf6f4313eccd7f5e435c0028919054f07c10c9d648781b644ecb09b69604ab7146ee69c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3f0995092c595311f57504fc83d54c144a12bd005c56c3fce76f589f85869f20cde88964e263a395fe3dfc93cf1c6e2b51cb2a2579a98576728d4315a790be2186bb941ac777ce4bd8626ab633e11f207004a1c16ccfc84cd5c89f73f033f6e49968e0aab84f5a7ec87357aabb761e1db3d68e53e2f6397411e3247325915e8e906980e13716c34cbc4c64b89fbc2113d78221152f991ee8fea8b74a2b3de1354e878ad4a6e7d48da179c931f47c6a53c0a2039ceb89f106f88b3ed74a8ca70cb49ad8fbd09be54092a7d82e24a8a239d351692e47ae0b68c5d0973b16dc75394cd2d12635dbda1016ce64b31aaf67006b14d0d860154b0da41a204824af1b0cf8ea673f2bf68f7a20b2bdeb40d31b18a6f60f44d5b7af0aa9c868b920269c373dd29f521da3a5d6b2fa8b57e370b89c4d163f14b7752676639569709a3e28f9aa39ec600d3ba863d2ab63172c7f02b5cc02f28844eb9a4950186ad6f879f94d7656a3622bc0a9cb7478654f2551b1bc6176f34afbcccf4e04b750515e15ee6d8dd55fe5c3f8d326d1d9fbdcff7b8ccd08984957507bfd12ff36ab6a00f59c29ec9f8c77cf9df1887a5c8a54cf8f3e5737c6d9e522dfc52c0248db53bc3967ba3290ad1712b1936d46a8a1af9740898a043416fe9adb5fd615a101510b5a29872f5ccf9e789c0f17541da58ba6223bc7ae596ea326cec8adebad6483af287ff9e4417cc54133737f710055ec0af2c10f1cf516c4fac8d879549b04bade2cb7d64ad4bb05b538c436e446fdf304c38410e2ddf21b5f00c9dcbe8c741a742f69a403e5278d421d34d3e30f6c15ea1a3674eb082213e6942d8eb9dd0dd526c1f9e11068ccfd8b4e6ef575455e9d626c48df595cc59374cb49b6a0acfb297bb40130d384ece7ca8d3c59d8153989495ac985139ed0f85bd5b18a25db816ba72c63f6a01d37b6517376f011c4b23b7839e9b240617b11ddb16e1aafac6fd6ee7efc9c45c4fd11206c9a2529ae638e098fda5345f456c648ec5980303e1bf6fa1517ad0a88d03847eb8d81ca535215da5ef21454893131da831854ed8c9de97fb72890707e51eb2b56a1b3bf4383f4ab88f7b5d6fae7c71c95a9d76f02ecf1154eebba8514e089f3c8e592412dfe1389bff96340a8c122c98be9e991e5500b16898f30abf5060a8874ff8db9675798652494f5d5c1d67484722b4e84ea000ea9434d40b49db16dfafa9895a1a38ccc516f3a6b7216addbd09e1e9e99d0c1243f96e3804b04e1030226ea378adae5cc6f819f1ec6ed7552d241018ea4388a86f02da3ecceb31dcbfece23e5fb6c58d71a7b51bcff06c5efd53bd956eb9d811fa4b6c7bcf25a0a084e8e57473791a3d019b0607b0af8f887acd193d2844ebcbb96c18c0bdf8ed4c84904e9bb9e507d475745972e16c3261b8a1795a4f28ed7995ae7902fe8361e996729d62d582fb93b95c129538b1753c70d4721f432ce5bdab876d94ac46f3d60f744bb87c2d3c6f8e94673976b68e4d8917818bb4faef3a51367b997121c4c79c86a6350883aec36415282a9b495d2740f65badc9c8df701703e03e88e334a73e915094f2f64af3e484c4550cb841fe64698d7c3830914c10f369a79552d72b2aa5e163b1e7bc6fd99395d2da75617aa69aa7e24d26892768d9d28dc3d30645c99e9706474cb83af06a4df1f585a81205883b3c715afa7513833a9705b2c1228731affb262a8c2a9c10d949f94eb328052af4b9caf32ead19f2474047aba2635808bb0d0ee75c1e0b3ce4a94bd4544c594a2ef5f4f3a9569b4ec08a1df9771f1b9f58e1638ef6442173008c90307e6b87ca1c611cb621edcf217fe567c541ea34c0639a538d12a1e02ef38053317b3aa9c478f1ea483621c70a6d8f882464ed179e219852e6f806835fb1db4b225d0eec510745612c4afa1904daeb31f37c7034f3bf357207fa6dc63b25d1ffa939219183bb5ace601cd875ff3bb7811e7134697ccd52c0383a2a9aba37b7348c454eeaa863ca7f49cb2f06352a145cba42e85cb3ed9170003bd6585324c85d5b2e58c914b33933cd77a8598560b744b29dbceda09f073f57bb16de8b8bec797b31649964e510e221caa2fddc739b327d64ee52eaecf9d2100dfb5ff2562f7cc32b3104d2f1e5b091ad0df0d4217a2f6e6ebacdcb36f5012dec93e6b16fd1e89c8311b667ff492819e9f9660768b26d18dd2eb267a3b4989b835439efde9230adfa9506506e02275b92353038a2c72332508e2b494b77341ad4bc2111306549ab3ba8dce680381a198bb64f620421e24ede843e66f24d1a50792beffda00d88a71b5afd2ecbf1c271624fad485f40161bcb3bd513228172961389f3bc65580c21b6e25a14fea053998b38e29bdac70fd0de9b3c1bea8b5205f72c65c4f9c6688fc4a425f49ec2efdf40df004c9a7c47f222eb2e019c8305110757c6cbd2a8b6582269c6adc1dcfe79799fea1d41b505ffe77a033f1a4f87d388ae8896923fde49bb311f918eea28aae386156d53809ae8955633a8c09cb0c2a1696c570c4cf32eed1da36aeff968519e78738a006095ef1775069a1ee7d43cb6ebc9e528fb513f3b5f7db1e6cc734618d6dd7c35624a8025349d7776a8b08b872217a61ac13e83b603fbd42f02fdc2398ed41e1b242a44df1cdad2b37b3d248abf6092cfea3d63ddff8e10b56b365801d880a91f006b8d45900114e21ab14e236544f8ed4cf06b10c9b4c738507cb222b58ca82685019b59f4885f2a0abd5f5b982fdceaa005f95b943956286ddf183ccf10141da200606ac264142bae192c9cf71081231b527bfbffa426c7cc032ac8cb79d9d1f8b8f75cab4aebc9df7b7c4f849689c91ad77288756b1e88df4461c4773a09b4609;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdbcc7e0f2e18af9b82cae438dea29e501545fdcb38171a68b3855ad4a61969c4460ee6fe6d3fb87958568d33e2c85dd87929906eeaf12882c248e52552aab78b6caff78ec3c8ec188009733c1dfc2d2934f6c384c03c8c074db617151ffaf747417176d7c1bb45b1cfd2269662b631adde561c3db840a9caca3ab261a91203d631728727b685c28a96499b141026aaa7bc06eb07054782e98c5fbebfbbebec9a6dde4b30c44b19b7dc99147eb0f3a4db847d0146c54ff31d911e0b86dd9865b1b043fdb4d608f00e705aae1a4e39818c3ca1a954834ca289a07b913981f161da64d2a6effbd8ff4e3535b6ccadb5a5c38a25e0132838c266ad037564c45fc57d4fa890f68ecb716aab537fad7bcfd36b90f03b07a47fd6533172b1af8c1e0db893ef367ec5c1326dde216edef46308410d4c959fe65ea9ae321cd44f487a24cd56814abe1a57c2c941c6d09b6648a1895b889c7f880e7a2a3b9348de64d7525b2e45b0248847c406db82c8163f5143a8991d8b1c39fbf1558ae1e23bf15714d1b6d9bed3352618fc8950668ec052141eb91bb5276554f26061c95a27f66f1a692d3d9d7a8a73f6b27975bc4461a57ebae8564153fc336576858ca9c832cee77562a3ab7e838f73590af2455a894c7b275cb0ab29ce588b00c434138b7dbf564265eca4fd3de6ebeaae213e45af4bd139e54ca3d2b3cd5216c1785e468cc96e6a560bd4322c1823021a19a0bb4c30cc497f0a75197df520ed17be096e5744059c9cfb987d52bceb95f012b81a908c2b4b52c9f84758bca759c1f63113a941db9bd2de3d6cbfd12210be36204bb00912d4e0233a2f07726add75ed4cea3e020c1e9a80448bdedcb31fde7097b922140924831039b8975b965ecc230ea2c058b60f0c72d2af3f50b175fc39ef7d79182f79bd4e84cdf2946c1ff8161d2faadfcf952a93688217c55b96e654681205d1118c8f701ba09f7a0f89d65f70596fefe1db29fa73a9b5008ed85ed257b43aecc2d6bcb0d545c24704a29aee6bb78901b821d13dc895292ad8b59d96ae235cac96d0d7946236e6df0bf9731acd88e6bfc653da7167bcba41a482e2a72cc83df22bed44c4d27280380e003c20c101e3050944b67aa62f312b2e975ce8bc25248c517c5fceec7eead3166dbc55f3df41d7aaada012eb75ebe41d91473a48135ffb98fb4fe49a7d33d90e52eb6325507cd1a2667808c8c50ed9d0cacb80171f7ef0db0c189396303472081bfdca98e6f715c1f4d7870edb447807aab30fa01123fa7da2f32b118d27ced160e9f20824c4b765bc65d14fb44efb32b2c8e696cb335580bde79b2e7141d0d936fb821f1275a9bf41c8aecdbb376917b71faf548cf8fcb0e77a8711db32837d7d3f3e2d89aa55a9fa4b0e569bd77730508b596483e2166689180fd3fbb831d6ffb083f8d5f3b54db43216d48614c89cc2ec3aaddb319d33c946634d249c21827db42d048f3cfb819aafbc92ae986276d1766e28675840bf065707f10c4df64d96b1878b1502f6f00243ff3eda44b1260f3354d540d56dcdfeec627173f57c3799300125ff259049de5c37ac7e41ce33d25866f9c0d81fbddbbb41e7366f8ab6b2dead2153aa3076fa83b6ab121bae5842af4ffbcb70ec45305a14471c0b8339a945034d0e1e0ba0428e91e9b91d6300ff9b166167b75468ecad5e2197e6b6f87fb5f73f908a42d115e23e1f7e6e93a0ec708480884488e8b0b98ed98839c9402b810094685b82436f66ad5ae919421516facb9e2519ff7f5bd77abcfd8b9618bced8f43af922abfb4b200aa64df8ddfe48bd7723d83e8c06fef34cfb11ccdc8528ef1d8375712620526d9c95d1d8720ff2f903dbfaf5235320ed1f55b10c6adc481203d4edc81627d8a0ae3e05862939c3bb8297d72e05d8f8ee73f7136a79667459010cf48be445ede52a5b401ed4d80574d56b8b27f7594c12c97a28ea398968ee3c2f8e87c47d1e6b77110999fe9a1007d6a02d2d354f8ce42bdd528c992c09841376e13726154d5f7c96f207b808a7ee83f4d47d95d28b5924a431daa4f6893402ac5c497e47985c499f15fe01acafb6da9892ef8ee31957fce70eb0fd706d45160b81c0d4bf5205f188e4fb6ba7d8d976da02d673a8627028303590ed9d2384c8c501b5f20c4658c2ac1b4e56f128fcfa2d8bd549f41010031c6fe58f61a4e628fcb557a00956727c8045272bc5e2dc986db37ad8f5c6ba6c7f4fb2553385b13df39a5148fc3521c67b15fce257e6a1d6f9cdeb121f3440c9341d2789b22dae718cbdf6d55c3fd99ce24200db2b96e0da245791888eaa615e72e028f2d24e992c0592f76960027c279655545174d383f7ac01e4a8b2f07fd0553d6593b46f6ca3599e0fab6bc0e341fa453a13dbcbe95dc7becd1600250804e5bc5cc57a80282794f9544cbebb6fd0b95a247f1d85661f7bbd746bc335de6465c7f6ce00c557972ae6e82ce119952433284d3248930af31a54432d0c9380e28d610df4c930648f9706524c681466d700a85b2208f1a52da2b0fc6051c37bf6d7336bea65d0831fca7cada86c8b4c34d462083fd8b10633680969d62eff8502701b5238d141d547f31b166fc6fdcfd804420db279339fbc84ddb58c7cceb940283a1899d5a1bd830c8c4690a4d46a68c79ffbefe4ff8dfb7dbb398afdc8b583fd3d917b26fa20f7763bdb55d672485423fa84d7bdf692f65fb53d11a2f94e60770040ae71c5685d53791b747413175f31c0755f8c393f6401e9c3d325340e422583c8e881e1ceac1b76d9ac9113fac6756d43bd774fa70d9e2c0ee73124ce412e3098295bf1f3c9b1d169f6948222b25614bf54af6879b23d396e1483ac701373c0037e9d9b3507eea661b67ff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7002f571ce17ecf509d8bf409fa22ece476fd6747869bf223efb9079e2755faff629a3ff5b1fe1b27a9044269393c093a8b13b2ffd0f03a7dd2d7b23ac37602acd71a67f99be994e5ecf47f80e3a05f9da6128730289b8a2af7c7527aa83dfa905a93269286943f4da73d3669525951c65ffa389dd096b0c768b3be994b15e05013b74846d1fdb1b69cf6b3f1c29379805f56911874d268c9cff20c97ac2a085e62fc2ce2dab3b6d1c006af0f897ae224663937bb2f658693af027e68ff4d96f7b900aeab79c687aba64c7f302667ca0639192c54a8f97ba08dfc277e55722bec64809cf545f582cd4b56ffaa68e292b73e73b5fb49731243e5900da61e3605b740817473b1d86e69d8965adb0636a4181ed9993cb21a868f1877c3a8d6ab3868d45a734cca7be8d2878d4cd9f20850ede4c2959be7530c0217e468e18047d154278c4f6c7801cc121e7860748f81e6a5f62631ff43012b3e084b2c82c96c517823af4f345091109409ed0360a441c39d214cc4c0465160eeb292676b668256cbea6ee1076e565e51237e7649bc1a9983e1fa1eee6d8a69ddc5869e2c94f0422f188de76bfb47542e3452107a9279c30e4feeb9775d77099db45763db6dcc949ed05d7e09e212f68c8b6b8a06f3ec24953000ee8cb1f117d39ecf5402b3fd82e0e43a1880f614eb819c19ade5e632cc8f250c59b676ab7a5db36858c07608dbfee13a36aa2507622ba80f293e3c19bb072a08c13bbe8125ff1853a6e2a7d4b159ac86bb1b22424894fc91e10ed2cc811b99db6c4626cf4cef8d67c1ea1dba25df2dd4a4250e3987f48b8862c2d4b7432bb2fe0796eaf0388c61ad37b09a08f29f60b8e608f0c27a362a8c360aaa575d168c193ec7d6cfdc53bff486168645a9a21d380466222017df16b396711acc02b5ac2f53b9c180ae497e2f169bd64aec9b2ec333b17782df272ae551c5551416cbeb6de51ff00391eb2bbbe9cf91ee8017afcccf09914babb69a44aa202c6e15acaf0d9a8c5ae1ad708c4a0bd826e389e09934ee0ff675ee7968d0c3b8c69aa067941d7ee41dba550f793c0d330cbbd6b546f0d67f372929497b2a887c74b2b908b73605be79231cc25da8522ce27442d07a4bdf31160ed47fd9be0d7442abddb26d47c403b1e717ec5f04677a549042501f1fdef0206360b68d8db8680517ccbb4f326cacf83f88165fd0390691bc0fee785869678defba7012e22d9ea6367c23728e85c043bae35775e862c0ea5b29ad208d1dc037098626a3ded56dd1947eb9f24299372cbd8a6441608373cf792e190d8f4b41f90e7617499d696b7d5560a10433eb39eaa97222c234cbf0480cb85fc70e64daf892a8a23eae5ef61dbbe5977cc507ea9d123ae2daacd56e2cf0d4f5bbab00c2e90a1b886d8fa3e6243f8da19da76fe1f6b98083f9259e5da1bcbff86daf705ccf8fe4f198a7870a59ed1d3f078812e69463b3012651eb0221d1688883e8fbb54a86f46aa6e14271572c7d87bc09ff13497ac49d7e1cfab7762e66950d42871abe88757adc168262573eb07428c3272f016243f10c42f18ff7eb44e61c13d7f8130050ae4eef344148b646a565737f61f25e58d9fb864dc8d2bb8a6bd43872d2be6048b01168cc425c6d05306587ca7fa8b15462f68ad0610834881a1eb38e5bffd2ad033952ae0a7a9ca09c11d4893c7a025d68660f7e106f3df1cea6f39fb63c02908453537b78204cdce95588a895250af33c6befc72593e05b15afafa40ab86b16998562be9080091394baacb233c25c68047748b5bfe80226f896c2ca3395d2e6d45a79bb38559eb432d0f4f3a000d2b5b26ac183e09a200e64009fca2252ea734d09aaa05981cfe9e74bacda8931847b37de9c8f4705b81811aa3251c93a1a90e583c91b23b7dd4b4bb85f459762493504937ed91d659dd5747e888a767aa05b22a0eb0eb11a97e172c8ee84bb1092b8c7808219dd3ffa30921e27833de164acf4efaabf859b937b06b6b68f0b051ebef1cf9c54178298b8bb41fb7879f972f9ed6899986069e4c07d97f8628b6d2167a18a1e3bd703c12c6be63388266c2182e040abed9600199cf27a29c0a4759c915f4aea7fa17b795754d12fd300d1bb7acdd1ac0b4122e42abaa7515e6d54cc279c3b382f93343e2f2ee2bc81f14eda083576562efdcbd31a7471ba8e576907382213bea16737fd6de2cbdd3dfd58e294ef33e5cf5e41c3af1be43de28fa4bd65c2281d041e513eb14ae909d942ecfd1bbd5ea34ddf3018cbaa9c4507d6b2f8776723c0f396174ca0c220dba3385faef7ee535ccac4b5e34bdf865298e87eac82c9ea6b1ef2dbd5cc97e75e46795193858d6c345c9fca2622bf6557e165101d693683758a2d8a4e7f3ee982bc75bcdb992e05a0997ce04dd8f1b5884ce359d23f78cdd028c2deb7e4d1d728d772120865be5143d5e72956c50156be68615566bdef5fcb463afb0b87e68fd711dc0524dc531c09c715aa714dbb1efa24b7185130fe4c2476c9b2339faa0f664bc5ff0bbf96641a1194f4c6cc7aeaab9b353c8db1a51b94701fe9c66f42ffe82b072486e8d987f07a48178b8c99cd40581b58f728a0c5d82d597a5c63f58c0bfb4f8bd722c53a99b196126b4f1544b8e542b919ba6c3df00bb44621992bfb65258a9a74f7e056a11165240b2049e81df78a0d509348d7ef7169e548fef5a77cfe9610dc158b98b22d3e2fa190e1606775eabedfde0bb209c650c35f45d3ffcc8d0cfae60dccb965e01d33f5aad14c9e4a5867246650837f0414b2ff0a1f856871f63356276c5e43c09538a59477f9b05821ae0e1f67d4974dc759397e08d0eb33a54aa920948ce492d259983c97cfab51479e46da0c6f7e15da4b185db;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h9498d5229b3d81bc3bb7ec5b8aee6bb559eb39ffbfefa5a593708e4f61a14254f3be0b0656e0f88fe5d440f8b11669f17ffed6a7651c709bfdfb7eeb74af6481ad9f77a36b1c2af4e9ed78944b342aa64bf33c398d54432e4466c6fdc059577f9fd31e17066b1faac7750532498260f4a031227de4bd94e6356370de6fe8b8cc7e5e629326e09318f19305d5d6bcf37125ae368929428ea234b75e31b76b59f4d91c2b68b6c25d878f9dff637d935a77992bb68e69fe6e1a3a78c8dd8da40779cd8b73ca2a4c8c69e6ca68276ed4e2273e47017affc834d6e2ad61cb8d05d937ad08f5a24f65ff11805aa0800310607ffa514d183c3ee01532de280e40616309330585642b0673ff6986e1093a0ddf0f9b3abfc9014016bce44ab087835c691b703b37ac21941eb666ad0b324740b7e763638317ec6eb07db36a61a188192e8390f3112168486c7a90a00e5e9c7f6770ab9ea8d592fef47340731ca7e9e8bce8b500589da0bc843620745f3e3f6c2f524e2b164f7256f3ecb8d97b0c69876c449913199749dad836b91b8f40b87bbf39389a057ccf86e4306c9d5e12422cf2891af48c76c423b14e3adecbe7742ad4d43976a03e957d1c361be8ae914fbb049210ba3201a3445585b0976a6bd14e009de82c12211c0ae9fdd9c5a874e233cd47f8acabb52b666266be3c56e6b08e6b3ee9bd196b9c623589a7a8ab001653f1fa93d1d68e6246afe109ee255a6447d9e3f1caef748e955bce0ba13624d1b6a9506e9c68e6d1075101f8a38dce6ec682f2a7032cace1b6d99b07f95d53c61a9adb840e58f8ccd364705e7117a63a0139e3df1f56011a4fc7ce3870ad84aab0b0c20a57f48d1c1cba0e0f3a4a1ab4d87db2dce012861aa54d24277e4fc2853c1a95b2a2cbf7428b257601cf83fb02a6bc50eb00b6630848df27361f5a94910082090c0a386b83cc0998877d2fb86b4be8c5eb77076e4b98a8bfaa4d4416e90c17affac9bc26614cf5994d13bf5798b1b771088cd18ec1ddeef7f68ec271f7fa98a25cf60c9b372859c9f627ed3beb1ff6020b34202bd1a610bd2e8ed3db6d4f60eef3a77d6b1cd0909e690cb32fd6ad1cfff5b824c6ac0baacaed90d42d510839a7d56c5925950b2970414083b537c2d708b5e6a714626f4b61624fd7a995cfea45af01665d9986d1a7005f48e99db6a38cb9fbb870bd8b4c77c71356145c84a6616231ae7bbfc601f3ca2a69f5a70916bc5fbfcda7922db91d1115ce663f6d4948fb0518b67a9a97b369043f0de71b50b45216fc0939b0c7835acce3cdd6ac8b612cbb8c33846d5bd5c04d423b3cb1fcd148e70e3e43c669399dbc9c6b89dad9b03fabaf9e102f8d90af72edc05d2bb727094898db463fa69773ecf30245dd7d6bb20b1810ae7ab8e7128674da59d75818a135f63857c4b2162a0da95e50383547a057a8f1c1785c0060662d0c84f555ec1860a424a75f6315dda1d31c819255071c75645febeea23ec6eee14439847f701f28411d3cd7a789331d53e4403d9daef9256cd95e90b5406b5f6a088499e741b5915e5627cd90ff5afd6bdeb167cd6c6826630d4c8bae0e7673899bccf2569d72c3d4b047892bfd14a778849b66e9076b1d86887197e86b1a0396372ab446918a7021011891a5ab69d0b807e59898c4886cc98baa0d939c9a3c179db84875f64aaffc73e7cfac286eb195cdd5135e475a7d1c7781123129ec8271ffd0dd9271c799eb62e318838e71641b124eb5afeaec9176492fa47298623447427e4a39655491bea6d057ecf2272ced44abe759edff5a47cea219cf4f6721c93814ab61bcd2b6c0df40bd0b20dd1748ee7efa183cd7d95988a58441661e477863e76927a670205d12af634cf331c9d3641e8a49414c92d06012ae6ec26358b4f746d336a6b1f5303928ee6b5a28368a55bf2ea84db9b77184638640002574ced5c2f63073621d1e9fa218192eb75f1bc8f0ff96e3b0f7de93666b0ee1fe0966e16135042c5d8a1949a067c299de832fe67707084467899b5ec77c629555b7ad74effc26a0c0d5b28bbb3923908d363f49eafae75f6ff8cfe492bc604698e6e344b7d08a065570c0e4775faf3d0dccfba1329b83a040078006b96a9f5a298bf8fc6ce89d3f8c4130deb1b25e62f6009c7b3affcc1644951aeaeaae5c76fdd68d19e2a3c35706a405e57bae9241fb599db9ed2a968b9d153f9d827d72a494525689c1eda38fd8fd1edc8ec4de914f92a2d02870ba19f64d676ed2b6f3d9f3aff1254749fe5f5d424e6cb99abe42158c8f87e612796077cce762623360cf7f04566fce574e5dc2441fcb5fa89f9e00b027be25704cb1262a846f8827731bcdd24f56bbbb381030b4899e9b24835c00714db4f9c15d6c1c6281b7c773dcba11633dae253b83d77bf6b3f984652c4a559be25aaaed0e61bbc48d9ed59713b25458abed7477e90aa63a54267140ba9b21c3c54504f666dec0974633758f318687138461464aeaef1079df92232c8de47669481b3000b19967aa3939d51e63eefe7be0bef0b8901ea5782b40667f15401198d2670c05e51311f3cd2fc4000522482f2aa4eda7369a7c5b81f8271997497b752245a4dda54d9f1dde717b4b8c6210b0d8c4c7571ee754052ae13c4bc1eb3f6d14dafbd6e9df61019f7eb31ea7e21e3601e53312e4a966660060d81bab3d5fc2e160f9cdea5db029c53d574753f7173d9da8821217ea98db88057004335014611486d63c49d76e1ec0628c3720413f64861b0233efaf4a3eb34fcf475c5d924e623eebfeae18e458babaefee52ec3e7c6462eed64026ccc36e45f6d7f1e064fb6185cbe162986534f64c1282cd90ebe33017a907b6698d098e6728234e7725ae4b9c1580f1fd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5930f472566853052c97d9f517ad6650d774581e7be8fcc3f6549c6224201e482a3789eb1fef5c19948cbeeb22e58e5496b6075556e213968dbf9de7d15ca22602b84cf6089416b1d7a80e9772803df1025b7c55cb0c60912b0c00a391d64e97f7b9d4b4f7bbd9525586c920d7a6cbdfe146fd8080c8400effb38a36586344f02c9bd9f77ccc0faeda95ab8bb37534f6508a4f03abd8f920974cec74a5ba3b27ed5522054346b4526574e27816f80d4aaf462ab991faa1366bf29f28596e6d32da3434314785bad17334ee1087bad98ebe4bfd4f4410bd69ee32224c1ebd54658b75848e0ab4107a9541bee606b973779c318f7c3ee6f663aaf52c6a91f635003c9b11daf2b46b049ac8aa515a1ec4360f1c1b8c088522d945f91b52558af99c5761cb5135f8c7d30d1ca1df4d99a3a8189923171ff6ccb5eeb490e532d924fa5c093148c7b9d97797e4bbb78cfb9fb53dd030be085b69cd5a4e5caa274268db2a84e9d692bd784fdd72e30237e795f772c5964b95bcbfad6a5e6d1291aaecc6dc1eb2fb7b73107a2dd5d16cba32ad2801bf8ef3d8f53514cdf6ebf09d71600531a6f9835fee5de476a2e49af072219654c3650295bdf07d411f13de90c6528ffbecfb23ff7601b26534e8c69e81e543a141cf2a27c23cb7159971238e0ac8fb7f89b314c37c9fbba5ce7cb2b89b428cff18b4b3c4383502b7840d1107db1e29d3db5b2883a61e7e520bf07cc0242d0e1b51a55a2ef75e5e25379f54a95cc0bfb5e2f81fd746abf2186b8cf24d2e3f0d0f22be21d6d5eb54cf74ca5414a95fb5776110af4e7eebe2a4f904d98ada90f0f216432800b58cfbe9d1a8144ce900bd7163f465e9dc8b88806f44235dfd471e6d9aca5016dd7b7813067553bd0ff1c6bc4fe78e05782d31b2ccfd681183c6f8740811444a43ea527c1da6debc37e0ad55fe790f7411745dccb5ae967bc3caa57c1d0348f30bf0b085455fd74417cb39227ab4200576fc612b0bba5dab3b1c5bf5d4e36824a6e05b2e461f1eed62127f8ab5927889cbe2893d193c0e966ed539d3474e9e7fa29e3754e98a0e9587ea168f127d3dcdb581b215c05e2c9f6d3425e3c5f144978b0c9c2fd6c4a0cb863e7249270f0423ea923d572fcc1f89d39da67cfe3cfc73decf3012d03f867aca40a2463cbbc3b51375267813c45ddd25ad9aad22a1994cd685bcf06412966a4d4c8faca2b7d3d215e7855252b08679da1c81b38dd07dd4b0b292819d386d6b664341ad5be96f8a0a01b303fb2e36983692e7d55016462b8872828634882e9d989de66899d6694efe692152ac1e95406e3a0ee8d06f762cdaca40574f767fd013688f112836fe12fae569c6c77e2052d92cf3798a9e4ea17ab3dc5a38a47a788494d56bc1c1a90dfc0e4b9a063bfdc1c47b155999f7bd62665795b19505fad6a58cc8593aeb1cadc65c2baaec471338a14b1527ccdfa7b02fc8f979d36c24b2b7e9eef9debc1978ac7618d3e727760f8a686660eacb721a710c8b8628706b82a65f0655fadad3cd533b15404bf4974364df5e0585e95cf0962439456546906e7be84607e145f471a12f60f89a385e6261aadd503f60c3659a8910f4245ad3a6eeef3e3c2edbc02c271ec72f216c6a923ac8dba0a99e13e32de2441366bd01d67e19c684ff1f6f1c3b2dd6d7682691ac1118f86a37bd003a142e1451848acf5435672bb80e0c486eceb2cac7406168c42e6eb995f91ef6813f7c24578ea24f12bd819edc7653e0322029f8cb87a141752afaa7b029eda5a81725d6d652796b3dd4cd64b7de2aecba9559ec386302eebc4ca4611691e392961fd4a547e050a69b8de679e63ffcf1aad36e77483f92c308230241fc5e7afd6f397ca57ab68705ab976790a55a4b86fb543a8bfd2c739b218095942bac04bf792fdddc90db67ee4bc29d65c11768cf664b478f687926367b6383008f6a944cc647f9f98431df62aedb58334c83e45ce76b2644d7c25ef55cc80557ad4833588345123065bc4b335e85caf0fb46ce6034683224bf85b509fba0429c547631f7fa5aaed86d3e611d165e917620913eaebab8104b9bd9a416a0f8d6d808f08207a239c6966fa7c732dbf0ca9e648eba0c17b47dd72308a769e9209950ce3938d546443f968060f9972c5b337739ccac910f5beddbf777c9aa937822e621347cb6cc7e7b575d54a45ccd22d743745c1b23acd54de123c98c181c64b3556f78a2357ec57a3f7db2ef7a9245c4f08036b439551f3a82ebb1c514ce906949ea9b82e2c14ce71347567b2f4ae7cfb97fa4c0a0d25096a8dea7445391af570cc3b28f4599fcca0827a2a904fde8091d56e00bb91d92aeb15e019d7d7841975d6627e576e925ddebff7a97233d526c377cbb39a0795d5cf80087ce545031ee3c807107cf279d9b0ab7ebcf41ad03dedde959546c23227a2044006869f15482dafe84d903a70a88857fa54caa5f15539e5ef4b458a2b1537a028b0f458a9e92286e9f2f0ac509f19b737f9b5dc4846b5839e6ce01f9175ce7df63df5369153d2f1cbb216dae44a777934d3ed2452527fa5efdf7c73cafe5f093a5cd3ad66db7c7226fb4760b445729442ee94e300deb17be3bd0fd2147354755671aebe877ac2d0e79ef31c5ab58c48d4df2ce5978075c234f078b59b14661cc9965f87dade3d2402b674053dccdca9bea7d6b21f54207a25e594103a8b3929fc462a9fa2e6c00f5ad5822ebc4750fb3b90b82a23bde67875a8266703d97b2943a8b5f2ad3d43cf679bb5c68cf18c313632ce34907be96537054e4d5133a2c892b745f4f1ef09e00a2bd4eb3c8d31b0e3347ec5074d9af09fee74a46dac5332cd955ab669a52df882c6b713c1e3790df805a36411a709b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4d6e35ecfbe822449c74517f13acac85dd5324b24fcba69b938f54c7249d0bcab6d632a345cabaca619d35dc162d92c402dce3dc89158ba6b11551334b1df369cd80f3efa8f9f25e5e1ee1371831d06c9a9e260298b096b497268349225e984e603ea3d5dad0cbca10e77a27a190dfe055a9030b932803b49ab3b8011706188c776bb9b656e8122909d1eae909361f762b996d9bef1c9d01d2ce07c102b3bf2ff247ed12a09027adfffae87880583e5847834a9a66a562bca7d777cc76dddfa5e6dc716b6e9d8d28a3a172726cdfbed14198821717d3ed5daabdf47259c606d5e8790d7b1bbe4076e3d9833580c006d7fae0fc347bff6eceeaf22e904c261620fb0584996aa10df452b94407cd429bc3e6a6512d1766dcaf6476ae778a7ce2f3732d4d7c896224fe008a4e4344dab647c71e7245bd80f8f34ed249b840ba83cb138600ca54b08840dcfadb06cf7d20dc3001de0acf7752dd6a320451ede085511153de156eeda3db5ada9fe9ac66b70bf0136545bf83e43a2b613915d4d138e2f7506b263fb5a9b648f9cf9f5e0ce1b3a802a3c5d33acf23ee21f4b9c7d6732b90947f81a067ddf036e0a8a269e822506147c48d65c4811f2c7f39cc35098dfcf6ff848663db68361d7652feec6943705082de605436410e1534604df7ad5d975c3f1369a83824f9725ddb6a6c280f4659b4caee6a433e125b8addb167e86aba77e73edc214747a1a6b436118f39f2b2ae1bdff481d8820296964135fb483047dd26113d9957bec15cd754897d3d99baedfc8186635e93a398cf87288fb237cbb19146450a4f4fbfbb51993a94656ba7726444d2f66539e6c726e190beb8833ca2d897c27fd14c31324753cecf6a5d1ef52593d92e4be8ddd5bb4cc5f37c3e94cf4d4ab773463c01eea382c26b275c70303347ec7eca7ab3497c099b7cc2ac9f7acb5b0605fd2504a573705129ebbb5232c0e1218a927826ed988284efd63445cc6548690853ad9d336509527ca2718b7685f4bcca3df5bea23bb052656f2422fb5f9c026f9dda47bb9167034d22f94e98108d580e175d99300d04185f0882fb02416da81df12e2e6fe6058e15f2f185b470110b74ca3c19ca4f1b20980a7b2cee3f290429822b7b27a6b76aa372949b25ef0bc4a59b04154ba1677f37afc2397ac1c56226c5c87dcbb228f9a4285b8a222161c263f46d9681f250b40d236d06b8c2921bab523d6be20257aa41d35fc6634bcd3a000cf9478d56004660687e431ecd37f4c5f114edd92017d99d45c46a6d661138dd8e57ed875b7a0685910a878ad36e6cdccc3d6345a578e75284559c3461af5c8d0ee503c7b0a811971c6945ddba0058a1ae6de76a00f828f9e107c6c5fb3331bd83cef6bf9a36440ec919a19af1f967f3d72a323642ba31888ea3fc21eb6d39a6f744d0a45e6c0b2b9934bacdebc6ee9337699d6476f360afc3b318205c724235a9cbc511398d425886be6f840f1a2f38e99e9758be5a472010ddfe9c1a35c5317bd7cfae6ce5a3f3b70cc24353fbb1e5ef4259a8c046853824cfd54e1ebe43ec118090c0a76f7118357d186609e12e6165046e95b22c605fe67d796327d1808bb0b317ccced538d56ba0820ebbacf59daf8ca010ca2eeb5953e786e18a1a69f5c4cb4e644e821e28eebf3058565169e5241124d64e088f9878a9673a97a01950d5977e257487d8bc92a502a97fad1d1e25042b84aea7e148dd9486a2942fb2ef5a319b79eac1d6d2f69e19a8bcbf506bcfadb4fa759cc2968038422357677595da53cf3450cda5750bdde9202bbdf04861b5bdee70db20457e16b48146ad02965b695823c89f3a48a542805b79e1d39da16c3859a2cafbe1cd7550adcba5dc84e803d4f3d2ad5e281d551ba95b7bcabafec7a394935e8c4decf38edd51da118c7fbbe03d6fdfa06d52a339f66ade25bb47cb91cbe4a3fc5ff8dac0bbe65d4e587a06042a27d343cd3a321bec7cfa9e3f2d6bf0e5efa249e0e9c3c9f52b0976c882cc8fc80e131d7fce08094330ca93abfa0778b4b0dbb11ab091eb7d0affac7b8e11fa09cccf1c35e73177edafccad915721639b1a5467aca3454fc527d8955aa55e2718c5f2eba0a7fbff25af1783e16243621bfcb1dde432fe1921fd1c92e8d6e894ed724d41c0a083f682259704f6e1a8fe138473286661104ca179abd070cd8bcf2e832c30741870adaf2b68c8d691f73efb99510e1cde6c6e014ca9c4d90519033a3366204109e2efa99b9886bbb9c923d5f66f76aa8cc3f7b22a344865a266462ed74b38b1eacb7f928fa0f8c1c48ab8ef353f7a2de554092bab3c6faf68e915d3817f8a0efcd18611b56bc67d9f85fa9d26a6787fd0141baab2b36d4faef930efb432a144fc297476337ffe561e14b9c757fa0e41fee56bf97f64d567bf5d1bda66c4668f2355ee7e9f1862b2ecf03be3ddf1454917f2283b0b8a462481747875fd7152097805a607bc6dbd16c78be27ddcc1280af81ef39c4f2128ebe0eaed32dd24ede75ac811331a90afcb914b829c2b5f6f56040112a8b5d4461f292333c03511d0dbd62efcb6517ee0a41db5b4dcdbb8de7b1a87f2daaa3e70a6ccccf899b938549e5713c5e6be904aaad88d00ff858f5731460899b4e5457ebbfc6ae9123c0237bd0eac870df6d299b97c3b7870dc525d723aff7be4b3b503eee22d48aef5f87da733b9fbb2afb7b5c89d5dce31c2bec2d73d3cbbed07f16815d98187df2b7c59a5a8aa4fc8016715443df4deaf33a5c7809534ed5463e304f8979f534e0b23ac0b4bda4d6ec7d5ac652e261eb659fe33f130fa2edacf3ca8f5763819cbb5f03e724876ad4c3e72ce52496d77b59862573693cccca483b29b460ec3dc1aa1ea427b9b2d5a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha9aff31238d3be3865bbc2c265d2f75a187f179c1095b961a23d1d97ce5aeca70733fd330c3c7deda8daae07707f2622b586b1d42e7894ee562dadbd6be822990ed9b13dd47020e0dabb48344a8b039b8dd0b9c48f4ff7d1f51c20bc0c153991efbe56b71326370960df4c1c649e00aca4649de421584cfbe24570ccdb0779adeac1f247a6d742b83a884bb90b672914bc082d11d3705e8d974f7dbbafd199669a732a4242220921a53e0c7d81d29816c1cf883567c2fcaee8fd71db7403c250877992557f3f35970efa0e90adc653992bc739a78a92486859bbf253fe0a66ffc8d824d8c663bb88f9ca77b87afb5ff84b014db566b3edf88dad3886630adfdc56540b8421864f697a7faa41a9841f228c0568ba13425de55a2849b437ba08035ad062b7af677555a9e466f74e7622cf9ce7bafe77246a823664be6154b41bdde4cb00347e271efbb1a47b4819668ea99597b5df817f70905cef3c8df7fb47fc4123bfc3c7fcafac9fa01ab73a3009998d020366f3dc1d0bad0d1b97fc4898696335a9b2f0751b1e7b91dbb388a73d4edccccf09ca6c22327ff18745f92bfb17ce068fe188f4abd68d7dfa4e38eca0fe0a1751d6e2522002c397b99ef0acc568aaee711189d5febe3a6e4e70bcab8624d6cd6c3f8b218f687ad1181f4e45b07842fe9fc3547d8fb9787559f9ea3c29a77023ab1afc2d4b094a9297fffe0cd066f9cc097602bbdc468d999b03a4f4ec05b6944259445607e3b6065b1085199d276a036b890e133479a80e34faf2ac220e31b1155f13c7e3060f390f531a4b42e62bf671ef2ade2afbbc385155fa6357aabe8280229b9ac144adb9aa02461f581f96392a7192ae41f6237ffc069f13dc58b3e08200150537139593a42663dea9d0ad52643b298734d3b1600959a85b9f9d884e6ca1d1a355356435e4c147207ac0ca96176116f5283a218bd0c5a2fb058a7991d2671cf8ccfb35e1319a46171bf3760416f48bac51451156edc6c90ba489f85a6ea33ff461f11292d27f94ae52ad83bd383525d36bc2fe3d7737bb4934e94dae2fc9ec9cf0a6efd72f6ac9b75fc8ffffe21cbc9ff66d7de9517f48ff604904c04d6e45bf3f37f6e0746f394de1457932420ff7f26a37383c170296ef5957cfb39d13b227979f0be783dbd721fe4f6c175f28b50dcd79c3e53cd775dea80abe8e2a94b0fb37975b3b40e5e84459d36c64fa9712d4c4193597efa9c2dd8852bf82a72d0a0d8c4ebbcbda905791d4627a140c3f22302cf7d8e27b98e28a8d2e6faa1c11fdb1d68d37b6882b48fe7c92932b412f2a5f58d91ffae5577e13ac5263fa7ced068d357b5a10878d033d979c77948a1b22d7cd3cdb9bac3960a008e67ef81e2d3757436b8e6dc337bc1b437f622ee3c0fe697754816aca7f522cad8dcb0a41f23578e03402362c93fc2a954efae1ad9e22dfe7cc9df345ab5d8b8624292022358439094157129cf88952a78609b94d450c5310a61fd2f3f7a2fc52b4e29b00e577de3e12c7bec7374fc15324807009371d7c89f5121edcd6cf7906dad0d580015f89430170e5c3a2992c453ef97f95cbba7cbfe71f43c6ee6b69709bd26111533c1d565830234deedcc5cbea3f2dbee90b22e5b1941cba768ea1bf75e2897978874009ab3b27a71f34106f27a2bac0d0435b8795f2fe02366d1482d676e003830ce420a86ac49af4005acef1a76817072dc57e6c0ac3dba296e66f0c02a474657031fb2d89df5963c27bc1ac76e39c98be2b48309081a84925b3b9a0cde3e0552e91b4b58e5e8049d99c2b701d71a4216e9cd3abb1306fd318449d6679392131874f45079920c9aa45e506f644837899462e5c570c9125946df2bdee4a606af3fb3b9257f33100f2e3378295f36f1116cf1c7fc3d36f6fde98244985fa402647c3ae4ba88d010aa79bb2c78797b01a2d3a47d45e94ea149e4e397eca0a7100bbc2fde99d7660598b1f56043da560c0c023f3d9f3506aee27de6be256cbabf01837ff5cc6b8e99e37efd43f49be2ccb1161b945d1da6b4f87788f03643d0e31099854ef2740cb0e66e53e4255cfa7c8d034bfae94fb5f849f66dcc33984ee714937586bd5255580d611665803fd80f3a5d61bc839c5c9e504f21c2ea64343261a4bca527ddcfa88807c5048cc31c25d867b2e421949ba91fbc141ffa5a7283b530d5a821eee306a3d5764be4d8ae765c08f6d71347961113e5e66baadb77cb3ec03d4c26eecd6bdecbe075286ecad3980da6357a93165b3b844ed39d95584d4249a0ef78a339eff59dbffa0659b9e12cc6e9831291e795fd6ecc8efd3eb1030c8f3e5f0f212ef484f529c8cebd020c963cb2093281c9933412eb6fa48b93128412aeb9ad96e78383f0dad134045cfbc04072d03d44177f5f58fc36a6a59a4d4a67be5318578ef388a8b00709a20476b3e5aa53502f9896fa29f41a58d792d30a1dbf36ea70fec5c1b736343897967cad7299df3fdad4da1061182f62a016e948886461c980b5de66b959edf6716febda1e465b53d94105ddc0430553f128f1c7aba41a3eb4b37ea87e3c73901398c1f2b504ba08ad9317eb7998f9fce57d4ffe05e11261271c2b8d37cb2774001255f21247076548527f72e5edb1d1b110ff25f3b477f39c0d52582437ff4b38fd1f79c1bced1a3270749f574edd6f756e0eb0d165c2888206d24f060b38b6d9fd720ff1fea8031f544bd7a8a74b945ea4205e1be00d6f2b464e9d70407ea938dd3aecce91592b280fdc800811101a5143dfe3c413edf039cc22dbfbd241322665f0502e80fa6df71a371018ce2f989d76ca388e8c09cb36a296d9130309290267ea176fcf605538a64249ba13b0903c2d60d85581726eb8bfd8a29f63a5b7b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha4da44002264f6feb3486f54b172df73639c5c1df2a8af69507507b06cbf46d366cf0c5dc6578531e385635a0f8650525d84fcf18e3cabc8061996fcbb9bc03f14a9c42313a37fe7463e7dcca4dd026046e3d41b54111a8227ec9b210a17a6a5f6272fbeba651f972cc3c9d8bf032300570d25e7dcf9475778f3ecb4a6b77ee550980bfbb50c02cb5936fd4c0d8392c6236fcbc73f1d0df5b48d1a82fe2387b9b79141dbcbd38b44393d8de757d9aa3fc8776b9b3dec3b6823cf740d705235caf9b6f79c5ac9b31dd9f7fcb466a0573ebe67ab87360303781102730001a4566d3466fa5099e40070cfe9cdf1bfe99710b8731e0ecd39b11da9b8ddc28f268f7d30351e290fdefcad45dccf04bf6f929139719d3a9a02b802495b37f55ee75a96395d2f44c822b910a3ab0f1dcbc1cdefea4fb4bf0499451bec5c9490bb6142d42bc9798f73615d427ffab2e9558a66599fcbb7c8da699f9ad6b06a14132d9861d8037200cca753ab33c4487870dc0a0b9327e8bc558f48165a321f1a8d89b46488c6cc2d896806d1e55921b53765526f6b33c156ac2fab7e6d7f178ed162824d58803dafd9b919c82549aee02df67a4099ccb289b23c3bcdfcf96ff0dbc55f47cf01a1e6a28b90f9c5204b318e7d83a0bce65184c37fae76aa95c8269c9a590edd9fdb55aa10628bc7f55d8eea6fcc67609edb70838262c4c6e0ea4d64f70b5e93cfefefafb01948e77c5312d786c821cbf9a16045caa300b468b3779873c33030d748c9f8f1aaa22bab48d0cf6c3869c1481e3ddf1a2618200999c36ee5b37a2b965a80b314fecd12c6c74c71155b4b378e17229fffd0640272bfbe91adde3f983fc7d6b2f626963e7eaf01f190f91b10cf9a1e57b81cb223f89d8dc99ddcac7a386f6c4c6fd03cec313655cbbf4bfaddea60315898cbf8f933f894791eb39100c6b71d2876cc1d97888d8d2a86c2665b73c6ff8d79073e73cc8cabaf4af4cd0cc8f1f0cab0ee4c5d1514332e176044821ccbbdea10679281590d15be040b50e3debc0d712a9ac25c7650cf5919b6db5b4876566ef2869ff6c1d6cddc6aaf0e8f65939cac74ce250498efb5441c0ddf9bc6345d5d02947eff50d5fae9d3eac77ecf1dc07c645c7740cf2976bc31415788ab0a8a32276071a47b989cdce6f0765f15c140521688f5c007522116ebb59f54a7ab1718993c994b5a17885e2e45063ffb7cabe59353dcea0b391f33bcdec1d73d83541dc8a5efb1a385c1affffeddddf6737c0902d8315278974eaceffe706a58e8902f4ad8482eca063898c48f373c89dcafb4a7260b123de7a3e25073a6bde2c721bd5d6e525d7c75761a9737c7592adf9952ec1cc818dd526f24832b0d72219c7c43c106716b02e7e3c31c10165cc8e361d989ee46e7c9ab29249824197bdbc9889cdde8528bafe895e03bce5f891381764375020c641e353d39b447f7482b57f1601b8a0e74f258f5eb35f23c2ff2f1d7161e0567a1b15e454c6ce692897a5b2276d99168d094194bf1cb5e919ee28b6580b6e2e63f94ab925f974e3594dfb1cb9b0267372c9df6685ac7e06ff5717ce8bd548685a0676eba657761f2b8f1a8f8218440c15cf878d711f204b4a3cb713b441220693a499684112865d61e85b50952c9b23b6a4722c5cf0c90aca7476cf6df54e225cc0e482ab9c070ced10330523903915a81cd43b7127702ed33fc3c56d471ac4a15a299ade250112f439e7ba6fadf259148a8087d1cabc41b0154d8a7da8f5ab48eebe975d804032ab87efc96149f5f4f4a4aaac22a22ab3bf7c432bb93bb328ec2e2eafc4442a2547d3c4a8ebb44682d7797beced98a626f627dbf14af729d1f2fbd786e5c4a6a0198fb48f9eb328c39729d24cc7d199e93d151e624c124e0e8ff5f550eae838e7e5795f9b494c1afdd64ae42a01daae24e75346d6b62a4a5177bcf192241021a5853d462ecaed1ac758d0eb85188644d13b2c117b63bd9c3cacf125a82a7681f4b7bcd4677987cafe4c8eab837866cbfe314745bc191ef2b5668a8a0902be89750b47a33fc6f5e548814ac4e3772c1bbc424f8d0aa7d18fb1fd42bb3fcdfd5a156703d5f6ce148aef57d0b0678951d4e64d9db58ced6f5a3e111ea5bc9a986176fdc8b0b608ee04c731545257795cee19f7513dc9457672c4ba94c596361f4f3ba71aa4a2728ccae76faccfd3aca4b3db13db2dc7974ebd9b118aa194dc9e22e596d7a44ed7937d3a1710315720bb8aa9b8158541fc503b6740e0b05f280a7ded1358c3b2ee9e3a91f64b5a859602cc0c9cfd86087a7ee059cd76decbe489a37b7cbfd78ef214bf376c44c2aefab9d5567d6a975c9657004b54fa30b3de336f9ea358296ebd10bd0ff3efbcca8ff51857186ce8a9786b415acd174aa7754b7efd4cb3a10f0f389587eb25f48d84ed9c5628df073abe72b089ea2905423bcefddd15887e11a7f8ad13cc8093268ef4ae1e3545bca9b5791f2c54c24c6ee9029582e5b976313da6318d0390c8f83b7d6f17f25e5dc2dee4e4386b47bff7990be26f8c7a0f7fc4864566fe3ed1ffb19f3edf10e7b86c21a8d128289d9c61177fdd6083001da1ed0504dd160a8afbf9d26bec2d3c5471f0a1dc87ddd9ba2152456c60f77ff6c78cef4a26092938fceac242eea517d9938be84da32fc67db14d9853b742a56fdef4e0402de8aac39c206feda46084932142a751a0fcc6fed5372f125a470aba2bf7c63a2fe9d27f3ce202680d6bca124ae05c6a548fad1e5845d1a696c53732e916cfdcf7df529ae95197c5dd13650755376c59b3abd40b97da6df627c47ba8cc91d98f66ae8e67900c48fa15586b5dae0a825da4a5d552466245d2c3b46665dca0d989a39c62f2cdafb026637;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h76bdb46f64aa51f7b3064ca0340da928770d8c44487dd8416f2c299d00a7e927ccd190451c5db2d03f4131ac790fc0ce6575de414328eba23ae9d031a94c3aedf0fb6c318a3a03e68fdc77bdf0f692871284106534d5cd475ae3a45db0ffd860d5bd3cec007327c5e7f6673e5e7ae7cbd957c1caed28f6b6d6268590228274fbc1cfc28cfad63385c88be27fc0d70c5b814d0ddb199ea2a95308298dbc4a4d3362fb8af66a9613a0976317a8e58f049fa41e958a85aae0ec086648709fe2bd3c956cb9b93b68b2ac5bad4db0172f3e248a38169ebd8a2f813e1e5600b909efb636869e6e7ae5e8473f142827f214089dbdcccf422609a5ae7e2d29fb4976848864c27ecc04854bd51d33206b1fd647f88214cc384e89d3f41a2bd23a66e68c561a0c08e40abf482999b2c01f7ba88d0304e37e5f8de078c38199801eda13eaaf87770f9dbe905e878257ed29307ca4e2025cf2607ae073791d481bbd1ee7d8d13aaf83b19a1c235d566576ea4acb9e7df1260f78637e86b2f15769b3644bb1d925cbbff31a7a01fa6141e97cb6fb2bcb28e5463b5ad16759b05671f63b5dee0224d6d0004c8ecaa3c090038a9ebca27efdd3d0033032c9ea49318e8b585774273e4c48e19218dffa2d1f0e3273bc5c39d48acb5a79c161ec10a025d86917a6b07fca4db33b06b7de60b291a4200a303eb3b7763ee686d7e6ae045b49c762671f74a0ad66d1e1b9034f656dd3045b1a0175ce025b33e0af529a4ae562744f508713cdc185158c14a1a825e84d574675caddb1ae8ceb6b738db79261e4975df1897e40cb0a3ffba820b81cd0c41fe49537822dcac742e3bbe7037a82f23ba431e8c16c514c00e4ccc84a3439ec9d3f9f37ec45231ebb2b14361d05ae9eb2fd7f1ea31f977c79f9bdebce3646ffb58ca5b4d4d73a6e25d5d89a25f28fcb13498d4fd8c822dbb92818a5d33f651ae2ceaa9992e158529dded837063c130420eaece52d3abc25fc96acf830ff292f5757bbae697afa79659ac6a20733b3ea32a24f313d2f65b506824133d3320842d2e05ca3e1aae834a4fd73a0340ac176d87b95c00297d7fcc3e516641848a356808b86eeee0f89b6e8cf280f5644ef7b5b921d31434b1b01f28cf214b0b85344c739f778a2186dbbf6e9a6086309a82311b0fe7a1079e0d60a806e849108080a26487ae316b8cc206e0fe09016433a7fd470c5d886346e86827db72e9c69b69fc1e587bf67ec7d47520cb791cb50baf4b17f5069aac79dae3aded7ddeb51e567c23099c7a17b6e97169569d797e1242fec51c66d2dd858bc96d00fab69dd4bea24a81308ff7d59c452fbcd282a0940e8b9b5427c71c85cea1adbd48a1fbc6ee833a7ccb7754f34db4b7f9409f99dfb0ca21129615debea75858223481826de1ccf169988e4b6a352c410b5fcda7ae2ffbf7f045ef023a89402d9940332d619793a8665aff7df8ba29198cde4764e24aa4db93fb9f96e86cd47eace4a6f3c7f8d313bb1b5723ea99329269e12dac1b433ac9ee9c05fd96bf5f6fdd9a0a0f8673ab40323e1e4c03d80b35bb567d7403ac05771a4436096da3a89e9dc7d0a997b9162ea0bc076c0301db7fcdcd210c90cdfd0728db4115cd1a84a0ff74c7854868a5d66777bdf100ac8ebb0a032b419aa5f991d5d570b00d51b3935259bd0128a6d6e4b2a83b17c7a951c54b6d342850a1c857e88c5670102c26c06ab28c46ea281e4843925ebdd982c4e04215abc8a2eae530b56eb12f10fdc73ee392fc990263b0ef3a3b5ecba4f26a60764d35685aa9b9265a9fbde8ebc3f7a59f0553d904770da34d3f7a89ff522bee7a8d88b0658eec9bb5c16529d0fad33384760ee5edae8b3aafda3ae097d06694fd18e433ea547811ec4b6591e4abc934a02974a7d657228988712d3c2410d63b1feea33e4ff2d65c8ff1bed87b2f4bb1c219093db8b9d1a2f2ddfc3222aaba2dfe292dc738ac166959ca63a331ab93b9be493f4d706f7623d4ef80eb73e388d13426c3f07adfeb435d4fbf64dc71f0a37e9a694a5243d6bac087d00f361b939454e234007857406d842813bec62713391e1ce91fc2c791f690ec76794808b39fc2c881e7a8feb521ebbdf270250254b2ab90bc2e607886b827546c9e8367f8491efb531103c8c76290c96ee995b6318e7601b3d4cfa3ad7ad3a27336598b616bb127c308a7f48c4c9576ea179f16b33beea224e047bade627a6aeca384f07238706a9c1bfd1ce56f889c4c0eb0c4d35a5903acee9f4c9fcad2697678f2bff73d0230f47a847fbdc09d5eab0c6891949cae35e7e1ae61682657a0eb4db2f47f1769ada56c32e8299bab1041983f8c122137f5066eb0745123b43974e3342d62c97b79ba24271d7c55a36e706cf26dfbe43e32f4a3d29c7ebfce8d118082bbda80a643daca3b57745943aca534a4d9934b6d74bc347161969ce7ad36bca01d15d90e3967a09ee5cc8e2c6803e07775e843d88958f119ee2c3b6c033e4e5fbaebcdd8335d3eab799d8233c7d31ab32bd6eba3061aa25323d9801f977fe1c2221b9a8be6998cba17423e071464657005a2451c293e4a7ecc71b7a383c0617846eb75330a897717581ece1ac5035e42b835dc8f6f7a81fcd919136124058a131689066b12273a26f35a1ba4c2ec897ea8caa8c9d08b6c1c68d1c845d8b1c0dac5d7600efd9b5ae1c31bfc14204b957cffe41abea2bf9fe239dbec4cea02f82068b284cbe2761510690024d64be6e2f20ad6e5a02a8ded665b8af98135892bbde424706b7cf57b780b23aec777593d2c97b619ccf639a5e2a1d4f94c8bf1340c8f7373ae4e5120f10779e507478f212e229becc1620768194ee937ad5af375c2589bb2eee02ce91531d3b867f0b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb9dd3c780ed5b42c0fefb03cb9455c027502ad7dbcf32218577d1cf8ad82d43120aa6461e32758e8aa7a245a2db870a07f0e1308d263b6f2ed447f96851245dd81988dd72f98c9c18abc8e091b75bf3200499fc81e28e962f1b486428d447a830080689bd7186461a512ad0d7fbe176aa7268a26571627cc9c20a25091ffa1e119d539adecb80fdd035ee5dd9a4a0e3e6a21a4bbb9e2186ccc40b75d12b7a04d49dc345eff3ab860587c240aaadd493b0fc9a18caf5d8279f6c5c491406a8ca885620189c64288eb89e7c7a997bc379a2572cd12d029e2f059f9a838cb60913d0d78bc73acb7c9d439bd4ac9cef13306c056c70fa35964fba09a8d0c166dcd0e69a763db5d0b088b403ceee3375d2e069cbfd214f0c4e6f8d4c0ae5326671fba3d9bc042548fb6ece171089675b7d493f2b5a5c886da6161f8ebfe1a6c41850284cb54906c999f13f581911f9a309065097d00b2cac0d376e0c973a58e5b9aa1e2298e55845c0c00a7d9315a4cb5d0562885bfb2496b237abb7f01781e08d7360225c58d992b15a3ca398a9bbe9fe7ac089c4bffe095570bf365523ec99c6b45912093b4a4236859b63368ab5071ebedafce1dcf4d03db09df7aab157bf760067029c197ed537012e7f0d43c896ee2f2da28dee5f26d7876928ef2c06f1a88695e781fd334b12ad7522a298272a104e71defa6f6f40f57921de396453cbf906d132248a9dfaa321033b37240e01bc49601ed39e3c2f84fcc566785dd33cfb422d8d731a727683d87a9bab99e53c866c0f2979ce99c7cc2e85d80d1d15b3b22502802f8d1c0cf5a64b9b2dfcbfc4ade2e1e5afbf98d6e8a4defb6c21eb1e30a5258ba6cc995992e24a30f1d55c6f195da55d662370e3ccff173cb9d27fb27ee6848995d81db82e03c874f66eae791ad841896a572d5892e861ae1fdc742f5cc0dd994e8025cef83d4ed77cc11c7a57cbef91464467145254c614b922e34296a2cde96637c8df81a74208c74fe2e20bb846e8d15f165519586e757c701ed396028d30d7ad3c795b33f69e67d7eba0f9ef5693383754f82f0bf153f1484e9a0fa74de702c9a5c9c9db0038968797bdfbf31fb17e99e9d070c088a1d40f1d6fada154221219ba6ecef6a9c0ee08ae47d2486f102094fc03c38b4d25b43f18cc4769a9da95c8b67fe461f0534d86f212d2087aa4b73efd77f05b0ff3808f93db854e93c2094d26e41b0ff3c98cc1c9dce3da640343773d8a85187744ccd3d648d412baba2ee65d70ac8086a28c687789106c151b5cb24810a39f57ee9981e728f862d36d7c03393199b9417daf520e251ed6ebbbc58bddd1f20e3d9c474f0fbcd16fc74765b2046f6399ae2b21ad6aa255a15a84f07de7385f9e07164ca8268a93a75d54de6b9f8d9c38d7fe47f7e7321698ba30f6fe7fd16d17eb69788086a05494c32712a588fea1252f31abd7a6911d6d5d3f42ae86932b18be062b6db4cea17e1b84960e160faad1c3faede2d2357b3a38cfadb50d58f523d72b1051888c1edbedef38b67e92bbbe4cd480f9ec6384539969ba8049f39844abdda7cc0f1bd9e18a8377815b2dbb4d4df44f04a21db2c898514423260669bc28104224c427c1a2f7e41c7610317f6537c30f839fed14f83663cb4a08bc62a213193331b03dbf60cb40ec97ee89cf897f9213689f6e3220f2a62ccdbf8098637700af17585df87d5df7bb28dd3cb897dad481dcfbbe6f52861793804b2f9ca64cf78c67089e7f67fa78bff0ba4e443bd502efc6ba6de0fd4eca593ddab92e361093b7ee73c1c08e8562d3f39a7e99cca3ab5aa09a1a12d5cb61bb3ad510d6e32de5b15c6388d949617bd2f399a7a4d3e807de074feea4e711c120f37c063327a8adc8f97ff6c552c0aa0608236a98e3fff95541786abb0277933e691ca6e6114bffbdb62dcde7c41330f6c4b6714a9cbca91defbc17a38711a2076c639ae6a06dd01ca8965a380221b86bca82e190d761c9ac46660eb3ca7597e81ed1e7b7d7ed654f852347861c545d69ba839edbfb21fa549d3a6ee61154c49fefd9133fdb2d6894e84aa2bc38c3e448e002424bf471eb89805cf979344b1d293a3aea1e008c7b4c28269889debd3693c8287e43660d66d07f0e094e75718b55b8d2ff892eaee154972311059a798f0bd36607986455ddf6c725f264ca6c01c9e685b761a6c5482568f2ff1ce292ab55b30a8bdff087ad6429d8132bda3a08df48a714e7a9970a55af48117ab1dc76b88b3b400f8ea05f6778d1ad1cf5bf7cce564aee8b51129fe1954d7e872277ea57ea3984b520984be02a6daaa1a1f4f92bdff4532496610e254254188ee2f46330e1bd5e13f5604d3e84b16824bf1496a7dc96ddc6ba47ff31b277ffce5e92e4421dac52043da2194ea63954aa0ce247e93d32e7c11a6bc37557e2600d6299efddf40b99663069f8e55282712347110aec5fa9be4df154f5bdcbb9d0b8a7c8e193dd41fdcbe029973c62be468b617e69decbd4e0bc8f4e0316e8e91f60e7c0242aa9019f689582db5e3cb883a090ed411a6f6f1ce078a23ad326c3c25e7bf48fed55b9e2212dbdf265fc41a20c7e460ddec11a9018e551380a371bc342363ce1031c3b18f5b13d49e0433fec8f221aa5b75b907a95183644fa1f5ca4127752149aee1f40fe51bd5b0eda7b8a4d45500847ce1a756405d49d0fa620a58803865220ef134c88c54816c1a66075845a1eecb46410f1941f6b43c8ac2094919c4ec0ea44344545fa82de6d650d654d75552c477763f0b7eff8bdf4968161d8a318bad1be604543be3f708c40d2fdc4a01f532716cf83da3e13b0414ae6e1594d30fdc56953819ae47fa8bb6f507aa32c72f35e0c8d448a61a7e95597c039a8bce;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6b38b09930cc5b1524030899ebbe6e2938884f2fda017f8d89fd873811013dd48e64f5f0513e09e4319f979c9635bf50b0f8911514ccafb0cf55e97067946edf3d839f5738f89cd04b17d045cb8b720e325e9b24c60ae8a2a776d6753ca33f22a7dcb1c46399a8fbc3b4ca552e5de8a3ffdc2e3b15414ba28eba2548edd6ea8ac1a6a230a0709416e0fe3a66041666d29626809dfbeb6220dc7d5c287503054edd828b62a63573748caeac6dfe882759da1bfca5b36b5623eb713d3f29c518640f2e192539880bf4d851e7761f667a5b46c90ffb81d768308407789264b838c1886cfb4442ca707d9a6be0e19c069f408d2aeffff9885b4a44dd767f373f189f7896d9a9195390f2def50d5c831a2b787f1caa13b3d2e84eec259a0164b4ed59cbf015ef4b2bb069738d94a9a852df1dc23c3b8f79337f654b4746c91e2762b3892c013fbf2a56946ce2979fd73b34909e99050eb8026b3e8ccafb1b4a49a8549ebe5300dcc51d6d7eb74121a4745dc9a6ccb735c231c0dbe8c786d111fd7a6a26bb58ab9cc08c04b71cf5d57237e585fbe3bac2972a9e55a0df6aa2e27238e51a0ae487d87e72ed740c4c73344321f2e283b91a2eba556aa0389c16feea2493bdad5fd01ef1a35464690d2997b4a4fd38ee84d82c889a6d42397775703b3d0a518b59bba0151ad945c5dafe9760aa1bf17d71527f80f0fb24911ed05b9adf1729eb28b2c5553ead676addf885b6a9bf873cdc1e2c36506c04b9b31fe2d06ce02a9e97d04cbd3c028fcbc8339cabaf71f16398a29ebf6b47eb502fdac97af3ed1d95436785c7179981f4cefe1060681d6eb55ac93f37f98f8ef6ec4d9176f79cf610b11683c20b7c3516782df2283bf3b0cacaa4a1f8705b055fe6e601e5c1cd42e99ad85e6064191bdc91fa8302862c746f9be78ec502e39162581c5353a9d5e457f506f8e4b0afeca3a6d405f6f5350d85e415daae30b1f73cb78abe3d27d97dbc4a890de2e74ad70adb8d634c7870c759fb31d1670228fae6844e01a676962efdd851e359463a2ae51d4c13488bdd1915dd290c91d754ef05442c23ff9e040efaa7198a98b169835df842492ec6a492e293ee09345f34024317cfe78d3952703e56eb1e062d42c2292f9f2b20dad7a206e94c9f8a99209aaddb246aef8cf9b28ce8870d2d96e42c43ee094e54e32129d478dcc2e1924b334707453f537a957c4c65821ac9881304f5afc239ae8c32970eeed377dd0ee55cb4de4dfcf6ada60e757d858972e16b5da2f4eff9c3e263d4277d6fe98709649854aa26a8c0c5dda1b82b5172d8b8938f715b158fdcf61607d119e7ef1a0b767892f2d3ebd761dfd62c2fe142d92c169b81851e7399ca1a142bce516b1b9332c3d2c8127b61c94a7b766f6b4bc10637ad8bc0e3af08db4262bf2d438ef682615c2b6f1b4c5234897cad1c7cdd4c8050c5732db97851731e18cf9906ac011e3ff0a3218ea2468b53839d451df76598aea1610e0e8863db16c9f94473a90826c5f5fd0702025f73fa3383a39d9322d6cd50064459579126aed043d3db2708728a577fa5b0887b7730daeeb9be442d9cf46f8e4e7d4c227c0cabe3367f1d4c73d25d4285d2763b3ffa976743dd69fff16498af05fe2f51df885d313386bc5d08003a9da0a6b0f31ab2667f75aa3fe8bd23915157c59bcb2736bca0f6ed6a7a37efb7aac0412c5cef1740acc86d3d5c9920228a0705ac8b5971bce39f9e24b8961a409cb5e0ac3f618bfd6f51d608785b603cbc3cb39465c4acdabf520ee293dc03913b11e96f3b69eac8b9d746671854fe1b65ea2f8fe5ca4ce8057b370d01c6b902dc72305646ff0b9ca199a255191ae79a4df0ecab4d21c19fdaf872eb1f9ebed54baf2906d03dcada95be25f00aa6e9a9ebc4d91b035bf21d6028af2e2df17deeb0e7ae059c2cda335656ce85ad238151159e1a6cac3f3313207cb488ca9612bf6d455cdae004c78abceee0833ac6aa03443c880d4afa25b12e5591274d9a23b94b3af0bf425644ba75f73ca61e37bfe4dda7fce2a14c17b007b71f1135632679541bcb1fdf24d9144f13cd92a877fa516ab9a380604ce43761a5b6d03f1569c83da3d92a1ebe1fe3b61f9936d8e351f94e7fcba0cf28a3b8468c155ef7296bea1062dc45b07af43f3ba28718a1d4503ff304c4c4e7763f77ff9b2e230ec4ee08aa32c72efa81c64448c7b60e4cfa55e01ea452f3ee58010b4cef08ee6a8b860f0374d22930b0ef18db30e522c3dc92e87d2e90e21b503a7d02e7e71e7380fce3c7ce4c4d490639f6611945f4ed3572e6759fef8c259d21fbc7f63781d60dc5c3623de7530e62b7c4325c5f19a1ebc65355ada46a0107580a9ba6d87cb8dd09670a3f469f7902f6834bbbde9a34270d598d7be6bc260c72f65da6ad8dd975d5bad23519f81daa1f463e5a1490369cd694ccc7a834ddd5df6937a5214d8ef577d9f93b93b2a031813de64f1292dc5abe4af4c15cf60dba42d0a7d06f93698bc23fbd4feeda6c73ad4d147e05063d6ac32ac55c0de183081d5af0d803074355d7b3bc3cb37442d6f534ab9b5b84b936468ffaa07d595e599b856c2fac15749f5201bbb42ea21406d7ef4a076e6126cece82d8094242df25bf2b2bb3fe446756ace059e5228b239644054209459b59547fe44bc8ba007a73348eae4fca7e3bca017db795881e3b3c3b06c0e42495916b42c85438370e6ffaea9951ac26e8ff4b98aa6666ad48fe1ad1866ed256f0ed423794003ed67435c290858d90cb99daafc84f815284b0c06fbb9375c6b7c20d308de582d7455ebea1bedde5f9072bdaa868007145379c350156608d8dd9db23c19a26be132a67753742022bce4dea6d2aa563607f158bc54fa6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h9ceadb08be984ab7d58498c3208bb282c61cf990264cccd926f079ce8d2f0b9199232d905848737c4146aae00687e1d4e145da0006fdfb8a2193caadb733244a42e5e38655da79d6e78facd7cc4aca7c0514082e15746ea0b3129b323b60937c270bcb5dc28ce27c61b24ef689c8a350a49759cc8a0f9ed8978df236c5068302e240b87ea64ded0e57be3f4f0af21d84b40ab478e12f78b7610285c2e84a38542ba312b8de26d36c4ba010cdb5cbe787224bd8adc11392f3398853c8f4783f0758bc5519a0c724a1d12141431a85927cc9193128d635d2fb41dfcf8248138b379f3b55b3c23d2fce1a6ab716db7a0926ae0d471c258a489f6f046165250d1523c0aa3a9daafb95d545833790b33bf1ad23561d60b23f79fb35369956c95d7a63748b9637d5b2d3863b04ebd13f24cc6baaf21430e1aeb7f3bcb72804fffd1c1d88bf57a7e1d1b09980be6413d97179f72082ccadfe59519225753ed6f546f2e72b000fd4d2329cb9d93a43f7ea98f90a4c783306e75ee79e47a68994b04f52a2c6339afc62d0ddaf4687638082f24c5620cab20db45628bf758f87111183ce464c13967370ad35d14ddbabcbfaea08e74f274f6c84e40577ae34189c5cfba2dee5b2a93f436057d1e357d2011517bade41aacb654a20d65d53e3f8f18099e32936170489b904b3f753b23b05d51a9323ef87b8ed5ce1000006e8a1646b3fa81d0399102d60d0e09a5d0f2c061d9c07bea430c94a28c022d7be3665e6e38f7e1a1f85922f8f1668408d03b77d0fef6015a6269b19d3363c1866672babc61a210aae958d098db17513bed3e1e118ae907c82c6b985bb61ad4b3120e7b168375b727efeb6bd6b4bff38695a00b02a3d916cb40729c1c007aca68845f51337ce67ffa113676baa13f6b5c17030da502881bbf0d130251ffc55ffe1fc1055cd0f69204e9103bec4206a05e76c43f6aa3a37a96aa074903f620fcf989c3e96d273bb8efebdfcdba097a6fc585d018a03240c7ed83dcd6300c754f7d861a051f59a3624f9ac5df9a3abe36b7de369aa32210d232568a324774e3c5f5afc272f3743ee879b09ee438500af44f06fa592a02211df962748005724cc51bb78ad5198e381914aea908c81de52f7db5b4ee61981fa332c052cded028f5171ae971ae7cb36d447ee16674444095128fbd061998928ddd63140c98946fbce9663eabb3708a9a32ff2c81cb1bb6492f8470340b0903628c1664f36b24e22e4d1b17ee027e0393da9a9a12edfd1ecfa615d2902547dab3c809e8d7f6c72e28f428eb5aee247467d38eb2e26ef24d1150c885f6d59b4bc2374adca65bfbaaa3be3827975b76fc5be92007e51584b9f168f695276ed407e58da916ab1430c23860fd41e88b08ceb480897139486c05531691f9ec2a97fcc771856619e51c0262e1828d5f5790e8f17348a45e9faee8129247fb3dc9da3e282fcebb0e63cc2cbb2a0ca9bf666caaf5d11a8b845529496e626021f1ef6ac1cc51d7923de823fe6813e60e52f90c58b19d29840263fd28342b9918f4449f100e2351389504693fb2f5311a345234c624993ab256e5b57d0cd442aa98f950194959aeb95f66d43093001fc08f8a66cbc6d3db5ec84758f3c2228c9638c8b50f5396073dfa46aaab8a6003a976595a3845dca07690b10bc96a5ab27ac3d2cf37f8631794c5b0123b71e966348910ee3206f3a0e654aff7915b326781cc3aa0996e51c27dba863195c683e1746fd13733204b501709b6a676c5744ad28ffe17fcfe8476d03999e98e53a80be611bd8e7be94c59345082fa3c97546a580bc69ca9e61474d8d6c58ef83a8df62dd276194f2aa0887972eec7c24fdf4a28c05c0990b290cd8cd0796dcb9ac7f684c4ec4812841eea18beed2f9acc366eceb6134f456a7b0740de1de97b6b863143bf9047a2fae4c9b0e939d9b4b29e655cf7d310dcb2ab9f7794dd5ea48156304fd1243e0d20ab9a88d6636ec9c6ecba917d670090ae1d34e1108343c4eb48cd5d5097263290fc6696327548cdc9352995f5661138013a82e2e4744f55d2b35ef93abaa1e6fa20f625b8559f16234867f42c9f1f063925bea2fa10d747daa6cf709eca2ddc05716b1b6f50736f80b1ebf55994f75473841bb0c267f4673ccba0fa1ca60c65543beac51b11a5b064288ebe9b69b46d170309bd1ea8fc0e957b7d8707db0046302cd374aff846924fe29006c68fb3d7dd18d95b5b05063f88294df4402cc115c47b1e7fa4438e8eb491fb7a5e8556c4bf045d0715a2e4e049ee64aa5199e5c706b724c57790d916d7a092e9d9b3ead0ae66302b7d4cfacc0672504e8dddef63b9679412f56a5520cc330b775e3bd699167ba28901eff6dd0cd4e3f977d2481ee4d46d3a9a76e9d048281507753b19ed876ed16ac2987a5fd0a1b5e2a01432f982e699908faafe06f285472b9831c89598faa94c1e431ad189f6239f1ccb40761af2ab8a0a8aa36177ff9b1e1e6b19ac55a191c4ef37107aeecc2c327119d72715c4850ac73edfe604b537afba84d25e24686c31e852ac825a315f8a352000c72a2c83ee0e9443340a22372da3fe50076e0b7533be582a7712ed3b7a8687a9216e4b45f09a24d93f5b6ad6aef4a425ca50e5ba9cda1e2ca0460481239af6073d7fbbad1fcb2506389e38f2743fd6d3248d0c349cc9b33cd963f2bfe21b233e4ae88ba22ffaf545fe33cd94a5ee5c12732f65a7511da28729b312697e7957c080075162ac4ebd457a60a565743e957b57f400184dc926707fbb42a0fe906d1b914a24f625f92d1d13e975d943fb797e05fae6b1d676d860376cebcc74efc67e4f574550028bf079fe240a34ea6bc4294e532cbca6579e3287c6a0d9e3b30d54011aa2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4410e0366846625831769ee74b534fd13b37e00d194f2dc6e5543882625827b99c56d5b5448af7addbe535719d9472adbcddc6b1706e767b4fe8ed3bb475d99ad5e4e074ba4bde31a514f2b3c2b9e302d0ef24016f8e98ea23e844a9ad86a58160447ba2e95804e6a47c8c9ffed59f8aa80fe7fa93d6ae22c4eafbbe5f62592641f804b1593363a61e7319de8291ddc9e9677c3d3064463a54ede518e4d79f595db24b8a0851fc5e8af1cdc89a1956b68b7c6c528326db8475a0e6bfd7e8e420cb8b398c0ec40e4228c7853bd2c3ad8ddd3e407738fc0a04239bbc87ae7edeafd6678d15050c98c9facd4df2ff0d9817cb7e3b82a8b4bd34c9a59103a0d2610626181e84c456c683ea29f6f09912b2480ac971f0651880f549b2b8ccb49fe385fee7175ad1c23d5c6122ef27e2f15269c68bdecbb69c98a8407ab819c7fa38e4c7c036b8ad915a4311006c03e9608e6ad3078aeb2f3c2fa1f225f1cfbb325a75450f8131d2b4091875c2932b437ac291bda6b1776a4ae56d6fc711ca6b37765709f69b8929077b8352141b8a1649414be01071f21abe5b69d9130a212a70b7a774c5f882d7551a21a7722da0591c3633b1c6db0a6100212e1b66b1f2bec52c1bc61f7bf489168d6a6544bf38e1498630e43291249f5feb250fec52c2c6fec7c1a934372403635388b94d9fd78bd27ae8369628c51dbcbac12a0be31f9765ef232849cdd41aa3a55ffc6478e5bff42b5715d911afb7572415179a50969bf72ba16e86dc06cae1c624ab4419528d2e450bd7c21e1cf58bf27d9c639b6881d17af6f633acab765ca802fcec32eabd042c337690f3260227f6ad7f3a743cc85750d6366078ca5f3052a1ccfb711e72828312838e3b6c53f1080d93c50e34e31095965d3f75c970e85119c960778c52cdc82267340f0c34c3575aa4494bc8f3f1ab7cbb8e33dd68e28e4b9cd70a8785c850bf662aeb2a65509715608617c6d617a1fda94dd6d0b41b34ec6c8292a2a7a5d4896da993ac681e8f4bb286416ae22a77e05a5be543304a42b9979e735ecc4267a143c72de5dd7bd5cdc05d54ff68e59b58ed7c6e247cdd46d40b109eb60e4489c26979c8af93b50abb55de8001a536dfabecaacca93ee417c688b474ada8b88b6541ed21c78785753019e444c219cdce5de97c9c021f16b619e4377fb9e9c7203c7a4a6513c9ffca2251e1bbb03e6fe6853d2d67d3e0b701e33df532632d1b42034732898ea0393987efd595319bd1de7c8ff148ed523fc12af52baded0481589364abc39371c4276b4be30c392684f242949d40f6b16a21ca8d5d6b528792d0490d38b0cf9ffa34b9f7414b439d39543524c5dc6a988a5865d79ed3b5d3c58413229fc0a439b04d3fd00d6731def3cb647d6c887ee58114907e8d9cf0209d7661562b9406ef78f070e77a282ad7acca0520c84a9234fa6fbb56c19f2d939070fb11108da16dbf2a32659ba7bd033e41880951e3d5e721c871e5b4cf41dba396fbfe18c9facf64c8ac5e7cedda4eb5bc9ad2e58f8ccc8cafdd99b7e56dd64640b79eb81e5b8a8563fc506c4f7e79ff4884a4ec2b983672cefcde073ef8bfdb8befbd4923295cc1e8fc6b16f1d74d5cdb15da7ac6d45e7c5aa06db67794c4eff3681e89733daa425a5068408879be5d47120e7a44ff2808d15d2f1d5e860defd0fcfa52b7d0ca0f45ec6a290096ec9e5ba718ec7b2184a1c19052ec6c67058a7ae214ddf07b25095048505c336e4ab22002b0559419ae1bc50d35ae711e856564650bd2719c3ccd18bada3dfd80dd951963f3ec09ed0fa0cffc4899ae3b5008a635c6cee145e1d82fd65a9ec5b6aa2c594f58e6970ada13e0c67206c48acf7f8272abbc42132e5985a3f82d491e83abb8da9eb74aec4718e1141c216a58f5d847ef82668852534e4d165c56c947d66fa35bddc872563a19547904b6960ce3ecb8f8fea5bf5768436ebc9496bb18e1461702fa17bd508d74a9b67f801bf9222b822c12174490a84f0b2c25d9f47f0f6e5fee654a0c9d1632b15d6985cc5c57e5b83a79d568395af3edb5696bfdd11609df44e43ca6d72bf0529bad601b6a5752460997088ab39cd9213c107253fab02dac1bbd82fe1492535589ee7b350d8e884c9f912cdfd21f7b994556ade148aa524961c4160b8d8210da0e2646adb5e771e72ec11bf1a963778cc1014ba1333bc871b2b2b7eebde7b54b1258b07971161bd4fb63ac2505db0c07154b8966634a8190e9371b58e88c6d73d1b526eb377acbba8c92437fc3613c1fccb0b6eb8ba8d6230c0ab9e881e6953ca31a307c4a57f351b0e7020a4270a1ea8eeb1b276a784105a21d23698c6a2dfe40a9a6bd328e633bed2d1b31da3d1b5db60d7edaaecd6aaa8f67237c2c5f49b6a173bf36faee3186c9a20132b528ce4be36811d57bda6e1902938aa407fd954688746f6459a99901d0fb728ba080dc54249f08e8eb4ffde19f70de497514db93c776da41b85bbb0181aef698ca21e5a11ff8aeb4f096f4345d887383a6f567a6903526ad128798471133da96de73c023eb055f9a4505c9305211933e62f6581df1e99d1d686ea4d798d497d97a10a254c77204b395df02074ad9815b6979cd242968263fcd229a8bef5019609c5eca99c04ade197a95a7144bf5c6057e28139b2b400fdd476ce24dfd23a1e0e93b70ec67a488fb67bc8331ed8de9b76ebf8a6d7065e88aeef4bfa80de8a505c06d59f36cc8b26535ed3d25d276870a8e23d965b8f6ed23ced586c7ebe784cedb004bfc3c39fe78d969e225f0405f2d4312f49c7d9b7a7d80c924b730d1799ef807e53a29431ac70b493c46598bbdfabeb2463d1e7ec1d53e49d1b00a28ccfc0d7911e6a67dde5084071c8832;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc4dd59d21ba494191ba32594b63194099453613bc4cc525dc909b078ad2f379e96cf4eafd49c0f644ef4f1b4d226ddec5785f4caedb138a2afbfc88899c3b0d6b6d1716256fb367719b7d9deb53f1e42cd9b04c9df5a14d7d52b5268e20e20adc7f5800e37847fb4117b17d2f00928ed0eeefcfea1284cfddeb71ab130d66c6e8ddb3962f442df31757f2020acf3650080fdcaf5b71e31d6927a8cb6603a6114ff71d0a967269e31d8151b22f6b234e5abda55bbd346519556559cad25540b2ed6a25f6b4cd6d65648a606580f586c4c2383e4d55b3f2f8cf4b90f1769e7635297f641d0ce3f7d5f972fb563ec30dbb05020fb7315c891279abedb9e466ebe65332634c3869d88f376b3d6d4a6d9234300e781f64397bf8e6f790660394420a6a44b331d36c355ee09ade9606ad54c25ffbeefca2c20c4793e1433b3532ba252acc6c0e9ae123503114db8fd286225d4719fe5163d963efd25d8909276a29908279bed3a5c6ffa6fd1c4ee6ca95d7a748915dd4e9faf56fa8ecb788d32ddadc9b71bafce0795f0706be722a0ecb84d98ce52880460b091a384df18fefd93c2a6492d99daf8d65b6a38c3689828adc859cbe069375ecfc9bfe26558bc51ef179aa4a3839c681e16cf39aed161d3ae6ae1d671c381d125fb5135229b10734f054969923bae202a7c162cdceef51c206464fbcca8d96dcb215d69607a582d27d6ac93f35e22f3c030cfcaf386de7a967321db7203e0035443ed46476f94c12fb78c64a13d206539cc87d822f2abcccc0ac3fb478702db70a85ef506b69384295c7d158a8476ea51dd6fe2c9c74ac0bb57eac70934e4bc9ae17e954060a3f27ead38476917e636f0e49eb78ca83c9ccc3d46cd32c70f48b82e7218ac8e41c9b26583b6c34074b55cd346b1931f7950acabfd736dae0e530b8c42aa33b180abe6054d1cf723a61046c0405856d091af852ebdf241afb2e30c13df5c320a29852efb95693e4064fae798a0803455ce1005722efdf8d290951fa64624581f75e676b470c28b0d94dcfcd5ded2f5f4afaa5bed0cf934577b801b1fa3e62fd9a752eaf21e71ccdcabd9326d2c2abdfa64db9bdd6323f75c33fba63814cc25d8940db7e356b9e96a16f14719108d7a7e5e1b60686b6aff0c64a62df460833129e929ad468c622b131eda882cdd831ef516efefbb763d3f741856b0be298f73c7d485219cfd15458c4071e7c025a7c155e0efb45af0cac1f689868dfc33be92bc1e76981138524c2961b6e72d3365674735359656d5e6be420a2262b21d1949818030c923692302ac1f8b2d29acc6d922d33135238d0d898ad7f77ca9224594d0e1a23a70672cc721f11774ac0aec4e9ae2b1d414643a9021d973da512608abbd1ccb845bb0c6d03860ea7416da6f80226734a4ca6201f8a18541e929e54c74d8bc4abb61a3f02f7b9ca972beffbefccdabd04cec3f595facfe10084d678247a46e56adadc9c4d8701ea470d6f57898952ee30a9ece6c62e8081dee913c98bca1d9b7a02efc19d9406b1cee174d078291a39b63c839e4af2b28d74f642828f1febe7d16a49a2447da5a980b0f1bff54f34bd0b6d5ed95d7c06515b0039286b5b7e88c22e3635c8a3f9859b46f45576b180d0311b3b4233277a4fa4f0b6a0226fe09c77494539ae8fa2886f6c9e0a5ea1c2ba66d80f8419be244288a98ca6602608570c5eb08e22204a82370ef605fd581ad1cc8669ee1589e21cfbfd93c287ed1e2c5e64ff81e5592adf3e7856c03a0d3aa0e06252f75aa67a48f49c2ce53e7a06cb4f00c3e161c81ba0200ae617c23005e15027f9cca082e800b6c5ceced39b55fc373d05ff157dcf5c448755b2454e8f03f50f6e80a16d6d56f7bed3a2f0524d4a85daad733c1071e3489e4ef74dbd653edc5a2ee4563149d6fc7c07add20cad0fa2509070a84f8e9397eac5272e35c2fc3c98e186dad9f0f83a62383dfbce302c1f6f65cc39b3b5f13fc7d7f9e0382060eb813b0328f10a834fd2730e7185aa125495bc7ebe6993005eabbbe5d2c10ac79f3df6d2459c3fa91a5c2180f3ad0c697eafc0925f2ec14d71dca9a7941ba398a82d64e22c4e93da68ddf0b7ee89d35ee6efeb3de88237cdc5cba1f58abbf2a9df53fa57631708471a3fc7e4448bffbe3d1bea1950a389eb695c3f136b88ff22349fc3d7a715ad61849509c2fb5c7c4ce0620d4af6e15012adf05482e3e249c6455bc358eda8513b1d736292093e181b4dc46e96155c50522577a0467d29885d8dc885cd233e634166ecdb462e3f081300a1e997e8c494be06191f4a5f7acf0ab9b66a49de1709b794885b00438defb2d256dd649aa508522a5fd27bfb3de76fc40a28f9a42b8f98d95a9a32e58e906a739a12754c14e0d58e5834bd5feec0867db3266f770fd034a73929a7c285375e0af2d8a7a15f9b959dfabaf297c5875785e91c4029e5912fb3a615d859f17a9534c94ca4856180271d1ad8717f5db98b1317ddcfb4f7f243a4e5eda5c458dada020a0f4f12ca504ec63a1dc4c1c208aebc00c81480b07d9dab6ae212ac1c8a0a527650d06b882275db8d419a5d57b8c05dfde012d82fb6772bbb1109ad16c82d4f54a1111f2f0409804cf334fbad851a13b60d0af9634126ac02febf82c5baffcdbe34ef3149dc628bae51ba17ebc51868963fb57d3efa04a53a57dab39a3ad9d88958e0a51bd2a881896c8f7f7067d05dd20acef3d738f37f4d4053660150eaf3450b4388beea0eefd94b83516e3eb74080e59fd4204b158eca88903ae7b29deb14735e4a5f5b041ab7b593ed3c72d71dfb8db07e5a87cba3b83891021b72c16b299f4012e570061a555dca697883dd4524eafa4f56f84f1b315faa1196d39cf88941c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h414da9e2d4d4c3ba4e1f8a8bd95534bf25de2ecd7937fd5eb007ec21149cd8b14c0115e2298d451b6c4a13c4a6c83294c272ee3ffa9ded2749fcc7db4cd6cc67c0df2ac74a8fc8db083047679aadcc32d305e45011387da22ae85c9499c07bd23d459d83c2742c190610098db5fed5eb79647a3a95333969b7757a4a4bdeb358b15e506c777a134c8edae635f31e5bace4f64952b78fa6d44006ab3901efa6fb1b30f84be22a28a07591dcf87ed2fc7146ed1a850883e711e7b4a90f258e77183183588b37d9aec86e4a1cb4a24e07118d96a308a5d57b8a3bbd1226d4fae133ca6a81a2b0f2f71182a6e2a67229ad5ca7626144632984c3d0704ce7eed940f6b94642ac8f04c5ec4ff9b842a502a50547bdd9132760a15aa9ef14ad8fdc706849715adcbfea85e41b56f5c97f37d91aaf03d9f168caa53fd7821c30e18634a27170884528557e619c8b606fc36583ee78137017e69a1ea98e12a5f15960e2b4ff337dcc0690e11e7f68357f1e925fb69c2abf6141ea0d63ae00edc8831917ee2073867adc390100f079b6e7c50d5a1aedc13c60fb5d78116778bcb08b7d69db43e30381a81be6d6657c77241f2bbe55038f67ecac448af0a713f17cd72e6e514a08f2fe81a56919f9d4d716979c3f22cbdfa7574281f191bfdc0cfb7ac6ac4c9f16cdcb3e5aa4f6aa3a70e4ec5473e6dc62d5e1962ca188eae49a097410bcebf428abbaf1dc3de20578de4f5e0d8bd55dc3f8b25c6e9f8aa551e706ab0f984f94f7b7c49319c6d6c13462535d66e6016610d9b4f10efab092076706eaec7dd3867c8339e84d86f1375d7e18da6e24f6aad8a334da017509aaecee701000a3715b440e3c0c28171a24f1bdbb8a32c280b9d3a9bc70f63b036ac638ca128ff295763fa66bf0f5a172000480dbcbf9ec1f799661d142d909bc18d537aaa0ecdcac7e8525bf80fefcf93dfbe4e778e13e1579427555dfb437786668df6791977fe3bfa5fbc31f72c515199342fe3a709400bf694f8daf709b2c64e448caed301d8d71f928410f1722054040b3b1b3c54da5c91b109b6f85fb8bf645cea451c4abbac30d25ff296bc65b7be64a1c74d6727cee44b5e9c48758d94c3883a56e88e9e14519172a8e427153ba9632c7e3e9ddbbd0ff85108688616f35e4f7519ac68ce6f57937abfe01e8075529a15b5a970d165e0c9eb8594d437a230319acec0907ac1820ceef590854458ade07b28ef7e80538752af1363403e8ed0307dc86e14d72990745759a0117d5436b91553b7e2e3cab1cd0b141d17122b6e81934f264e16f3fa5163652120aea75a7b63a1f345e038943502c17ecb8012d402f786754c517079cbad1dced74439a7f985306e8fe034e18ab056bb90223898d366cd80bf16b04d82f18c64be56bc2e9d5cdaa7af3475d2a99edf940a45d6e7259ac17ad0b196df4b2e9ae10f43a9fab3ccd750350124021dde1e4baf9270dfd1e601f0b21188fe4bf65c3cb40d9fd8b3f87177b5029864be5e27fb785268ed8fc62a56e354a2465091b6d52141ef9429e4c8a28ff9dbaf9ffb7be1f3a0ac85193970255a97fbfdc5763fb993b4ceced03768347ca26732168767cae9ee031aeebd51ec00d6edae67d1ee7af154808c7fcb676c4169ec6548f57e8ac944206c57ab8a4df8beacdbcdc731dcfe39bd874110b850d5a32a75a9c7ea94bdf1cbac6541fbb9aed17c82b0a4ae9d0bff6e4bf3637dad65bba5da9394cb8613d39e8f129f2a91dacf1de5b715281003dd27c1ef5d588a105ef2638e0a0d01a70dc13a1be1abf0dd928152c23cbab04a66d01ca542602f063087e03437474d37707a41e72a107da384eb0bc7ea60f206ecd67b99321737528e92b1380c7e37f2325aa6768281971db5b5b0c37a5c7572731f266edcbdc0227682e96611a4e134dd78c1f990774ff3ea9fae49e5098a7a4fea07cc6e07fee429c6cff867be87627d8819994e6c517234e3e8c6c40a5b0d50f39342dd58974606654ecf5d3293ea57777f8808332ff3a8ca20d4d131c06a3add5d3005983daf55d04d5a3cd37fcfb4206900256d0247c73edab3bb50b20983b6077867a925caba18e0692ecaebfbe6b748098954604394075143bda0dc112afa10fd2c0ac3d39145f831208d9123f1e6818ddbe192a514f4ed2668c0adcc80dc181bcb5bfab7f3cc920eb8d4ded15ef26dc17a4ca38e0929cfad10415c548664d20c6abb4bdcdf035250ce9853853b2dc7ae7ff2f30f64fa8f0ff00bda08a547ca5af198959d9573c1c4072e928460dd12f0f0ab9339d3008d4377d7f70fcd2ce2406bdbe6844e5c4f423bae0e504188d86d612ed7a776b765e84c5087000b8248612d74b875a1fff2564147de288c49863578f271d8dda73c22cde2ee1f5e8b71eeb6468b92cfcf20351437d0f50f4369d716c2f5783db65edb6280fdaf5390ac8c8222f980b5062a64a66668517a7b602ac4a774d9b8a176b589db9d2e4d09767cee5ef8a104ddefe507029f5f72867d3c02867d9c1e143ab2f1131bc4edbe3dd964f649a88d8c53ff07aca6f9a2a3db65f610245b35c9674cdc4826f12feb6555d66b93b2d5d2fe63a991940156e5d3a3ec6985824a8cacdbdf552bfebb50c4f86e4a25be096bfbe27c77383bef94da36558835ffe5e6ba80fa81510bf8ee3b19e0bfd8a8c76f84d93a929053bdb138b64100eddd723671d07025ac25dbf70cc08f01bd986e69c3bc8891075e0c7a9aaedd6efb11c715aa5401e649615fcb8da0ef14d461a03aedba440f325d68a8e7f70ecfb2bbb7386ecd6553745f1c8834ac948c24b7fa48287d9814970c9aebdcac506ec88be05c67512ee02aec6c45b1835ebff2489098b988eef8633e765f9cf0ebb88e825cd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf0a804ad8e9e0b1db07d82b5d77679f002e71125602ccd92f8b1a779634cf89c6459a5b852dd502a42275384427f4a4bcd62d19244681530986b4ba1100f0d758f2158b2c60a73ce97689229ebd088101c4cb356acec4e440acb2c70b47744db57213e7bc8f11ff8e4581329d540c2c59aeb96cba9a4ef7176d84d4510ac4f4d1ad905ddc8e7d4bc2ca038f019f6b133ab124f542fa9a319d01816f41db8528aa37ad1c897fc471d3c5d4c475c93d4a3f42957191b72a4b85f36817b60b5b4f4e5f8c385eef326512e2cd90d283e998998f72f695307e327505d34df7b44d8ae8a5da83d3839af22d96960c36b0942133ceb10e7d89621d290bf92e2d21156837015f1a04c45472c949a7eb6a7feef16793d215f8e2c29d466e5045664119e69bb44ce396e803f0ec11212e5dcb2259e9502773b1959dc5e60678a0ac0fae9603fa6157666168b357949d00e109e2010981af5fc161a2ef4524d689801cf6259f370c146e85a95f56ae9ae74d4f0809c5bc70532f4331f22d2b47491db1c083a63cf83c754cb9ef5c8462fc5b99d12be09cf5731e5aec698250c7723b37a6140e6edea3dc20a45b321571e0dffb7613b0c128ac4e2e4ee8deeac75dba5755b760c8cc6ddb6428fe33c33af28bd8df41ee65c9653f2be1b432d834888bd062dcad3644e5b4c3f1da0c97bd9c14c888fe5d502761a76faaaa5ea3d8d826e1bf70d7fc4c0325ceeaf9159591e8aff27afa66456469897a70a0db01245a8c9ededf5f1c1b09f7292a31aaac8292ba32b94b7ac3e33d23ee8f142f4baaf994414f9256f6475d809e9f9cca9ad6be3616d2a06c8e4a227b3278fce723d2be19d54cb95f6307464ea92edef58de91a363081fdeb53a7f6a66cfda5e0f6dc21a742eaec6202cf1079d3c9c4e6ae5ef4f9eae6a17a9d4aa1daba4791091e51ddf3ed096180d76d83dbed9b7d28245cb1e1eae3b8a42aa11c382a2604e45fb89e6a910b08647bf4172d1c03847e3035784af04545155d3626c9a8aa4ec594f76dd2345ea9096f349a8270b43d15e3834d4d0350160eca75dce0e03e46018f77c077152563c649fbd7dd40c317cd7a23a839fdd3f3e828d902f14c1aafd54aed12ac060fe0d7589030522f78039dd1fe815e02862de1fb83670e7f4df5ff9620701c24ee3a3420e86c66cd1a0940bd88583b621a48e8a41c54f0e0cdc20e87086f3317c7bca0b1fbd1ab1f69502f965f02fa8960dd9dbd3b7219256f9bd4d2c7a713d431e1b6c8d466114c5d052c60a40ccd4a0409cd2a62f7be1694c879106279f7f00fa465e3045b31ac7ffecbb973bc6d4a2c1562727d80ae2ee6892694a7b084736a1c670f869bffef7bc600b5fb1a74bf5f1727f3147083ee310568784a05df9a34530c189e2cca8f0ccd430520053c6e39aca26bdb2e067b3c9db7f41e72ff8b04b3b84e2a40def97236ed81444e52532ba858ca23d2a5ac7688cfbf4f71873fcdaaee13c59a099a5cc4e95758a10d3405b35e092349834566fcdc3267990089d91c2567aa9c291e1252493003bf026c1a90558a3a3308bf48d8de02ef34aca91c47122b4f0a32c3d1ce3c45a28634230e159a66ea87022b63140102d6a5e6010548c123b76060fb8e9ca1e344c1ae6b533205dc82c79f18d6320b1622f54471f6929954b7a0131f2eb77090de4779a2d9e35cec6317048cec1e369e46fec070a71bdb96b99dd6e45d1dfa0acbbe4c494332c0a2135a6200e2fe184f16a20cfc25b39d1bd650a77b51f475387c39df95db62b67b2007160738f4ea7ccacf74a44edf09c81a0632b7ed74b249dd04e7084eb1b27d07c99bb43cedabebc94521c498515a21107262bd18dd6c7b43f8bf36ea7b443e4ac8bbf8d2f2f35d583a67888e6014fd6a22a7944b1972d8fe9612d98a5747334489ee350b22ef186a774f64708eddb22464f3009eaba850aa0d806efe0a3eb4c86cd543d5ce73f26a8754547e5e1e097654bf09f56630f688d2c9753b5a5c1c8fc266c7880fd54f742c9a18abd045f020e33ada8eb587a8ec7a7888c8e02658fe8f88b3782e46a597b167110f4c4e983ba62a08b2b37935c1434e4510b6f8156318d95c1cc9c5fc69eaddca5530da24577b60f6caf1d9c5901730234577a815e883ceb4611c184939a74e2337c81e42a52b04515cc9562ff25e59ea1c2a15c639b9cb1664b8439ddf20f1467c501952abdfb167b73455099e61b726f50bf9b944a8db29c642be8f00e62cef370ec250e7e97a8c1d1c0b9912b0a4e9a7be54d15aeefaa393859cfc85075d37ced26f7b279969291acf5e37c66e898dd148d59f252a8f0c63af81076b69f45917199a1f0b981dc7d8753fe0c2d436a5cb24203784041c1370bd71081d4516f039c9ed59e1f69bf7c9f2bac6443e3508923067eecb904121c725bb68a6084238661b7c7a4d7f46d8543059971dd0990b33ff52be173e9c727bd22a5c3cb17653b12104145b3763c56ba15f8b42f95b57f8d93409e19fd5af1d6c7fa910752fbe3f946f52ae4df05f5b6a9553dfaca52d82d649886196093a91b60bb4e9697f51448e776d5d35d9ee63e861f25eafdaef938ba3b4d174acbf0102943475b6d42f75f7e932b18f5e6c207fc756cba73c4691e477f369bc6f1169516d7b1677444507387556d6751a4652bed45c8a7d3d34c962fd1e1c712e83b3e3c924d65aea6e78ab2defb8d05c93ef1fbf26ad11f8b3a4242d0cc754765a70b7cfc2f583e2453db45369a20ca5efc603be9b3cece8447772e3b3ef0ccee6320103e23857325bed23bc2bf156a1a5784f11ba36343c158ebc86d8fc92f5c729b55e644cf210b463930f93f7d6b486595b55e4ac1c5b0c64365979efeb832cb3a5ca8859fdbfd5cf021;
        #1
        $finish();
    end
endmodule
