module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [21:0] src23;
    reg [20:0] src24;
    reg [19:0] src25;
    reg [18:0] src26;
    reg [17:0] src27;
    reg [16:0] src28;
    reg [15:0] src29;
    reg [14:0] src30;
    reg [13:0] src31;
    reg [12:0] src32;
    reg [11:0] src33;
    reg [10:0] src34;
    reg [9:0] src35;
    reg [8:0] src36;
    reg [7:0] src37;
    reg [6:0] src38;
    reg [5:0] src39;
    reg [4:0] src40;
    reg [3:0] src41;
    reg [2:0] src42;
    reg [1:0] src43;
    reg [0:0] src44;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [45:0] srcsum;
    wire [45:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3])<<41) + ((src42[0] + src42[1] + src42[2])<<42) + ((src43[0] + src43[1])<<43) + ((src44[0])<<44);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b95a7aa8dcc4faf7df06d94a5195a2fa1eb2a30e78eb059bb67a272feeecd1c513d4f3e8673f02e3559bb7d66f343456a34a3412be6c7b00d8418c0383ec759940c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he03c47f09d0ad9a74b1b8b593e9b41fd53074956b96c986564bfe41c5a8ce5135dbd7e413eafa3dd159eddebfe6fbb65e49f8a9759f0c649b945fec6e1faf1ca0952;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf7a6c9f441ac35574ed1c3f3067de62bb289d12082e56358676e8dde13d3d807adc2bb19a492c5aefe97b6f70e7a95291e895b7e860616adaf5c4dc2ee4a051e7cfa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf21fb892fd014a9cd21934730cf3da2c7b9c006f3e6de550154d21407e5e989ce83f0603488b02abe0d9fae42fde08c88e192638332eb9217b85ded7db2c86e1b575;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h286af3176e1f21b5e0c1bf9ddb4522c600784196e4ab07c38a5eb8cd284a9a82066911312421e248fced777773d4f87d935cdcf81db5ab58eeb62a88425d31062027;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11a6a72812d95894b377a80645ee33cfd77627aa92641088e3b9188f0d67e3f3c32f5fc1d1c509acff0787511ad0426045ee3971f5f4f84ba2bc7c36e17735f309d7b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2456c88a91c14e16ba1f3c382e09ab282d77c424b356a121ef82d0f7e57e38f0b91d7e79fdd9eddd737362cab4721bbd2dccad64927691f9460a2402a5dbb8c98065;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17aca3c8c37508e9c438d6e9578d7ad7a16633a0576a907aeba52f1f5c56d92262436b7075701d60a24c3830bac10dae1985f8690a9d95dbb9ef8b4710746a69704e3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e28ab6dc17fa926b0356a7534ab98a47aa1fdedffd87b3f990700f8e7df1dd104a98a5b938a650ebc3efdf156a8f5444a319c260f4bd09114d91d1524881174d6aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e46d525905503037432b730205b201a5a5b136fd030f78fcd37f523536e9f56de3189084f850368e65bac99f4cdde1de7fb285720906dc470ffcb6aef776404f049f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8cb5d2b07fd90d6f3b65694f9458a9c7796906fecb75cd30383db923b371a1bebdc84e6fb3f537dfac689b08e676de0325f547d9f052ddfc8e085c43db827ca7d247;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19de07ef58f8fac8ec0648866b3d1fd2b6588b87ef170db9d6fdd68258003bbe2860dd3c9ece04f08c4246edbdbc7e5cdadeb5cb6c68367b1ed310f7035eceeeb47d6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef0cd57e06307c24ac082448cda3247bf4918d52a96ad3392b74dc6cf59c9a515a8d08a05a5adc37c334d65dd8a0d3b9f1018f99f494a7b9374dec7fc08a7dae9988;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb63556a414b9ee22c28691f12252f0bd477ef40b9fd89022be821a475f53bdd39f475e73087587141a895809ec0cc52d974c062995f1e163f075f67287f805857231;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f1573cf2b360dc0742d4bf05f017b1a0d3996a143cfb662b57bd7ba1f9003f8177b5bcf454c8c1825ef7c4c72d4585bec11bf9cc394eb0b9eca87b8c7ae09e1f090;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba3f10617993afddc0db67ca64df458c521df8ea29d9c8672a415c533fe004ef8327dc876c3cd7ca08395c2e0012f32c60c34ce8af33144c7029072c700ca94b2028;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1273dd4ec906d985aac1984e3afe88e80fa0f076165323b22941ae3b60284513b44cade4576483ecb8b80f185c206daed11718dd46ac2f8b4825814bead7ad6386f81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd60b46cb3d0ba6507a5083cb277e660be078dd5056a4b3120d5a21a208938141b2568c731753e1234823758a4e93568a29bd7ae3f150e3e42955692afaece86d02c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbcc2e56abcd9a9a7f047b569b53c00cfdaccb866f69102fdc6f4d8a65598184b13a62d403d2d654bd308f84a9eea79f7beef0adcb0ab785e033bd430a47320484fc9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he04fbdd57ee7da7aa02eefc49ff0fe36961bc51fdebe5bdd44e4a68898059dc846573ad11ac43fae10b6a0d2bc2c2ff48e137a1b7dacc1fdaeb67751ccf040f4c850;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a12e30948c133bf75714efb3bfe6ead68030afdb7bccde3b960561ba30dd23dbaec42d291bc2d8d800657c775118532e2f6c2c46785c878a6f1f3cd18ca9481fa0e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h131aa8693ad34657d98332728c52d8460658cd8fd69aacd00fa7e6fbb53775c19823a8fad773f27740d98ce4e5e5461810425109d293d0154095d01e001cf65ad3539;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1884297d38a10ac6b3e97034faea1144d937297ce278ab4c0340c05bc6ae21e658f3e04e4dfaaf634d114380753fbd8ef6c9fa84a3718899f33afa938343cb85bac83;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28dea3f800beb05bb0aecfb0387cbe27f9c9f619c4ae35c4171c946f088f26654718be6dfeef0e78bd9290875f916628b1e1d07e95114077aacd3004d9e6cf1c0594;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8ea041feba57b2e536358212adf1180b5c7f511eac10177fc4cc0b75e1cb9751504e740b1c5640b199d9f86773463ff083f0a3e0dcb5871ab32ad4a18b5359d0c57;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13189cccacc640e006f0ce88199d101dd1a17fe460b258a1f970edea8c777a0c45f9d98828e581c9b437d4ca1e6dfb222b4c91efbae091b4aca869abbaa5747529707;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha9d651af71a0a513e4350bfa4d348cb1fb345cf51c339ec565b0ee83c2ba3d2f6c9bc6355f30ce2ec6b33705a8863d64d38e6dbb5d8b71333d4fe624338a01d1e7fd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d131c02c8996165339a713ac9d8e9d31f0a08124f970d28cab9aa06ee125c7ed001836b6b545c8f689c984c0a0224746ee07357c717a3ea66ee353ea1fc14733aa3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d69aedade388d93f1be7f2b647b0a9dbe08ceb2885e08a1371638ac73630700c7fbdf4301735c32211925a2cd0659f71481122853c079c99a4c425f9a81a16dd5937;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h248a5be67142b0d55d955d654d4835ef6ec48e7eb23e3253ddec97aaff97a3659db60ca70a715ae8beb812e6e1f0756ca913e98d62d2248109e3f3763f605a806ecc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb56febb702aefe647ec91e161e45db43731b897a3f206507be6cf822885438af8c910374f79ac73ae3224db4f4e656e4abaa68ab8a74476bb2c6320d8c722a35c63c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1075e8120cebbede104125d7c8d089b3ef52391a8ca75a1b9fad425baef3d2d4dbc1df46b3beaf88a61bc16302137027537efcba6397cbba48beb7571a3b14a270bf3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f21051a639f49cc4afaad016d79c61f54aeb5c16e5bf0b5f02286b4724ccb6f57217f1cc0f4e0e1930c4ff348c44e11b418f6b333a8c830a50ae933db90464fd54a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97b53826bcf5904132473122a1148b1513a05e2a7c4d28d5549079cb0b2ac7c9c0e72d5d3dba0cf435af3212031138eb623f488d3d16ce9b6f9fd6c19e2e6e7ebd09;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d23e5e063f9b670ef7acd7ec74f8d1372b37213b971a3aeb4fae94893f3de0f53007a77c43cfc2a4920a57948682ea31a6dfd62f574dbe1d052babb624b813dd02d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f4c57e6c92d357e5ad9770ea95864c543699c74f62283f96750ea3051991e6eddc4ba17215c1c15379d6a3f23574c8577aa9591de5a4d87d8147a8585d305fef9b64;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71cdec8ca776f3bbca000575ea90e96ea7bd868e55f1e2cb6b2576c18b0d806a3e6cd991b8be7ab9ce35fef4728cdf97707dee25ad131cfa6d61b0dba0bf52793975;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5327d621cb6c2776826bd5bcc86e8e5afdc9cbc14d6d393b484117a53cbdb92fc75145558702fe62c3c69dfa7dd7030a7ace4c8dd670794e72e40cd67ac5f6211d92;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h130e70ed6e7338cdcab396b3853c27afcb2cf383fc04d21f7f615168943acdfe5664f83485cbaf5c7780955a12eb55537ad1e99da6680fb3730ac7ec20a838235f1de;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1747294102ba1552b5f657099314bcdf176f3e9f64875fa3a5c1038d9c972846bf8638fdc29440f9881f4397589f6db8bb180870b4e2ead82899e1683ea4426167a49;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4d06ade386d6046cf87b5f4f62fb72ddc0ee0011e28084f3c3365a5e2a7878e66d1393b1ee3019b56c58865bc45bb3a16f978fc5fbf19474cf670f5c868c74e18a5a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f5d286b1fa5f9427656d14c410fc27b8bae64dd091f6e16783a729ca2c000fab70e4c69326f5a1eb21f58c8c3f7cac8338c962e75d3b701092c015101882ee21b303;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h596075d22260672eb87f212eeb5995b2bd6bd5b694f5b59f7e5064566caac133b9853e7a25fb9359137fc31f285ebfdfad5afb2460e7bdd1cd64519f889ddd0d8c91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18742d10725800b0ce5ab6e2c563d36f9eeee9cbb8a8004219ecce5988dba4d26b6c115ce59be70fc2dbb203bfae5bf3b3be85956305f4056e26aa47e30031c73ccd0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fe6ff5ae705b465f6d7ce56077efac1f6df0b408b26ab2f4145993d00ac64048e99e2bb02328af6eb65757d17d06576a405acaa56b171a45ce241313e13015fb2504;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea46b813c768d88afebda497f41776b72ac72c135f3fbec9cd562fb7b75cd3d149edb0972d144c95abfe0daf7a8d87e336343fa4daa958a9cd403a2cb6726e510bcb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12816e1328f556da09832e388d186b09216a30ca8fcf448f9834566fcf88f0bc14a0187ff084219ba124a352b8f5af5f88b0c26df7db541247c8dee163afe97ea2cbc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd5a55585d05d76907ebef48ccc01601a5e5e499d01183b61c4a702aa27dc5269e2d54956e9891ad01beb7886725e20a19b0721ee8fe96fd37fd90c56305f1e4c33fd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d40ce19ce7f2613101a97227baa0f01c968f57fd49d218e5c565bee1c2ee8e16c61c49c13fbbfa51626b5d1c5b5223cbe7976c5cca7e4f06c2d3fbe52fc4da8dd14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9159ec4f015aecc920967511d9ec3db59bc19db07af6f3b12f26e0fc5c452135785dd1cc717b9a9da298b6284c7a041b5c9b3830a82537b3f1d200d3e5310644a738;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a29c3528bca9dab485e3f10601807699287f97af5fc75c329c1b019874829a3f6d42c1beeeaf834740bd7d331e49c3cbb71c0473c3448e1cfff9f8d08748e5e79eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfb0b6d13f31e081f9491ce6cd350b3e3f1f347e48291c2b7011c8c317f31d616e1bdb7352f9576ae483d6121af751a3dcdb29a357bb929b9cce12fe3fc6ab6365701;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e1f81e4b87207ff83bdd4f3f7bcc296c4befb84a79b14a8a9372a135dba73b0f16a6c33089398b6e2bf7bff85b1c1d0577759876910b8be7cc3825bbefdb6eade284;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h826533d7b41b6f8a60b35d59df2ca3948402097bd2b2711a09586a19608e61b5922fceaaffaf25a074226571cb55b1127319d45a3ef5d9a2dccbd0677478cf4166d3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11c0cbc288ded93f7401b2b1ba8f0ae17929e13f8b0100e2102d56bcf4cfe35b8202289a3c443b77aef3f4e77c231a5a4ec3679272139cc909c739c2358ad7af3b66d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c457381e64e79172ad1743522e8f42e0416d0756c48ad03bc4d7b20285f39d0938e6e9c24910abeb98baee3ec13f0b4f584d76b8479eec78fea18861df043293ff4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf05e7b0ae99b227555104c9eac2e38dee36bb9e3e9e78f3317c3a18509440d9886520c1987d0a62286cf29d2d1fd7b264ec8b16f2b6fd1ee4252141c74bbb8754012;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d72ffc9714a0fc7ed4d0710d63a6c418882287f731760825943da297d1a532817f28b9e29e2f8253743b34e629f67f4521f692db9d77b6afffebf7fe70c92aefe01;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb632a12ef63eb17f1bad5f12140e8062c35d7ba37827e69826bd48e679dbbef731c945c39b33f2a17e8ea51cc2c1014d51d0ee58678539ee69701752ebbf9ec419e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7dd12f2c9b2513ad3d40e9c5c5f30ecda13173b5068f1de538a371539e663143efd1615acf845369d08ad77d83c7a1720d9287bdc489779e01bf7f658a35aebc9f03;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1db7372be61b6ebb51eabb299247b606a4ea401e13f7ea3770f9d89c36bc30920f046ee8a06819df877b1759d1528893ea464b9334d1d012f0621e9c05305c32d1c7f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86f75ed93c7e6f8675c580d73f427baf5732f23b524cddc21ef7c1fae5adff4d32bac25aa5a8f9dd08cdc7d648e817bf30fc6ed6f460c9ef5a718ddd845b8211031d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9cd9d17da0d2a93aae5726b47eb0f9f8e5e2256f942aabff4bcd4f03f671823a53824372a0df6b18de19479755485ca0290779424e785107389f1e939f85e41a8ec8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2faf6618cee73c22568272f62b28eaabf95993bd5edf3bfede59ff33bb18fbf647edcb0d5644f5c77c676a65068dcd4305776d35ba02e2e7c0d1c3d8fb171502144;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc4a1bdf4c1bac533cdfc3c8dbd55e34a383fc7071bba944a27063b1e606806d22d5f8524237e57f62652297850acc464ac4174356a9d05903401a17657783c15bb41;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d5e6a45b9061abb6b7bf8c105ac01955b3c81741185c01feea5caa60750d8d041e6bbfce7a42d5888210bed70910958030166674d0a7ee4cafabd55829068b1d71a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h160e2e4b154936f8e465f04f67bbfdc75af56b9799e58ef583e3f9618ab4b5d6446823db88da630e7ee5f125d16c7d00b5c9b6b7625971e81cb8936bc1ac9a4edb633;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc440fc70865e286d4db429557e73c484297fe04585b0fcf09c1267aa7c263c42184c51623995e19ed4a5dadb96cf292a6ca83474beffc819131f398b5f63f51a4aa2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc99b7db4778ab11bc1b140cd8c465eaf98e0f741245715819fc3908a4b261c34845a5f4872975dad055d77cc605dbe57a0937cb31280e39cb4d6559311bbd7974fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he8006b9f9e3dea7c20651942f7c9468aa3b0883cd7254c4949c07b2ab4074d8a5e356560052796cb55781b60d93f99d6ac31c1e0202fc230e8329db1066bfa40f17b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h98c03ec6a861425c0b10c2cbc1dc85c405d1dde6008cac3804b2676871078dfa616c9eefbb6961158b8fe4ee96f47e5a3588a539310f6cc6988461df974d6a3bcb3d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15ee2eb0f96a4d32c48cf413a77274ab775d9a98b164a940f94aeef6d29cb496cf7b760842f3624f092b8ff64b6561fc188b1c846687372ca079cae94ddf1007218eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc2e93696c4e650038ec01310584ec303c4578f8f39ee523649f55f7d73fdc84d78b57fce0ae32b39da2df169b579896c20b36af96aec39374f440b3e4a9ae03fbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h102b3771c4bc4b1c015dfe8eb0f7167698a304d61339220ffd6409844a439fa3d05ad3988744406d0340dbf8d0fc26b6ed4bbb45d5be1bec50f2842ec1eca7ab598af;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb0bdd0843a3e10f175d16b2dd2a5729b3f02eff31e5a26d2bfe1246592c35213d6aa6819eff778dd4883acd56786b53987a4b5927ea7d30998353f83f1cbe6cebf41;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14f2d87cef2f6e43d031096041987be385a33d6503611a7a41e7413ff1912b1e5d24225fe06d4da951c05a0aff14745babcef21cf99f1c6c81f58dee7fe8c65b04254;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h745ef1011feabd22e182fbf022146fd598aca2a6d0aeb9549de05269a86564ed9bd251e0d14ae20d18f1710f53067e8ca55df8a63c0343e485a948ebbf41172bd381;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16cfc289f4dd19c9bfe809b533154b660343822bb5691375f0e852dcba0af4e52544b8339d6992ab63ace83e1e5e07d2c847d6c6aa2159054c7aa9ba07011df60b176;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e88c0c3c6e3aa9aa1bfa8493aadf2641d18b4897b8357cc58f142c875a2406606661a03efe717a5cbbf24f03d0cc0380ac0afce6b4851eb3100b294a54816a9da09;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h58a47af1ae6653eff47fc33c71bbbc8d364816f19c830c8a63d0334b05dd639237b0c07f8a53471691e87f1f22a16db05b8604dfd081730a510ebbfecb44647bd53a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h918b4dfe164c3b968b3f8a2b476c8f6fe0e82da10809f4c9b0de120ea5ac550fd0f29eccc9b4cb4e4c0ed6d8d4a793867ffdb44fb79e970ec6109cccd6c11f6195a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19bada5975f3bacbc4d402d0f5d47bd8a2fe5fd7ea0f02ae7b250094aeab0fd1d0d48cd2ab214e8d97f283e9fec42a214670c05cee4d594415561b8a1639e03239505;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hccc5aa5b12d5f6d428fa6e58c863e1ac6be8840686d85f860846f7eab1a988406b83e43910f53093cf71096bb6bc1b504e15f86eda5b276d73048abaf5ed56658f69;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2845cd75950e494c9a3bcdae40e2a4a28ac168249e6e5aa51f05f37259299ed8e08287d58bcc5021b614a2f424902aece9a6b2353abbbfe8d1e419d14f7d54fb492a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h160086ee22e661d97747e22a232d74e50a8a087e85f18374217c462cbc71eb94b1fb544838362d9fb7caf7f4239691536f7a417c920e67a7b0cc316857f6adb234b91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f7b6f89527b915502959aa755ffb2164d144a005f3afbcda2ce4f02a5e4f558bd2677257fcdd3759147df41e111644978a60679a5adb51f53c7e6eeb9d5ec7d0882f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h40d9a7a01fb2c67722e33aa5ae72ba0b76151c2c73559ba281e6e57ef2af82291325dea7b29788fc9e5e1e20faffededb1b5140e03b66672d51e74347a138cbc1db4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf46468ea793c03067dc3ecf1ad0c1dc298e9e567a909e92706df1a5e02640630e5c76e2e67091d6b999d4bf22bd338f5ef5fd4e4364183c50a0e17929f7219674a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103a2f794e16c3a282871b649c134521d4d2f4ee0357ffb880fc5d7094c15f297518a03449aff1bc31ab44628b738f3a81bdd2a6acb196622ed4b1204b74e10a0dfc5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1574a48952aedc2df5e871ecd636a23deb54772a950aaada69cde10621a951abef42f733e2fecd46abc1f01e7b323d0672b62d36004f2e6274a2e02092c26701d53b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c2ddfc6976df6088a9e2b52d9d31c04a3e10378e5e6fa96fd2dc0479648d11d3f973109f3a7d8580b3c3e08816a90fbd1c388e5d60a008d9f66dfb010ef7d3d5fa0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3264fdcb75f2a82ed00a6649232062a7f139ff9c3d1989dfe2ad6a78647544144f6141d30ec51f69ab43fca9a5a4ded2113bd0ac0044f6129ff3750573a1133f97b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6aac1b7d6d2ae67f9360aab91dd96f82d36ad0e858ce442ef79b25a1ce630a76867280515c6fdb3ee3719af47f29398b026d168f90ede246268e777b1fca66b4eb28;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h768fd8505f42aa5c74d563fc7535461f115b000442b0a7002eee0dc7e18dee795fb8fc030c884e68c8496ee67907e02315bfbc3e71310fa8e97ede5cebb337d09f8c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf0e57c784b4b34a92ff73ecf1ae0ca5b20e2c88341c028b442dd4f1442ec01d2788d74b4367fa42432b270ed3b0b94017323a8234704b0179a599d9a9b2ada0826ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11efcb0900c2c67b5a1ccbfac91ce3fd27bcfe15fe9c5dab6f3a01240c6ae040a7a45235660e7d1317b2ad4c5187cb73a1b68d261d11be7e7b4b4bfebf044b2689ff1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf613b918376e080466bbe10d698cb7df4e872ec2a3ae3be4d10c810238dfee8d2552552b8b886fba39d47baff9d943f93e66109e033f009f4265785cb2e163f74504;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7db4406527ebaab05ee87adf3706da572d2200c340d285d9146d65d0e8fcba1c41cad10ec203480f30ddf3fabd171d8192141fc96a2117d204186dff004ae72fba9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ed1b51886a3063ebcc47473b73c34c42768dcc4c49a96569afb73667d185ba4f14fc6af02112b11e103c70635a6875c3529db95591b89495dcd07dbcaebf2fcb9ec5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h85939d55f1892f61d897f8c2a517094a17a975555bdab9cdf5423a20fe19b32819e01d4271767ffc8c04488cea11f131be3dea4ec45c0f012d90613f5c9105a31e5f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97dc1e2ef47ce458bc0abc8ddbf963868aa164a5c78062820037551191a5c0dfd905ed0390ab8973ede67c84459ada40fa2de6c6682fb75173ff3784745cf28b6fb8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c68bc59234730d2945ec0a0d465b9cf1dc4d24578a9fb60232ee9d72b316bee5311ec4942cf252b590db24fae1d7f5c6bb1b9c1fcf392d5518785a32f1b98d52b39;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2f10a92d6e7ce01aa47094e0e465e1be7ec6305f60100d7bbcd5770fc6e5de53b631559f41af27dfc3074a615ff390b97587dcbfb878c2f2933dcb31a0bee4159b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a14873ab5b19f682d5a1329622eacccb33d192dc11f791dd4372d74d8a5b671d5c2d755ec8722846cdb2ba0df93dc2b2859f2c486053ff75472637eaa345c6be466;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15fe27e9f7f59c09093dce4c76317cafaf4b7b7cd63aec98b4c6e297bc9e74023da60eac33de68ee3626af47b1ccf029298108c704b1c57f500e1c127d312a4f4463f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha98cc91be44737a342fd9d4d15c40d572c37c5c22d2ff0a5ffc0d6ec7568be11149cda4bdebaaccead1c1fa48ccb593631a365dd86482324716e0fb2dfd2cfe40eb4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h216d616c05da34ff1c128d4b049794515637869154fbe7598ec0b42c638b1a0c100100dac0c00466cd6cd52cecef833ee4437b158dc80ccf7be969f4a67981820e78;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198751a12cb6f717421e3e0106f1827fe2f3f8e20822cd9d22ddbd29d4ec53a7880b0b9e6194d30f442ce6f99cd2ddc72af4792347bac0a85b8d38d0266ca5560c08f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11dcdba82be8630f2de2355f950cb5f4cb75d85132b3bdc9b3d997c9f7f9a3cb4050a7745de0d74afc3a356c6bc0c8e56097cd2fe5b39e53d0db3b5dcc7f36baf6d9f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105ca9c0d80f93a7d0376768753fc5537ecd73e45a8612afb4ec9866829e47e1fbc9cfae247c67086f4f36356ecb4ee18ab3cfffb36a8ca87e203667aa17df211f4f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h552f2917ad0c55e649296a949022396bdf63f5e0972f81eb22f011e4842cec55c69caf090995ccd34f0af8c6bd3e7ae9be9a889e4af085c69413ab20b3ca7829cf4b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c6faf09d05cc8c60b6fdeebeb99fcc4a8e3704b09dd2ed09de30c1a72fec697e61b0d3c49754cfd59367050a3f97a91aef12523ad3ad31559ce3b0d33b5d667e455c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3e098d63e75302ff2fe149d99b4f1efaf5b5cec8ce9cb80ab598a023559bf6dc27c3b0cb887a1fd1df80738b114a7fc6c963ec38daa338faeb7c63afc42234c9b9c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h176ab18ef693621af9a6b39395fd93a992a1a74b9e99b245612055304fc9669e6ddce5923f3a583b515894296cea5b5582e067b8f877cf32d0651f77583fc9536fe96;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1308ddd344d3f8ec3a7aca5a9f50c8812f43fca11bf38d82ca2bcae19399f45f8fe4fe0f64f6d257f127c397553e5563bbf3e1080305ee54ed83bacb58b229a899fd2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1caba3acf8c98fe30978c7b615f7f88e9254a27cc591763a55172226fe721b197eed36ecb8980d44be5d6e0a77aaa0505a210940bcb4f3299a9e560fdd6260b5f3f89;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7df658a6447a5a8cf62a07f760a8721110d18e9717350c103aeb4cbad188266c161624facf0cde5461ac354ee370c03c065caa6251aa07a8e02addfbd099fba08c36;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hadf154182df26d1242670fe89ca93a45d4b08fc47f6783e7a2c90d70d698db15c7c539c1ae6e8755939f4908a89428f1736ffd10709e0e1c43313659a5185a560c75;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1388f675c9afd6eadb8eb66a69c2e3d53cc4fef9fd336073b769b3610d81699b9a57725039a3f011931c0dae0a4b9bdf98f72fbbf95769614bdc7d8a7e555f2a49342;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ead8bc9ce423687451597047f826c15ba7ef62ffca6cf0ba3ff9828402f7642de81e97552af1b0d4d369932a53833649502660c5a59ee1179c878b147bedad6af28;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h116081d2a97926c4fa063c4bf038ab554f95bcbe862ef04c8d9acf7808f78534ebdec45fd00d123392d0195384c100f1340d5c99fc2f0fda76ca363b26871dfab211;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7af1bae28c134fdb16d5f159b4173740fa48398c0bcfb86eeac566a999499cf0bf798cd15bff4b394150596cb5ec49442af868c839182058e6c7f5bb4f4ebc88adbd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18505e4ac37fd20e2d3b5c5af8aaf13c04626d82f99b9b5db471ece876f722c6c757edbb868db50857e892e1df2322313f0ea1c8a12d30c883c6457e6301c775a90b5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eaf513ac4ff82246c4d537fba66689d928fc0ace6068fb8d668c37aa5c39264a8bee090de30f2a37df5cb5ddf7755f9132eb22983259d5f8790ff760acd9d53ce665;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ca3180967ffec3f3e6efdc59959e5497af9b4aeb1bc446ca2ac8492bf813965b18b0d63bcbc1532ae4680b7f42052a9164f4a4e207913adddb21e94f54943298b863;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c5b49a51e2e149aa818e7ab9d1c1d4db333ad9f22a48fd764c763458fd2132a19a31cf68acd6782edd702b1d3cb5402dd68b29188a4804f5b1c23fb961edb945007;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86945f9018dd26db095148f63bace4db0b4bf063888517d025494c4e405071dc4c663be664acd924f62f0b69b4b0dfa9583f88e66f445f4e490c72389029a9fc5d9c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f466091e7b2b7ca325280518c392678a201c820f381cacc07ab5916ebe4339183ac244dfc636e87b95003947ea05a6354b37a8976e60880469c33b03fc21696997ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h899484125e86fcd6fcdc59a8cb82df64588af980a06b4b968f6426510b0f9ea1d1e4961cccef8a57b3348a4afa8d5c921bef058bc4e38ba72f8bf5bc7c553bf683f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121967a662fee1aca4fdc52c579e23fce18dc82c4af711e0d01dd8c0a7355e33db01bb29e7a6b9e3d717f39a934e9304356a1acc845006aa9b8623810f874ec90dde0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h125b5a264588d4c39af9a5def744d79ce9c9ff694403ccb5a6bb3a83c665df79d4bbe68f61af628255dff7251e9e023a1a7fbb325822e4c971665be861cd53099100b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae62272cea8085b5a052e9a6653c33e7832a0dea69d8ddb888101fd5e6b3c0e88eafcab2e32e09da4aa8e2f254b746208534ae10b44fb00bdac61671d4da3ab332a6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f63e37b8045983ce6026a38c869c90baf3ae62be96a2dab9491dbe5e1b77ea0855443be3657552b662c9dbbe6453cc1102d5f3eef8284494a6cdd14ff7ed35f642b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a5612d2ff77d1acc598be943b30aeeb9e95d8bfbbc1f1c477c81ce0c1361ed8c3d40f5dafe60710e6da0b58457babb31a08474e6a387aa9272cac82b96866dcc29a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haae25ef7074c35b902757f7ec67fdbf535afb96588d771d379406770c573d98a68f078a442ed10ef0d32b12ceec0e1dd3b20bbef68bdeaddc15f900f614605d2a318;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h181a550198592140697a697c90e664797b654adfbdcb5ed8ec1cf684f51fc5642d42956ca36cbcea5127beab81b838bd42406602f08d20ff9b89225d3b2f4980749aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h174ca089affedd1b96eee7ec595ddcef1801d1d85dff46aeb7a3717f34ab4e9e2dce1fa0526d18f0fd51ee330db93d9f0a6d48985bdb4d2e6c981c60d46947df489fa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34ff90318075af4560f2ac32991c38522786eca508e41515fabc563a9e373c520ae8c389ffc08454173b9778fff2601a5b716dbd4f641a95b3775ffe69595f5ad3fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e9de412d739fe7dd6eac97b7da8292e26c2261ee3f90538a2ed7a0b4ed870f703e5adbc4ed19b82e50308a6c7af6b1f2367694c959dfe0194370af1888cbb908d1a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h132fe0ef8cb056e31c942b9961189b4aa95337e2d998f3f6ca54ac91a60d71e0b1da4be254fb3ff70d23feb8e4394c72eb02d774713a74c4a89a301902eac3e45d379;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0221fa26cd960ab8f2bcb5a8ac53860b1319270ee895a932271cc01af059cc4760cbcd2b59dbaab5ecdb8d03f739a05619fdea5e00314a274a38fe78c0e4503aec8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcee3eb3a03e7f131c5c1142e92102d5b5b282a75a2e030a81cea3015d299cb76b8c74bf9016cc5fdd7742cd02344bb59b1f7d3d15dfa8a1819e04c44f490baf1263c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17b52c38886c0e17e1d176dc3aab76e9dc04a2519598b32a984a6c56f39a75ad2d91569745c55545fa2ef82886d5a1f31bb3a2582928c4e2b4ef5b10f510580477d1c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1003877a4e81802015291a7707acdffef9105c0e6a0c402a8d7f0e2c860d135dc18d8ecf9f9c38205100c0214e1d56863763664aa0b6893d09aac1db1fbdd1f464daf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he837c0cbc62f89789689d1fa38df80b2c2a64a3f9a339f643e6a1fc46a0ddca26a90b174c0168e2e4e9f0e449f8cd7d4a86f7d9e962475492192cbda5f172082d1d8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe951f20674fee7733eb17e187aac1ebb8d7cf480f64ec407cd50e70ecbc29f59fed832b5477f27a9135ce2927ee10ca0de1d745d90d7b8231136cf56ae44e6848ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h85448f26f56403ab7a9962e74772f58adadffbca291efc6e92d2544ba7c3f11c30fb3e54b7426c35c6d2df50791b89bb7c7a886e3877d01ffa811fdb70c08280e495;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6158bf59816cd07368c4b674bfacb81e972ab8c2cd721734c756f425dc62b5ea6dd3edc041cd776e05702b2051ab44999a718cd624eed9a12be527fb8b0587dc2e1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h140e65749ea4038c22add57ecd8f677b0b7d7a3fde8e068b9e6d591a12743dbda6399c759e32272f8ab8c3f5472ca73a47dbd317a5d7c42b0fb61d39b3203c38ca488;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17e1f393857122fb2946fb737d1b881e3cc53986e0fe0b11ae8a4b686a3b1f515637ecf00a58e890cb6b48bb2adaf9cfbbd34b3a685d265beaa8133d65487b2a362ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17e8218e90b03dab4ec505768094ae66f1bc340a762a658b68262936201620ec0a78ae6070ea0e8f9cd2aad551c727b47aa729229862e1500c146903aa6e7099113d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha09cfdd87b1a36a58414884f406ad6347f52c132b23deaff86f26e514466c45c900f70c551880124f139fa02ce8fff95d3b4ab1857e2f0810f3ade56acc8bb068445;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1013508364aa440b3606ddc415d9007b8be9883b93266ee7a61a65606fcedda88a5984f8848b6fc0ee309d3eea20b37e6a734ac3c40347f491fc1f0e7f577c27f6c21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1668699277950807e805e6ca2f406e0b44f93fdb39e109f627510b7c3b9af24406670f4b16976d427f1c5028be9ee7455e02a4a838624f8fcf729e60acf336ea04591;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6cfdc13e3830ef12a4647178a9ad010cb32f0e806b79beb6ea13a9c798ff2748a64c97ffe6916ad7a82958ac5c46e3c5170097f8d6706641db9b958ef7b076375b17;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h887099d51d304b7f9932c969174e11cd05d5f377ad7d07c072952852c7c26311e7b50354ba244935cd05c4a20d5bd4ba15e5a8855d57791a94b1c605f52b5f8792fb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12d9c8a1a7d3b758daed8b5445f0350800052f2ac1f0851823868d7287978e743f07eb14a40185e547ccaeb1c120946e16885ec563341b87576be905519deefee52f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1afdf4a88a16aa730126fd3663878d5dee36306b5f29f7b2f3fe4a685adee03f20cadd3a24e07263cd7273b5d095bb69d7ae09144d271d8c0fbe56dbb2dbaac4ab854;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1210ced5934352f0dcee5ea2919db9f3271fdcffd1acb2fcdbbc4791e1de1bd8722dc5d9fb8df169c2155d018ced46a600ffc909c8092be1e1c24157af31cc9d09e34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h540de0d94f7014bd652c94db84fb755606e517a28962082e8dcb38dcc36b168eb23c66ce4282703da0abf4c5ff8f35d2caf721889761302e2355995bdc34b6b26b9e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18fb294af92ee9969915d0d77cfff52f6f3515e78996c82efa3f53ab9145f3be94e9a70e4ca05fab6267bfbaa0ce589c58a2dc98d264665328f7b019516769b8fa032;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a058aa9205197b352dc2448716de5a483efed38ffdb5932e3ba7b55bc1a1f18995be8a3079683ad406f2ef7f9adbb5120aa5065b197270e1ac6452ac441464c2386;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b085aa95052a4b65a7fe46f90a548ddf20a5992188e473ec453d40c0fa7163e81bd4b34f5ab039b6f900506a7233c8a73e8a8b0c5c744a2a9c93f25eed472b6dc99;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he03cd59cd5b858783e7f91049e4a2a645c36bf0d28e4b7907f7514feff387511b43204536a14b1c9d393fb18d6640eadab5835174e589e0fceb2dfbaf6c19a05d3b0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7ac9bdb397185b4fa6f526c45bb566ee1594011334343fadeadb0437dde1281d65671b1950e9d309de07f95604d024b940a058538cc44bf8079223c55411ebc98ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1245562c87448755bcbfe567492e23606f3b51513d5feb727e8d16a42f3c26ad226f92a6a2c54793fcd1e23d419c14b0a6aadcad6a265d76a2603379847cc319fe94e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1845dc25ce9468ee1f97b74febac1f96af7b4a338f317da3c8d8427dcd83ac7264465dac4fe130166a6dd24c16ddc67df175a22eb834f474c04465a295bba3745e999;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h33c6853ba0d0a5dde583b491428a7b3651f48c926eb063b81231c584d7c0e4a291e71d9fc57ec88940fed7d3fd45575b63b510b340fa8eb9ba5928aeaaef52a20cae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180085359dc29874cd5347e8181267dc92f7659647ce7c12cb25f96ade208773449a302b8369a883c7c5f5f2bdb5b3a9cf6f159879a4a04a2ddb218a0a54423533562;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d7d1862dc3dc3a5107f8c3c42eb973487802d18622fc2b167065070e5d2f236843c091d1929af730926d5b3b17647f051798ee3394c71f85e4736fdbe900018185d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h153176ee4c19844c84f0cc73e2b65db7bf1b88f196ec749bd6a3b81057233a57d20c3567cf0fa81458a78c44a6043d998bec95c5093e6ee05157b1fa8f079704bd2c2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27f46be95cf979b16771bf991fe54eabb82a3ce37cfbe36e43d302c5a15a21fd6ee1496721cbc51088ada6b79a76b0c26c85070d69e4fd4a050414097874e6c15c8f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6eed8e69141845348066fec2a18ee2fcf7e7030d839b8da1a65ca70ef83777ad54a191e8b441c5d1ff0bd5f6e3127fff8c40a233b2402941364076194a2ee037dbc2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f20536e3fb086bdc2b7b40dff82d227cfc10c10b621bc68cf65e529d40e8001f2b464327db3770ac256682c157b2988c24c7f205f778b9749d9d7ac5845df0e124;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h158d05f5d14636600a4e6bd83b8141dd149046ddfb0c22fb90ba017a43af701540231103fc33aa4eaf7cc4a15bb25472c298a2063f9b382a0d9e66ad1131a2c70e1cf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b0c938b05cfbc662de3f8ba14a7f5e98a2130d65d4055f3db54f0fea1f9254b4629dfc7b0b09ef8d16667d0fc2049b11fceea95e44109a929316657a421748e427e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15bb4767e53cca9bf2eeae9ab04843e1d9fe85f8d4c8dfba0d12476b4056317eaabff22f433e0f5e8fbb4ce671cf4d05899251b98c728590b83618d7806baa2e0d67;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc1d749a00bcf84eacade2b7c2189f3d086e3bc41253be20751c57a5e3df57a413e87d624a3819acbeb8cbb171611481b8788069e3eb75a17683739907fd1e272829b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a1d6ca54a5629dacaa1940cf2d22a7f63a07fd83df60364c03ac27c79743e2adf06f252cde4ebaeb371784a44c23942d86e1c3bb0f45b90fcae53ca7fd5e00774c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h137099096c085d498a6f2da030f9b418b481f1445f8360742b802c41750fac6837f2069370992e249dde68985aba72fbffe8f7256a80a082a0b6dfd3dbea09f7e353c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27558953d07015ca721df5c1944c17f0771ee4e42e978ed36c3507c50a19192b4ac1628a3e2e7338dec912742d6384a10f94da03026cdcf3fc3af26a876a82212c8d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f2af02d68701d81dde80ca9f47a3a5f7a27961608eed190938179bf48704fa772f32c6e389c50d1793912f46b3a6a34cefae1aa0eaa363b64abf7b5c120dbee95f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186a239261965cd005fcbf55ad8facb0d15a8b0fbb249edbcc6cf2fd8893d86bf9485dc0d4473fd787db9d87346ead41dd8b6b88cbf97719a4bad281068c2be3a59ba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc7db77676cec715b71e0fc2e707edee4b56ba4e9a6b80123a6ec571393a8558652292cb70acedbf20de84b76e2eed83b2c06917355b5be4cf86d8b9615d932da3a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f053b95b81360ea27ccf88e3dac07a90388511759249d7f5b07e463009ca8a583ff67bd5b129d3b046fc67e08b5b97b66af773580d76b3ce8604cf1b04edb8c61940;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h141db9d21cd80eaad52aa0400feb064883832f8bac72a9f110e34d254d05b2bbdea9389cbb7c18c11fa98c07921ff3319c3a33b6ddc57b9758284c44b394e4cb61146;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14986a432b9de3797c337050e9bedabe3bbb2d3b2105cd147015cf54ff2fe2086363bdbeccf94de61083136ddc4841adeabc39758f6865b8d686299c9404716b4e02a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d413124e5597368c880e28e8ccd438957d159ed6d8e443958ba7c92c803ecbb76ab90929200b5d17385bfa06092e5ae2329af262d1d29290b8deb16f3ce3d0768994;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd0730a11437dc36720966857561919f3220bae4b99381089618d907413e5377e76cfbe6e5d0ae1453fd1bc6c0ff282c90625a68fc18d38cf38eeddb4c5e826cb302;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdbc10160ddac3cd3e6e45fa09f94a2dfb99be6b587f726fe64e60d451b778e9e627d481f8d1cf891cb8352b6fc0e3e7160d5377524246b161f5052928c97687515f0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16496f73ffb8afab6be74024bf02ba6eb7f7f9c2fa5f74b60794875097abdcac80781d63ccda55d8d357a6223a0c097fff64631bc1ad7c9923535b482779b86079def;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h917e3ea63916f35c1f8068892234aa88aaaac41b96015a2fbb36a0d183c45d7301da3c344fa3f25d2712c5ee3a9eea6b336f11103756618de3adcf45b11693ab025b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a7c2b15f5d5a7813c1b18e013b563af3b57fcb658dd84b1f00f39af541ec5a9ab6b91bc4300e2304aa92ec4608bde0f4377d0de192cb9978e58f6fb6f286067323de;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b64d90bc6c5cb2442242980480e4659e3da94c95947bea565a85e8b1fe83cbbb86b68e0edc9be0e99f3c7e9969b2d416abfc0fc29ea4f9560c011a73c5db14c781d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105bcb097bf58a1a1615722bc8883e947ee5f2b4978484003dc05efef71b1d2a1bf511e3a58c66998c652caf83da69b998fcb981133e6a9f5d80586552caac502d9b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h49d254c2c1194b9655e295196d802734a2cede8b188872ac9cc038081ed732b6f6cce4a8a308425d13a05cbe9c52fb92a372abb70dbb147e61e235a3297177b63313;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h145dd3edc12cc634c181ac88f73cc7cd88a7ec66f68376cdbb10ca2216ecc1b064a558f7318bd2a0490ff465e5011d74a5e6f62f2e4506248742403e1a7cc9c2685b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f66dd6aba5f43f98e2f6ddf8c6151a156454f23ed49fa3556f6ac4c97184f4301bd8e92592eefe98c352cb6fc4ce7efc4b31d7cb0c38b06dc1ed5b029b922c711d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1616ee34bdc8f2cd61f318780a43b039543004487d8896c585deee7cd0defe705f44e0202125d1a9cb130e85ccd99f12a6ec01e818730187ba5087a70b949a6981feb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd744f0a3db2d8026f5e51c09595c401347bfab5d9a78fb94423c5dfb9e9c943300d96ff6ac30fd7cc6fb419c240f77c1796ef05d7eb9ef86873543585a4683ae2549;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he83ff528f55ae0c1695aa5fe2202008a50f75e73761b2c9e8d5d82b0884a66e43b3759cb275ebe79ef797a254a59f848ce57328363d6ca2c283a15f09fae5622bc23;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h104ceeb6ada705a752e86742f844fac5af4dee9783e6b9779b3c266dd3afb09e958d9cffbfbbad19328301bff2f9f976049ea26ed7dda2833bd659e963e8ea41065d6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a520229cc4400455ef05c576cc9265821173c42c732fb8146335e0e492baffc930cbbcc16e88a8145479637609e12a8226357896d54b75c71ef35328b906f5f58ad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h123ad12e6bac4a22a4744b8153269008337eb71ac9212d9988c4e0f2fa04ad97a4f6a67838ad612574b93155d44049a0e00d501bb026e39eece10633b8518beb0357b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f5e0d31f81eae56be9f1a329310aaf3293e99b3098164c7a5172c3739bf9747a00bc42baa8995c2e02008d2d32a686aea24f99efc22e8e137c8d301fc5790700674;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c5d9d0fa3a5e61645861733febeb0dd2cda66eea3aea5411bbe939fb9f8fe260f18d6c599b02c6d1c32cc55ce14e8f0cac5a122a7c8c96488c0c41f08bbbd812430;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96efdff54a027939b192cc1d8e4e40518ee50529dceb4854ac54e4c1a54e02acfa8a280611fc9999c58a103029ba8131be657ec158e011859cfd3ddb8a4f3a4ce525;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h166c5686e427d3936b8381ae29d9c66e3e8dc401f15fdc1dc728692f5d155c1294df6389827f219c9d5c9b77502f082a4c48464a8489b21a69c63af064ba6006e1837;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9892285488d6662f46289802bef44296c2783d31f07d93ffbf45c396089514a1b524b1c8e101c576649505cf11e1747b59064a8695bbd174425c3e7e3ed022a03e44;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf7c1b37912ffa29c71da68045f9c9233f473b2aed1de28c8d9894941eed8aadbcc92c520aeebbf767c37c623ca13a34451ee9e0ffde897dc756e499b8f40aec0139a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1849e202911f3e1517ba5e23659793e10a9d126f6f25c3c11c97ac79541661653beaabe8ee1745f123e56d645173b3387ad6a05e34673c88f866d0d5c1db48f497bad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e09705da32cd9a8528fe6c0e08e4e50de0095f73cbe5f400ad3d398526d5887d5deb8ca9e3a1c45af5abbbf00c5907e28b2aeb321282f9e2b40db543a320d16c83b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15676ffa5b9b338ed16595f6810b382135679a4b7733fb33982ec365158560f63188173dbd957c11fc5ccd888d318ae030d7d0ae96b3db8bf2fd9efb45bbf881757dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1be166bb5fa84a07c7f26238142e2959dc3489835f663ac1cd575a46ce6883ac0b795011d9e0afcdd6b70b98cbdfa640d7f7b572183372a646f3b3be133221e4fb329;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h950a229c57d906d943c40cc6d71e864cb7a738230054a737309a327df11226906889cd579df6387f458dd42fe1a3fa832edbc606ea21f14da7a1aaf38ebf4736959e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118377e216d89b052752c125c1e19dc16daa1af3455f5bd8ed278e060a5f885d9b750a35fda17ed35e47a6992e71ee8b3db1eee250cbd776e7932f55093abcc30fa3d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1236d46101ea8ad569eb334d93310288f9c3d44a923bdd38542ccdecac01aca5eaa07a0dd452468cbe1365f669fcd309348fc236290f1a95594915d0aee008947b1b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5911935ba6ccb42fc455ec6c90da71f729f8bc2c22b1d63777b35a34054539978a55d5f1fba05e3b1182cd1ea10ef40b85951950c7c7d81ba292cb39798768383dfc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17fe645843188b6492bc45c3a4c4cd5e3f381f3308bd45ca6fe98a913736425f3d76c928a0bae30ec8b3b51524c63e9f8e888de62c5ef34e30bbe51d9dadb4f128e28;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h178763de0d54d1f87d0906b78cd7dac617b58d58e58e3b0aed597a76a57d0d98cd13831f76e4a899343f4dbf0b723e7466c5c846d94aab9376a6ff1b2031f46f9c75f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1933fad3507734559c94df1a9d3cf936489c8ff865548ed1c60da120115fe62b60755534dc679454a62b8bda36d5b7dbf9af5f42f43e715320d7cb3c18f1125c8e9e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3611eab53b615de6bcb469474d81cddbd6e9a686c876d428e4051986abfb88ec2fcca5d8d4a6a410ce1c156daf3f96819e959784a70cf7beb068d520024281c8c82d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc700d6a0a0495c2d4818d3c952e02cf34ccae03696fdf353aeb01063d69d68a1a6afa1d6bd157e4e9d1c35aa86dfe109b3a53191a3d127cd86c1daa7db152207b6cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h115c55f415217e28ae5d81cdad93be1e9a4378957e5305f6e6572d47e9cb3962456cc1ba6d23e0c83ca1c85e90439effdbdf23a129ff368b5150ff2bd89e3240ae135;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h216d44605aeb3f82ba983e8af0789442f83dbfe698eaa13f275042b74b101705353180f72089247c766ac7f1176e0ea4da45c1fe30319c7102ba89df2e9dbfcf91bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h932b1581e6d3011587f413508e49568ea54a2922b93e074cdac32afd6e39d590057d17c264aadd1584fed02751d0acb9064b115e3e27cee2b7a27f4007ed85c9315;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120de99298a855c4de3a0c23142d5ba80d7b9a45d558de7a95e6eb03b75099cd5a26c44667d7e33eeea84fab8fa134674d3bf702b009402f0420daf534cab8b96079e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38fa7a98f17112738c7ada2d7a6fb7feb01bdcee8f66a1f5b38a89019bb7ebd300a12b81758c602faba3e5a3c626aa470980ba45528b090d84ca2146b1c1d71900d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a0644143302b8e2acdd14892c851852855c5b94ea634fb5e67d2ced6db5b59c3ad6cb76c34de21191ca996c4c7c9a72b1b6c77e45e29b9f2eb669894e35dbc8ccc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h755c02d7cd0aa9ad0663d32394370c25ba8b9594185931c63de6219dd519d60a5a3c407f5cdde48acec77d7980d51229bb192ec21e39592887701078e0bbfe8c349e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdbb1e610d1c622bf4d75c14242898d0e1bd1490d1f9de5f5a46cf810323d45103fe9ed1077268625aeba9cbac476710bde32471b173ad9f24435ea5929065f297f61;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f705b68f795ce597c1e396e0c0cc5249a05320e8e22fb43869c80f9ae9a5ef0ac6bfaf371cbd1984fe999943fd9b285314675ab0ff3a7d8c3251cf512f8fa1049b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h93fc86c17cd665c84a299869bd6ba4ec0a94c005e89bb2fa16ea88620ded4b6636299e4001089581102123b24f22cc5adf888ff244c670cf31b47698f35a27c2e898;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h184b00bbfdaf7ef6ba91566482e2ab948e55f686a7bd5476badd7e5e84a0cc76fb3a6362998668c6bb5ca6d53089de407ffbca07d22c3d1e4bbea2ddb404f79591931;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h675d0795b31354bd7853a65bcf659922ca021f41c2f10e29869077f91336e40408aac7098a3a96db67684de31acf7a853ecfb6213059806c6bec95741f108055cbe0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b19fec1da4285ea56b6f2dc3ffa254597b5259a6c501559cbe85dfcd212b5f1b1f4d4feca324c2ef7165b483aa7fbb178feae00735c1d20b807f389e61669aa1d85a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e4a3985231e3c0055f257f560d6f68e1de210edfb5f03155545a4546b6b3cfd4d5362336d5e0331ef09990691070e323b9a052d575a3b278ecd4fb99c2e86931f55a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1294e5a57c4948d76b31dae7df7fa28798cf031bf72a46d774db7905fded579ab768db917a69cddc7b7ee7006a667528d164be3bd1d0171ff7fad066d79b8ab7305d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h266e963ee31980145a4715aaea3d2db18731628ad3a425f4442397f7518747709766dad49b9fff7e8c9bd6da718aa70c88df833de48cb3cb4aac665fc5d9cbcb947a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1820ab3a3f99fb4ac12c3aed73fc29d486bfee9bf652f86cb3499ba6790f70ef479bd03642d54dfd4cc54ba8e651e36bc113aad81cdd01395458aebe4a160c721e26f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f62b4bd834eb55a338bc4673c19ad4529573a728f818fa7497270338c5cfca145ac002007caa669155204b8aaee2a48c35b076be4154848fb177f9d3571de008e168;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h177b274c185e45569bcd9efd4dc03207c7e95e6890d6b4bbaf4939cd493d86d03120f5fed7345c7331b40ce2ea7a784271d4c56586fc6e0c49222fd4e8bf5a40b341a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15ac5d75aa564e340a9aa4d78a89311b7679a244fca3e797a4e1b05da320c8ef4556d98c65470b1309d91be477d50da28fbe5238023ecc559530968afaa79ca9d787;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc41d51c8717132a7061074fd523c0e2f61cc1dd535a84a620317c4d5328322b72341ad246eea81d0f0e8d17ae173dbe19a456ddbc63c35e641cb23821b7f6655ec7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1852f8b86cc44d1d4cf81c24e3d36ff2e17660b4b92c6e9c2c74852aa3256d6b1600db9e7e039ebc6de554335c6eff7f1f4a2f5283b2ca85a4a969af85305c8892b73;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb8f9454e41aa0ece23437fce28a9e9fb392f4feaadbac326cf35a8705493c3970e55dd4ee90a482d282b114666c0884a41a314df0a0c7d208a3c95fd693ec3b2d501;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d24f948bfe0570429f6085a6c38fddc61b26d95745975d20b9c453f2790f4e7627b51b7c3fb98aa16b73f9bc68bfce24be14002452d2b62c28c80a6ee4586e4713d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15cf31ef2b1066c22290759bdf772796f70c584ec3f8fecf1475dfbad361c791d607b6c99141098b9e065fb741031fa21c57982e3b11142b356d7601ab2e453077759;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb6cd14f8af4d9769300764109121bed453034faf298848c7c3d4ead886799052f23ee558952c634ac5e8401d6de3089ae573ad77a88229e826d3333991bcc1edafeb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1089de43b2c1f7d6781a97a2c50f035f6248786ff6aa3b4cb3902ecf6fe553156762f7650c666d7068581b0624257dbde8509a0a84f27e2cef132d1abe37931a183a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h188edaf8ddbaf5fc5a634800786a593ff00bef41acb121b6f3cbdcb8b9f3571566c5ca6dd9fd9e24a8fbc8e168449cf012340bbe1db1a6212b2ef08b43ce086de4c59;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d66b9d308ebcb2187998f4d43637b364b17333680f6860905437e8efeb49f4c89fc546ade3511c64ff9ef28afe6190a66e8f543d388199454e0fefd84b8390bb0e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b6f200a249d21cec9f2a86cb20fdf679bdbf5bd112654fdb6138f3b4701a09a45e8d80b540e6a0edfcf1f88258eaf4f354f6312fec25f654d82f33f8b0d61d957ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17ba414e676e1372ae0d6ae6f1a96483237bc2253896cfc1a1a6e8c2724b60d9036c6a0c30ceccf5503a29094997b9a48c941ec5fa9e674203c3c8b4a2176d91c7e10;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h127b73681fbc7f070fb4a2331cc4bd7ae7dbc23e33b9eef3530fdeab4d635ddc060905390033cb2f5c5904daaf3ec1fd098b8a1fdfcf8422ce07ed0b2fce09e1c6509;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4910b7a1f52997711fb9df0be35d9656099d3b6e3dc5baa68ed596ab9c6344c3f9b0092e527b2af8f997d205e606cf471921f7003361042b48501e67964068360e20;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67a8918d87754a9ffe4ac3da841d95152423d5f88258ceb6f86261eab634b793cc56bc75b3b6e528d479216a5b080f24803d7268b28ae516ddb82fd77d43814def57;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15131866ee0523def8992da5547c58887d2ef8408453725b0bbc100e4b0d00a017bb914f0ee0f90f8bbca83e049881a8fe55ae422d5f549fb6ab76305fa62b46e56ea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h132a278b0a336d5971b53083c3efc72abd7f1622811a75d7b9971280d93cad1d15600d00679c96cb82103f6505188b119f17b7e1f112e07f7f69548d3ae936980391b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha805677699f68d4a8cf32d7a7907e3e4c1bff43fc120e3219f84ff92b11994d8ce34138bd5d50ee69e54aa20da818721d6f39531e8b1630c4693463a693d1888046;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8350a53a9559e79a8f54b86e42e5e3fc3538680e87980aa11f239c812efd5e84505ffa862c01d96e207d8dd94db367bae8a2ffacc57376f43a0a8fd76834f30e2bb6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c3bbe82e0484cd21dd52da4698cd588d79eda2fcbe0a290ecd57f889dd1a4e859c6e97842930d13d7859412f52921b999b0d71082ede27212cd3e1e47956528c137;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h22f07d26ce0702f45ca4779db694040660b4f7eacc88d57cfe8a9f03e2d6d4de6fe81133230a78ef2abd23a6f9bac4a82c0dee6fd461a56fcefb963a3bbd96e0eaae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab5c4166e67567bf90ac68b73d808dd22f73310571b68815e9b7799d4b48e39b0d9d8079785b5798b664167fe80da09ced96a7a3d241369aacce8ee319051727c7aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8486ac7ba8baebfe44af7e07a086b4f0c35e733b2623e25c59d79545f572838fbbf72d8800a4f2ee639b9cfb4deee9e22e437bbef3b5fa4af6383cc5a65454b97ff0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c9b9a6ce43e91f715c3366e06211029d82bf7d78e6c0e3eb94b2e70adbde3e1d9f0dda9c6ecdefcdad56f84ace98bb013536c3da5780ad7d32d5a7b93d0e30e0476;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb68f12f5fe5828849e1f00a60b904b07856bdcaab8d754cfa4dc98893b78b9e68bbb92e1a90a831eea64ebfc24ce3258a5f881cc29a5c1c002fd28b8c4539d0d2f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb66579823686e70441061a8b5b2aa627b0f0fd0aabb6aeaa3a688ff5c91b2b5e13a905d9730bb5d1fa6dfced54f7d5183a228e07637fa1177bc31480375c2f894401;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1761dd701008ee2394869220de1544aaf0c24b5df0e72f4c3235bf08ce01e3442f4c29e90a03f4d35930b2137950122ef873d11e0d179035cdeb422e234c30c4a516d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0a378afa113a823fe64a1e8445910c0137c935ce604d1e36669422beb796ac5e56176384ae2421592e77494da4e58c6352f4c2e6b3578e3b1e1f79e802ea09b7a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe0fadee881e404fd2d755e715c56c44c2305beed30cb2903145088e9c0f2b5dcec501998ce6e3e1f77837d87b5a83c962c7f481d9e92e05e54a275b683fe60df5a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h288921893f33b425f9a065597cf989394e52e8fb08b2ee5c09150dd3bff19a7899686062ee7ef49112df5bfee6f2ca44148869ae0cf8291c430fab325ccb74268883;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38b32b6046c6432befa7473af669f5392d61b3123341e828e28ca6b1b0425380f5738cc39acb0c28d31de780cefc347514ac645e7e572e9796171452b8aceffa016a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h146032ba24888e2b9480b78a1852fa7646709e6c5037b8053e740db5c345fc20b851a8bb0b6e12bd7bf8aa54de0ec958b049a0a09bcca8e8a0f43effaa3adbc98fa0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ee27630fc611e6e60166e14d402c9ae99c38b2ebe2cee0c36fce7cc052d91c4fab98d499d404948e3841f44f690c367f9b1c022f647db449a6108acb490329ea78f6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e463b38fe52c6a6a0395d3c41b1654c5aafa0824782e7f7620ccf87ab826fcf7997292915fd29cd8be54831e85a899ef080a86eceb5f02ac1b777724d4b5f6748ac4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19922414fd2c8cf72f4c4fa9bdc072defde5b92cf6c719669bb7aef37a320dae90e1e8944e7ecee70c2725124c50b260f6bd155f2a3a45aa4ec3975fb23698dfd1270;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d1749a8f5e44091b1801337a0dfbd0136837d5cb93eb8dd425f857ced66fb54f34acab83ef11d119b854220446bbe02061f9c6d05b0b4c59716e0cc8c197d1974dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h131d19ae920085f73e42c9f862300c180ff5dae67001f2267b3a79ad4eb15ce31ac7c4f039da674acc7091a271a40ee748150bbc2465b4f6284134407106d7769f023;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h173e9d63b22ed6f548a946536c49d9fd89e89f54c23bd5f2747e2c5f5c236f0d49bf848e8387e0a31e12be02098035196c25a163b9780eccb178d5241be1921092097;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd8d080d8ab69d870fc0b546040f7b52b8aa200690352680cc730ca16e1d2eb0dc0a51f90cf76935dbf4eb1d439ae7d41d0e8d3284337d312fef3f618a6e93b6a45a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb9af1111d12b8cdf9130bbaa6bb227eb293096d55156b757918f9747cf31938742e688096a51e276b05129edef2d2667a3c13153330f902a73f6505723774ddd39ee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1838f1b737a9d12b9488f4ff262e90b32570aea4d5b9eac3921422939632cc8f957887f0d4cc4a0deb2c345339aa77711106eb103fdacbe7c55e9888d02d38779d105;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1638d266e640ff43904201cfc8a5bac67addf00d5951645f82ff296363cade934da0e095a6da17ddf6a643e0c5f716713048bec8b4af2ad583a17136f0df6f9f24afe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf2eab5fe4b86656bf47370eeaf4853f88b69611a924645234412d7f9aaf4001bbfa027004c542ed015bee42bee22739f2bb9fa4c436c38c54f8f427d65c2c78880a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a265ec528c7fd5f294123284d248702fc860873a56b620a411c8a703a5d855382dce3d39e36d43b65b941606a31d18415b588dbf8a17a69b4c44fc69c097228c18c4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c822600cda2eff25e4d9f5c452ca6f464c848510162db7a9513ea82c8cf47a338617f71587388d4064e5732f0c7538add753028bc351caf646b7b0f25662efc150d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdec058b0f22a7ee1d904638b1dd64bf53d7fb0a29352520cffea1e2bd1a0795cec6119486ea55544612b642445ca7fa13d15250e2d50eb10b2c730eb27b018533e5b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bfbafbfb7d53ef6c8ca02f1c1bfaa4e3789f05f174995e08c97a8d58bd0ec7d2de52e6d91579f800c32db96c9e9f009a27ef162833c010a6e156378876be04caa41f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h125fe046631bb212f9d06855c0d347dc67a98ce70f961294745c14a3bde05cf56d7cb9531907566c4ab638d138e4fccf7231e5bb9219f6da50fb177300400e4417628;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h102301ec2ebb0aec39ed69253e3b817e8ec44afcbe8254b3cfece91767451f3a385bceb92817dbf252e74d3ed7729c5d01bfef722ea6ee87c9ba3a495b276daa87d15;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b537dad6e1bc527a5fc6526f38c67dbe8ec0329023c4f009dc5777fcb9a00f9ef3ed3ef1d80d30b00e1128879519d21e8653bb60d6e672528279ec82620573d7b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e89391b4e14e20902e24ee7adddc3913e5b5e166225ef4e96249176e9d166709aae0154993a98663eeb330c941014cfad5271d06562b3c806c32104887fb8a321072;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h50a72ff42462b424a984ab31b00ffaa6bba7b5cca6ecabd11e4be00c56e9250122358ce08a1d0544b29562ec224f9856dbf66698a31589a8b7a3acabd1a538e0033a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h95e4b844672dc433ef8e874ba2ffd60f82513d3c783e710620501b16eb8dfce423128c9897ec43d8606a0fa4781ba5098861ca5243ca8bf0ee94ee7815760421df82;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cbd9813684c6de38d3c3385a711f51f79dd26c2c3afa20d232964796e780713d9d20511c5983a78570eb9ef1f7b9d2731702bf86708e00a7f2b11236958abee09036;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7545fecec2272077b5ad050cfacab9b2b47ded17e1b6b0792c67ee9baa5913e157a3f63f31497c6d84bdd80179300b8aeb21388fd537ee4545771fa27c69ade1d257;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h20df3ad15fec5f683fec9bf21d3b733bd5523c52d2c33143e85f9fb9c08388a74385e962e68557a3b7df5fbd6368cfead527a17dc3a6c0b1caca2bf2d70414624c9d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h637b93add14e98c6f0090ecee162a49847196942a0c59c5f034fffa98822930d3d712b1cdfa71380c07a37b506aeceb02c1ad60bd6f5e394e510748e8a6816a1cdef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11309f8dd8dfca893003450574b56e6ba434a33abf983839393da520eea3021bdee858423b8d1dadd0e9701fa4d2e9d0e6c4b39ad80b9de5cdac3108880c916891555;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a09aa0b5d551effdd80d746a2fa0a0664ed91dd069e3f2d1b4a63a3b866f3ec504ce5eb3f58f549659fe29f78f38dc38882704bd3e753f0118de48cdcc28c391f475;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cb247bf8c296e1ddcdb41957875da0eccbb18c3203fd2183607044de0701e4bf002b515087458b2f498e9b632e0bae38518db0be21c749cd5f5f09d183589e8d142f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff0959e0608bee55ca08391a9dd7443b1441609060d4c5fecf3394ae2a6a8c38010625b89dd1c5dee29e85fc659236098e136385de5a29d6ced2cf4514ea3b03d99e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb791d0b172513e87a235656f7f292e6440e487d74976a8b1a4942e81d24c6a67e85f606b96af2102452d1cfbd053acd13aac0c0288c41d0c1f8ac53be09376cdfb17;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38549640e3b2f6ad502a8ed1d34d1aff01e7998dfcb1fd49c0f7a853e4ce78f40e7115b46985ec452bf6586dbc57ef4967679d4af955388538dbb29cf41ed0d86f1d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1adbd59dd828cd2bdf64834b2775ecbb3e0b315ce52f3668c021d049b6a11ac96490c51a40be390230e73ba9f266318fa892a3d57a1babbe264ea55e37155c8110523;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9410b880e5eb14407eba91fc384d0c5f27a315abe1b709ea49164380484ccba99375633753980fa944069bdac350919d5dd5ef4c54de99a5a59a4df9fe60eda94c14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165eff04696148bbb3a2362b002d8b9721fc4a62e63300fe9d87c87c19ae51bbd7089ad580133c409685be492179ef14fbe4221a7289a0a63d381d696880800c48a4c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a8ba02f38c2ea282431aed7156bade3d8a15e9cb49c81a510bc626530a0491231dfa2436f3aa65452b29c5741c2995ec499b0026e606f00993d77ba4a0e1d9450da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc80c8be6897be4dc58ad84985f8d06697fb41fae9ced3f61176226faf32510f892a241e17992182b4d2a23db105d318ec0e006a44a9007ec9177a006202bae9a947c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h123fac7cdc84a2fc483c74751e0edb7d49961951eb614abd1a27287d4bd6b776aedc69994c1ecbef4c724284610cfa0896d987ac7fab30b3fa71e5344d364816e8794;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e7ea8de7b3304e4a88fe080a3747280fc2c1acac4117cb0829b69214660e0c66f9608a7aec3f24f3736ef38ec0ff9ee3e251bf352d063142ed72bf6d1cd8391003ec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e91298aeb2f65a2ac1d9813455bd06a0b438e5a470df35ff7eeab02afdf870b62422c58634c6c2b7bba70a693f55e69364cccb773a8f1a4731308eb160a84eb5eac0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af57865fbeefce9607fb63e40f768056f664f52bde80d9889ba132d38f99167367c0b17a23ca0aed44a62a740ed960219e490ccc0ce04c42faf8a43797f008e14bae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha98d9b088f065bcecaaf3ae11657d15ddb729fd6824d7f4b632af317014ddb07231d87c94661a291d2cd6a5525fe3ad97ad55e40424c1ac210fc8d16a6f84bc97c3e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b804ba7ef7077ce0bac91273b8a0c1d8d32411b1f28bec522e7473b907a643fb19d13dc4216a6e249d0427c60ea0ffa8485d9ac0c8257540dc0f29bb993973598911;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc8b7b24a66f02a6d7032c70190994a7487968a6c91af533aa02cbee1443d1bf39d9adda02cabc48ee752fe85dfef650660838bd16586f6dd2b5c515c5ee1ff955ccc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h58292170420ad0705169cef079fc8d2f32de74fa902ee3cf59bf58788a4f3855e2eb7e19dc58cfe0845806d435323b8d2fe3ac4e2f8ceaac77a3e5364939d5184e11;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11a6c07f2aab668edf44367513052e36bcec70b9afe308bcbd69ddc7e8f716e67fa09eb32f7517190bfd926e17d4365c226edfb9af9acee995bb106613253ecca3424;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13b1867f01db5485485a053aa072ca575ebc0af871413fd9711d60a7f7dee0f239b317c92042cb6dda7605961a7492dc33240d5c4b43e9bf3faf378f2a6304e3c6738;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e46215f48a906862f3158a524ed6ac2fb69e1382dfacc54f932cccfb47c14e638dd2b9f948b0132e1826678d7ec3d0112df0b5e99cc19c9befd12203ebf68370d6c3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he15001876f8069e14cc61849c0eb03e5fb4a8c1bfd107445c45bfb36df5660e0158f8d17f197279276275bb080c369c661e69dc5da7c81264f87abd53aa3b488b284;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h82fd92d4f261ccb57b5102d0a98ba6168fc16aa1aac2bfdc85bf2f263eb47a9ddecac3bb87351ef97d1429c1f788bb58818febed7a8c0b80b69f64b462c13800f7a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha9a7d6453c3bbbf3b75fb9a11ade60f38e7786e2422f4bf2c92d6d917b029b5743bb5cb2d4cd93703448b724df380754eec22a44900d5dff1bec65d3ac53c99f7203;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha69e168535624a1ce3c820f4247ea9954da2d272e890314a79d33166574215351b074b0314952b5f9ace8cc2bd140149d7da83b9fd345a176267a09173217361ebf2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c3787ae505cd1bbe7cf59b9399cd1757133dd658d171226547995a81fce8de8679429ba536bf023a1541eb7811de2911ae7c40907fb9bfa8b4af9b56bbf112d88d19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a193c0dc01debad40b8ad715d03f1ec830b833d4f2dd8edca87260336173408f2c412198dff415866044413f38942450d499c9dcffb7fbdfa062e9bf3cf4e4eabbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11aec31217a3d930b743fa7de6eb0f656ba2e9543656aa1476d9cb60b87395dd99bd8d06fcf77fd8d0aadcb970250a39a0745093002a6b07522beb8594b78b93fd5c9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6bcb5225105aa1d7a97bad8a757ccbcd8fef38723504dd2a49f5577b06a56ba02f491b0cbac8229e8662b56f4e003118cd8f0b0c23baa7b3c31581fb5da67c6983ba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h92beda06e3347e71112425b92c88d7aad70f7c7fe9ed147a6b672752d187906d46b08cb7276761fa9932fb699c404d30f1c41899323a7871686af25891df167a4bbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h63d5cd1be0e8290b26f05f55bd72be2ee6c352b7cd314283bb05364e19d8d5d5d0a4f3d7bbdeb3930c576f25b700d40b1fd94750d5cbec5fd7e65cb4290d86065adb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13cd4eba5d5e778f972e3be97c204fb85b2245e9cfa1da80d7ea02c07564730a1382b7aed043d55b1882f7bca3f4bf114407bb250ccbab2c8764a8cf6ac4ac1f26b32;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7133180199270b574274daa04ce4209cb1e7f129897f9531e6afd8dba1cf2226877ac15d13d888157f4b5a714172e0918d14c366e0131bf6be8b793a169905dd74d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e6e8134718bb0f7d6cb0080d8da336119b54166262e3123df22d22d6ec08e03d8f5b4eb188c7d0caf240e0d90b7e2a647c12999216bba04d522e1ccdc565fbdd7f1c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d141a06fd680a2987c1096fb490b7b97a21b3da0602383fecd18db22ca34875010dc966d8b5d86664d59d8964cd9e1bc4fd0448ea9c40a1d3b83ef67d4f55d773ce7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc07d8488e5e9fd8008770f0c37259695202cb2eec819fec50747b28bcd8479750d7558706fd2a8ddb3e74febbef38800445d7db27bf515f33e40ccf392d6deb7483c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5a78b6492a5af2943b83ef7361d84b7e93f0fc685ca859508eaa2db7dbe8befd3abd6694a3f2f4c0abf4532e4907e4fade7f60969bb6acaf9f3a56f09dd2195fec1b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f46097f6023206458f9d4408a1bacedc6b52dd2427622a96f282b254eb8a98d598ede96a1a212f6e398da7d8e1c4d5fb46d34c1afcf1512d6dd84066808ff8ec9368;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11104507405e5ab7a3dfa1920882928f1cc497e595af08c9a21a8e53dfb9db6709d6398643c54af9c5c8abc8e9347e5e409cee49ed2adab44431bb35e06ce88bbbcf1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbdece0b9f8997d57a23a4f473a6cb292f853c6408cf683db726acf0a0c38bcda34c5c8f12a05b7aeb1aed71a01f7c7b6fbd3db109db134cbab0f3b3b13922b5e1c53;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h383d6d312a83b92c6c6b53a1936be07dae8906a5e6d9a2f445b690a6682da79f06470795fce774630feb219255333a27b928ee850ad175e688ccdccec48419aba2ae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha43d032f6a2916e78cfc4e043df70f9e56f5a5b4e2389dc71470d43f990235c4ca052f9b6693043ae86d7253bc3c274eb16b5d78680f51f5f86e2da8b1bc77e2bb8a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b204327a66385c90609961aa4aca1e4695f5b32931015e04ca4650e8445abe8302b36fe10d5c425540577c8c72c769d192b5711a17b45d9deb0fe91f7e809c18b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dd66e8665e71f6896600bdd85b12c860f7583955ab5a7cc323ceb7827c648f02a1b353bf313dd4efd4fd88491d52a63e65349a8727fabe69a2f8b45b3eb015e3a0c3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ec0e6da49b05d9ddd6ec3bac903bb9061d06e8456869f11ddfd96fd2b5de3a2e8f1dfe02865cababc231a264d99049d8aba3540a2514aa72dfa28791149c82bf6300;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h170baedd9cd3bb6ee55e48d639f00ea88fef5b6929d3e08c1e47e9ab8ef2a5c746d561fe59ce5e306e0fad103fc3592bfb766a8928c64851b27190906cc3e8adb980b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dcce1e0dbc74bf93ab190c0368cb46277e61a732c7e4aa65730e3bf98b8dbcdf6ad1fef88f9b27e108542e2773c3d2dd7a4044e4dbc5f9af1b4b3ace350358d8da61;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hebed94da3dd6435a78b927241ef368a4ca83e9d0db4730f981b568a54136b0e466840c0d19b800b7f60b31d9b41a3517a0157245898d6d57490b1e0feb03686f49c4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105f955d785ddee6c9ee9d847c9289164ec85bc3295d6089c8df133d1135e94c5ac1c5d7a30fb1c1acc63b222f3ed74ea5c46e11e8b216c6009dbe5fe4c3c5d0ed381;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105a462d0851e38243ed3b75b17abb701e14ddcdd1b85e697cec4cb086f6b30efec06974402f47fa022e38e3f1913c8861025d9e76d151cc82746725e39e5d0673cf6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d5a8de8c199d69ac7ed1076354aa1608b6f2a3bc399610f09f54aee8555a20bbede444fad65a868a580af91caf2bcf352cecb3d06efca52302c453cd0286db5a5c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hebf04c82d58a17a9052d4c42f1fa9bd6d15da12501e2c90aa0a95fcd970f664e2929dee2aa82026b70253e7775b2f4ece5b3aec66fa202859162d0582a4fc96f1a59;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3683d06da8b2ff2243349d5d899b4f790c2755c74d9b8b348a26d4d36929cba8e0fa7c8f9261d223aeee541f94878762bb2bd88c496db66cd669ad56bf79fde9ff41;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14c878537a975c1894cd3387bc43bc51e6f144ca38585e4a644cda0c5c28a923d46465682464180c7d8f10ba39c377a7b50374cd490eecfb8a26bd5ec4d9dcab62a56;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129422bb44a326b828ab1926447c857d536586b28a174e0efca65d10a74c0f663654855dccc36c848df87e2dae5372c21184019c2f0fd1cea537f85a8df05a9e35947;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c909ff8d1b48029a7de8f03369660bf3198774db0951075197e9b171d1d5200e120a0ba577436f2ece1e7c0e42a80598a891ae47343c1b109c85daa2709e66fb793f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1be3cda0dd0d22d787dde28bd01176240323cb8be9ccad5631862f3f765d9ad504461f0e98bb2746123ec84f322f3b4fb7f0b7ffad5551857b12ddeb77dbad1133c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1369348aef2927be4414eac8616c9915a67acb65ce4450943c7ce56799fd3f463c63432df6972254726302f9e4807b12139c21166aa573987021f2d830241ec57fcae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8013bb5e3dbbf208c880b90b61abef46aa3c5aa45aadab1df14188b6077b2d428d1644ab8c78737f2389e3be0dd4c7df3b5ea358eb3c294500786d43a95c7aea6f11;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd2e44c8c0e917c2c3a7c63d2c32d26796e467707c6df26eb8e70416ec77e735acc0e5f86d3aa51ed22cdfb064a63a86142eee354c0d9d049f94697bd22a2d1011ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9fd84a6450430e755103e6a1996b242a3baf5ecb0cec59d061c52bc5234953d9eca996a1b04e736e4660f0aa5827ccc9e9946b56180ba311eb666e8e00975b05fda;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf793bb0fab7eecccb97663ef553f6eb9cba441422a60a353d483de5133b2de26a3509d84c474e39b167cca48d493400b034768cd62bf27dc8431312e9fbe12be5015;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19039637f4ebd3f9c1efc67c66a1fc6379363c00332b7fd7446484af204ec5c68629e1c045205687e959a715025677d4daf8e08f03d3852b8df3e3b3d575a414cbd82;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c21d826f120db3799094e51567cac00947e17db83680d98bf135d281bda4cc9215843576ee4a3d2732c943d799aa2d80f4161e1d518f794e35b605dc8c7de13507e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97680a0c70345edacb37c04ac4a6b6f2c4aa53eb08a772b856d0554884bdcb813769b20f75fb92babfda57eb2e0507c40a8d334873f1c187077ff27e592df4aabec4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b0c6ccc77a102c5564f9db3982f7d07a440b39eeda828b960c4bd5a67473b3c0d3aeb4a6234e6032f91471bf366d9ed9537e4ddeda0c424fb116090daff357b0718a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6751ce517f1bdd3ea0b5774c52d6ed5042bfd804555a1970c81a8eb51e8f3a9e2b733bdf9213c518f17c2a0e86d968894434e720917e9e092f16f2ef894dbcb7e5ea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd328ac07381d2277b5ab41bb9539141df056f0a5e4b0da0ea0466a8e6ba54824747b862513f8dd79c2d68366941741f3ecedddbb3fd3252fa0e99fa52acae0d40a79;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdf5d8719985f44931073ea1a7215ce8b6f3192cdc73118eed1d2fafcbdc1110afd4de95c8bf8de053107e3ffd4565cdd3c7df42e82329094b788b55610fece55152d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13248f0f4f185f87fecad25af3f3e5597045b3358a77339027ee5caf5229a78b009938c6fef8d8f9c444783f372dea24b946d969a99964106310416d5cde07dbefef5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa431557587cab4ba3d612b8aeaf9b47eb56e9a5aa21c10ee097faff6d43a2296797d1b4ad482b787ef0f1696c0d9c3220db1e6febfe5c1550361ba8a619e6545bf4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb9fa7c5afca5fd9988437142d791c61041c9cad659d27787a0f3496883da1ab3882e9a2a6fc5d3e92afa5d2a5322a61a1d703255ee65d1b6e308a0f25111a7aee8c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5906592b4103eacaf4f009f4f36e4fde22c1434d48a881cc5852b699e78eb46e8af7538a938dcce5811619225233e0da8fda10d6fc1e64a6e793fb5513363edd980;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2a66295110cbe7a25acf78e968cbe87be34ed19e0561fc53e681e067586938eb2d5dd018560045d118a98997c9d77f39dbabe1b0872e9430070679ea4143cad37f3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3dea47e173cbda7b703b948a21a3e845040693577bc4a0136a6649d5ed01b7535cbb77edb7ddf19d47c9a175c8a9d1e0f24859e265d5885a0e616fb9e5684cd7129;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c60792088b3ed2929d53db156d6579ca7fc0e3f9c505e1a962bdd544f806a9acd7ae0647b4c504f96e401565c91c43985a1137e7fe6433258e0ac5de16a2edfeaa63;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ccb5c02e4c6fddd29b5fb3f64ff1ac81e559f72a480c189236928dbb43a057a87a4b3c795d7613d42423bba8ba8299d56f47034abf00f7f3a3f27d6b86ca6d455039;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eda842b9754a57e1582c5743f9d0917a56fd1c247688daf4786979a7206b134de23e12d8db290f4b667387ef1afd840ce2b6bfb2ea333999eccfd3db6b19fe89d3ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12da09562e1896b9ac8bac11bf9bd210012fe5c9471488d17586d8e309f3512a36700c47c077fc63660666e87150a681d504fddf0e03da1dcc10cd068fbc9558e03a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1304796dace923e30c99ddb132e2306e99aed338d74ae96de6346b5769d127dbcf2c4a974ec5962e488a900478b5c9203408dbf5040fd0011313aa1da7d23c070851a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24e6315fb0a06a828cc1a76c093016ec5a8061b8fcbb4a6b637746aabf4ca34629d1571b5dcfde631a9d13489b5f633f51df0da32442b4f7727811c583b6d1d5139b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed0c258b0165084763ddb3bd015b6eff0d89a35a6e70d7f1c394a298e50b97409c5e771b30c44364f8ff219d2664199f992757869288089504ff1e8f979f3cea2de1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1baceefa9ae0361d567a8ce4958c9822a11ada87e0b64c4f19a6fb8782e45b4e6c336ff75257fa7e744815ddb2275b5900c538d14978a6c36f584cf3c80108aa4ea71;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he588fe5664fb87fcb32b824911ee2d02f64b131241c64310e5cb632a18376c263fc62b57734f30d35aa6fc7488e94b9450afede856f3cff5aad9e7c47db6fd9c076f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69cd5b3e75d9d4ec620a06c87b460cabb82217a1890ff8489db1ac486f95e35a39d2503b6728d96e934422ad0290e680fff50a547e850909997d71e0727dca11df8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5041d3ffde55643ebb9a0c4815b1e94ca05d4221af535c2ca3da3a5c881945989ea2f7f788ed3c727d1bfda249199effe96841fece3ee0e3ad810ea72bea53359c42;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfdf06cc11163a275542a16c6a595e195f4123192f6316e4ac4ba321d073a33b7cdbaf6c82a73edd291fdfbb8256437a0399c2667e1585267fea3c915fbc6dd40669;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h185ca971c5c5b450a4136383738fbb1772ba30199b191ca4faeb2eb762112ca0048e0a2df8546563358ed32d23862a13af5b61558375a62ca11660ae11eaa7366a51f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12ccf76883f4376fa5c9ef53a33d3392ea906ed13881e0d7ac143f8451cfdb2123d982fbeab7a9a54ec53bd4e83401d1a256ad6162eafb175f8e14178cebe5c7006fb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1edf45343973384d66149bcbaebb2097856eed10d80dac07e638c4054e3f117c3c45153304db0b075c466fd6b9d946da45d97de161d610d87e0b3b84dd7429053f321;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a11ef77233ceab3c14108c9eba8efcbed32a4919fd41b5b43d42e1a3f7e7ccf865905b26fb74f80b03ce0751005a79150edbc11ae57abb513ba0810e30a0702fc582;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a11eef2f36ce5993ef9df80c23dde0d3147d9db551079aca6215d7b39c5390f5790bed5057e4c79577b2c645b3d0b89e7a8101655901eae04c0b38da14368e1fa562;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10151d993dd920706700c3f565bb3f3c40f1f6e0958340aeff8d4dd0445b7abab8eb96a7a1d8f2d5b35d835618efb5bd78c5b4b60ca23808f999939016d11891c1443;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f6a3a41658fc1cf967b5dc120221d85b4204ebb7be058b347e39465cb2d9a70840e0ac9520879ab7205d3aea48feb5cd3b68920925a611ceb377b7d023c54f32a4e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bc2d87c7101f8b12b5fd0236ddb59a11f6cae3f2463aa93374713ca9e3d5d612806b3a28d1509de9c2bcaeb4e590571dc36a2dcbb268e0a5dbdd24e0064461a440dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15afbce09ec9777c0934c6c3b88d12f05830707c6dafb0f572282a6e91a83457cfb142279ddb87e95451af01ea60fd44ccf7e5ca79b83fd1077425b8660bc9787cefc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a98be75c0e0c688ec0413121991312b80263b529f797e1f17a67fd7b801411ffd60110dd88fa72e64d3e4ed2cdf67d446a15e06f3a2c3ff7556cd754bf1b2e1bb666;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h26d3871bc23dbe034131d52f7429c4be46449fe123ed26dd775d0bf449c325a51e32e27f8d8f1e25a8fdde9389d4e9e72cc53fe6feb5b748d20e5d5049737b8775f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1704ef5b8a781f34f66a04768d84c4eef50b42cd175230b46f6d35df68b04246679828521439f992800a71c2d47a6ca92343e9408418fdec184e6f31c0bcb425ac63f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a2f6466e519a9bcfe721e4db6440578d91a38259d7df690429595c57d92d7fe7ebad4208ddb8c19d8aa2af8c0e27783b1dc4941fe907ee91797e2b6a1e34f395459;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11a85ae137df88e51ca56428bd07548c975bbb57845ef6f7893efd5f71eeacb5cebb7a258217e566541cf9cbb2f68a0705d83ffca6fc5d5362b0a190d8764bc02e536;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ba94293a6d3c6ad4cb03ce7b46fb198abc6b7211b027164084b4e5a11c7960409192c1abf2d901cdbbfe28144c857cfb4dbe21975a7391a6529de985faee5dca5e3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1debfe25b9e80a9fe712d5e89aadc52033458cfba2d37714ee566f1ab46cba7c36c3d09a1d0e8b50be3e2b13f8df432594eed9ccc0bdd47928b2d95671d5aec1c3049;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10071a9b6f14d3f72ee5b5bf80d01107e0ee266604037d821f5c1e765cb50d8ee51b8b125caf9e7f65fc6e4f5e311790027784d24cd29d5a1260b0c9ff3488332159;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hefc9b66e5700a96b4b85f5ae0de9a08e94b453c863cfc22cd343733a7f36b29539d724ad43282ed4c4ba8c89980008cd41c869eef4f45c2e01de17e773ac074c31b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b702f3767dd427960e0f2d357d55d217e963bde5d62e99aee90f8e9daf1f596a790ecc29b146aadf28bb0ed82f5a765042c143b768137dd4f32166c7ff4976cae07;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcb92a9ec1310a2663cb680158d4e4253ce4bb944de3d73e10231451a952a1d40317bf07449f226eaa366bb2e25b371d51d45c8e5c3f0e3c2d32421e9d9806b7332fc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he7decf28340b828377232a8f0fe2aeb74e0c14f7baa5ed329be7492a581b0217ee62dd26757e3efabbb3f220e9f0e3115da11401b0e5480e22adbb20c3f961e3ae39;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120038e72ea7b2fb40b073782e9eb548bb73b0805f8b3f7c67ffd0d75474c9860f0ae8e3d9cc0e16d53601aba979e88528ff29b2177f3bea1ecb9137cdd8515008b7a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14e5ce7cb3bd532fb6eed5093c4572e64d588d225ecffd7a8e42a613278daf7fb4f40b428870e3c840237a460b0b22bc704c617867808bb09e84d5880357714e22e46;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hda8f0938a0acb5d18ec303b7d6da719da617e735b5b0e22fd2402cad6544e53cd39fbb9b2c3d28cf5e246c4064af864f731bc36318c42f94b44ca890e42b470ce0fc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18025392113de2a259e6c224fd2ee21bae8bc8c29d895370d3dcce7fae28226cd9ee9dd0d1b4b5c49a82889bbc4db400b9b43d6f2bfb93812e66010127e561d2a5c8e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb11955177c28bf6b8dc2ad4087a095618b1f342b56b9b336fec8ff2ae95f26c0e994ae31376f2af18f4025fac31d229871cfeefe04ed358694ac635185b41eb8753;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69ee011f8070fc631868060c1e867330b439373cc85c677792a010620a330da525997e790947ccaba2fb41dec1fbdcaf24b988857a271fc4b63ec5fcf5e6f38e2c25;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1916a1c29bd4bbe696661211f67fc19005ffed5364d569f8b226064e07fccbd145036ff02af6f5edf47a15c3ab646c97234ba564c5df8fa7523bde29c02c7a44fccb3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60442951226918152bdc18f6f96a06d58f757b0762b5451d50dcddc341f9f305784976577d9a4401e67570e334c6f5cebecfef66a01c36c248fb7486256bbbd6d63f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80cbc310b27d63e71d6ee4be040e87f988e54458c5610a083d6120ae33d93faa69e5d159402af28f38ca21bc1a5e2d51e3b415e02e14c45d89828c4f5218244b17b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha1c56a2abf6d71ed556f2d1d6765ad0c08ecef5add7ac2b0d97887add6c8fe6146005150ab2c1b33d8516c19c2f63e0c230fc5d4c443e8c14e971959d215ceafbccf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13ad28b89f26686d667bef4d696e6f4a1c8918cd7fa7a9614a2b320155ca73f2c7f901f7e8dbbbb3d3c894d8126ee8ecd761ac57221ddd9584c61c7d5dd47edd382ba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h85f451b4694f611873f3ce39c021c9355eed0ef735c21cdf92193daf1f0a6c3053901f6116aecb5f7b351cbffab03e8c288cbb860273bd22d88932f061ea932014ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb36a0ba0ede7ba8d6ee82bd5bd8cbd834536046773762585ef6a484cdb86758b44f20ef8eddc25f12c9bbfc3f62f71d3338b77b19da93254fa54b7d521ab2e81c405;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16158543a6dd0f83869afa7af31fb24263612f302f235bb961abfe118eb541f629044205f8d0adf35c362a254feea604fae1ddde332be58f06cf133f8959f42019b1c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha59d0fa8887b2e8e0cc5730abdca48ceed364f34b7c34599d820ee1c4cb383fa8a19ed2d2a74d14fbe12ef2ebcba691f61a20e859ac9271d773bc71422e59300cc62;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h148f058562b8f1ddd9ba0fbb3352cbc424bf136f0bed58ce65585357babd3bf8ebe58b20ad85d4f4e3264ccf658eb39cd7506acbd6c125055b40933f5209aabcd8838;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71d82f0d7db5e4e42c1d10bbcf70d859cd14b03ca12eac81ad63b392fe0ecb79f01f0b3b6d7238d3f4d3d245ad8790797d67185636eab482224d649317a3e158fffd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb1e78e638a9dd639d228c09921087b19bc2a41c64b9fa4d4f59c5e772a3fc0ddadfd67ca3785f0fe00dcd88040a7c6eb67ad3b50e2123531834147dbf9df4dc9ce2a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e3c56ef3e5b8bb2a703516b6ffce524cca2a2f0af1171683c29c9ad4c6154b215e132ccd4168a132bb12a4321e6477363073ddc0a1bae8057acefc792c96d8d37a5a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1598976eb2b32f013363ddfce492700f9f299bc717783b985ccffa1cceb8f8c70e04afd3b4b4b17a50f47efbfaf3254581431775d380e6c40bc6b6e192a62336ecb56;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5636a2c49a87f8a056e2ed87a2f0a711b9c45f6d9d270ad2c7db3ce759dca74c8ecba5af287d24fc069ce8ad88b142c54c3b3a4c042beadd435b7ed1f1e7f20fd2aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b00e9e7e0152f46b5a09cdefad90924f8fca105ecaa56418090573ba87996190109f8676b0afc9f378e83ff80e679cb84b8c0efa5d831d13bd6ebc3ea0755aa31063;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3d0e8d3d3b84e02c9c6c936a12961a2da7678709e66830aea03a5e7b1232187a5bc39f664110303450448f4e4e87b107494ea4c6a48e06fc31857d8ba211743cd520;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91d10839af76df9f46dbd1e6b9420c5148d1acfbfa17f26402dae0bc35e3c7b7d33c5c259e02f83ed9a1db89aba5cc93b044fa121013a36a560a1f2b4c894ab5b28b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa7091c8ac3084800de192efb2b797bee5ecffb615886ca94c08910b743c7d03d81faf72d067cbb6fbc453709b6e42e533ce1cacd1dd8d7dfa813139ab4fadd0f96c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ec35563dcee34c500fc1b234803b54792f185582ddf2079384b37aae4d3bd0cc0d47bdd21cfabb2b0ee6619e4563ae67ec44f8fe8b7d0c5735be9ac4096fec1fb374;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h166d56ee1073c62daeb2ee208f14de8471c8b38289a6e232c6263ade34575a90f61c793cfe96d56764cc2e88ae5dc33a726f72e79adedc9b80af9465512ed6ab67ff5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h177105633fc2560b1c4b1baa73a57ae8ad8e05522fc44dfc4fb83ca982cc65975cbf608c7c504ec8e9f0d3833c3b7ba8821bfe5410931461f5da22f698dc5de2492a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc1fca74fe9519a2d9ed6fd39ac8fcdd313ec2bba7026738c1cc017d49912df3bbe23812e0c28681c404550e41e66fd94689575ab0512c07e880eeeb7ad68b6075ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd77c20588679a4c0dff8745d2dc1a3b87af7b3ab414db8122ae97d0eba80b8ecd1ccb420200d2669d1de9cd6bdc03e2d13f042548acee7b04b26a59accf489c88beb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1529d4d59d87691ef228e3b3ab56d49e8c08e3112436e30239a3db6366e8d9572e8389bc5fac1d5b74b21024ac98a568fa11650c2125a376454bc4561c8761f16a64a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1db07415f03c5f368be3d28c04a0cf2643feda4da230247c52acf61b8eb8341b05c22ec54a409717fedc71e38cfac7dd401216eef79b43a360c15b28cffc6720d3b6e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h192473eaf82f26cdfbd9e03d888954716d5dc092d51a51021944f6f9f5b9c5762b5cb858e80c8fb77f41c0fe169ecdff8008f80756994f6c6b564edc6346cfc99e1e3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f29bd44e646208445002a79401ac3e645b7a7b296d7ad516045f61dbc6e36e4aa599c3b2217ddc4974660a582f9f0a6eae095db62049e86fbaa5d6df7dce5f62f9b6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ced8988bd942fe36ca1bd773e5c73191a666ae2244a849df2335e3f6f2004ed6c9aead948d4d789c7aa32cea03c02a4da4d7f4372ccea3afa056d2ec2c6443dbd2b1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4ccdddb7f0b04514c045afed71287474f19ab5c972c09f47b9ac676c6d9b7628eb1368474ba77d3449ee3f328b80d7d1ebe8eb50732c66d08ef61cd4c7441c642444;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1120e98c9379c9b7d0817f28cd7b0f4d778a26f2c76be8b9ba3055cf2311a3b86076848b733ce6dadcba45b47f9001adc1cbfb6ebffa87b6b1fddaa4163bbf22eb695;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11610edde43423d0cfe20aabb46160403a534d3c43c8592c8f91e7fa8b382b62bad9b412d0c66f4a51172d74581368b34c5c96641e804d08b0e124a18460af2e92621;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h148467b70aeac2620ede8fcb8326c1357a62bf1e7b26018987d124e195d1cd93e1eb6f3bfc9f9ff9b5df4dcfcaa81ad5c8735d3b19df3efedf67494811b3fca318509;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c33f12d7bafe3809dfbd7b7d2a495870ae95feb126572d3a07afb0b11730a78dcc8fbfe94852812c3149f9728f2fc8ea712cb63c35f1f5e331cf96003eec17ed5aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b5b82c9b4d93612305da2f17a9038c820ea67d29280e9791c7d7dcbc2392e76ef458903041e7349742714542abdba113f8b939c4f24d4d94fd24046131efa28cc783;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3cf21131be958502b7f1ac0f3d86b36f46ffa2b90bfcc06c60f9ac34efb9c3d2a4b778b9a82d775b873aa88b6fa269f6f7f57b719c957e09804826d2019e3ca8a4b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d8620a27cc3925163bfc9b2d61266eafd877c333e074993f9a58f5cab9f62a1c0e122cf830b1c5bf0ab5f602b9892f6e11ec37e87f5077934332d1b05ab38d6075b0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc7054b63314ebde35bf53dd7131348c606dd146355af9fcd7f15cb7ea10bd58c98921b82063ea85891dec30e498dbddfc43a518991d33473ee539dbb1cc573b049b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h640ea4735fbaac06db2e768031c78a41d79d0574fc56d31a5698657cd079039267ac8d662ed1675a94a483e333201e7d938be2dd60645fd29fc19d455eba139ece74;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca9e78ea7a6d8624d51de2949e3eefcb8e9152fbe29b14328a7395955f329141ce1372e18cb4dba26028cb84ae47c3d909f4e7fdc35a5b3e2949f753b0121b514105;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f8d954aa2124cf4bfccb353e7efb4e8ec9f05e261d3d03043cafb8525ea62c04a78e57320713676b6c0ae17e63453be1a6d920a4860d7ff38ebcca56eaf85bb41a7c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53d99d89d8130962550ef8278437003b4125cb010eca1a68e366954003abc67adce727258af074e77307a4fd2d225402f9264b5f0c6424bd2fc83e9f9b60a2ed10cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14f266e1e874e3ae2c92034d47144b85c14783ec472dbce2771f2ab382de36c927daece6a4acb25c53cea0918c505ec857a6bd30a56982e5157093d0e76e8c0dfc2b5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h478fa5d600cab9d4fb3cde535c3a332967a334e24ff807ec6c835532355007924922dcc9b2e438425adb4c08ba5ffe9b25dadfd05d9d6aaf86cc00e8b20cdbfed89d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14c99145588183f1f0586ecbc80e540c08a056b7979c639472a539ca792f9c2646062e6c2d62825149adad7578922a1c41dddad04658c613d84a8f41be4e3dcf32cc7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf75446d8dd2dcc8bf17b7ccd93f9703edece9f0e17321f89a40527d4d449ed5b51028540d66e83b37fd798bbb9c4f96482442e4661e50f50443ac7eab8391368fc80;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd39a5ed4184d798b2c16b9e6d4e898c7f301b413a9c0fbd8cb2ec9bf92af1b27557584134032832b29b689d91dbb94a560e3ef7d6137b801b485d455f58094b2530;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1263cf1754d57372497d575a094a81bb4bbf1429a0e6d35dc59711745227714077903abba835259c55c3596839e0b773e53781b920b84ecd6ee94eb406e59e0806903;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150af5b81ae26c07df93ccc06cc321ae864f36e19e99848080562e71ef01e3691c01af0e844dd3ce7b9474e102fe72e8b3fb86ce21a02327160f45d93fe5037c69b69;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb4e87674e36e5bef0b4ac2412e8d59269f1aeda933e7456821aeefe498937717e7935c9ab5366c1d2836487713281735949320d66ca449a9c88b41dd1426acf2f298;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1efefe782c8010f4c2056aa0b2900f224f7a053bf01f5264bc47447fddfebe5818ce16c2227d30a6767c7b9846787ad2caf56f44c114e864af8871c6421b81a261d61;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c2f4ada55523292a0e62d2ddfb747a9f2a6c5c0b34688c1cf5c1c8b8002e5c528ec2f0a41a325566ec45623b35f76bb5178a92fcd65b6c0b32fff510f35f8ffdf99;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24565f5b06284230cc18daae65cfa1c70b4a7828290f3e2d0f561fedfbdaa54dbbe9921a54db934bac2c0583db3add28325f2a40966dab1635a2cd26403555c3a290;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6a56b961ecb70498d08648e27674e2bb2b287997af9b5fe5468fd5cb2017aee16dacf955f88b196ecff52fa2482849fb1b12bf922ad698d3c25654b971ba1a83168;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19736e9d0016a2a9fb734896dc8d7d656a93a3377ee85e9e48723f126c9b6489fdcee2d9535693a77d2393952e68ace5d46007ffce0e6f78cd6ce516e121c92b1deeb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12390e649cc36f751e94efdcfee8aefc966b710b57822a0897c685836fcfec16becd688ec747347766e1dd82873cd110e8522a94160706248c6fe728acd1b98405987;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3308b214d5aed20480cde0f2e17c6c96b96562fd4553c68a60a2d9c88a3998f3ba7214af573ce0e04e0a8626c7db014033bd681edb06fb52f3412d8ecd6d59a03a3b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9681abe63fdd5f2af602f4eed0d6437f849469992840bd6378a0f48fd1145cc5b0bd6a685f5ad789568340cd18f37804944c4093d301f64031d0361156aa644d5531;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha1d3111dc77552e082a4694267ac854db47021c2f3b60174082471dde9970889b2f36a549dac21843d3ac5f1e5f514451804e31f7229c9a0102e18cadb700d0044d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a952372049bb31cca4da2902e327d85b50c1cf709027ac290cdb311b408184269d537229b51336c3cfd2566068bceb1cadd713f38d46b6e3f58594cb74f09fc3086;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1439a9c3e8a817b8d02c1adc2db4a99e3aeda7b894e9eb1374d3aabd57d50673113b7288983e87486eb66d389f88588b29e03ceeefcbbad0ef8b5bdb6902610e96f61;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h111bc65fa48291303f8b39ef935905d7bb5ee9bf13421df62e404a52993caddf095a4995087ee0fa1812c8d67e83fecfa65adbccc3ae643fb69bbc05b919579b2f508;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea37cd7befb8e4716c8ed65b46732c685781b83911914c373a5fc344c823830441ef7a684f5053ac4cdd0a75b2268d781d0faec43240d3d31a18daed8bcc9a77b3ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h192e1475818f7661a776ad6eddb4a8bd03fa2a73d11c08eaf94b605bf32b55e5996adbca6e8b9784ab0d4da61bb30938ecd03ec52925e7cbb776c20228808f6661129;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d7ba20f1d8f9d51bba9017fd839f680d57e81c5ef24e31f8a8149a790f0866d3238f15a23caf4d49c0ff4fd340f51df0ead2a7931a2cbe200a04e46ff4fda3dbe36;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1167863b748dd8347f9afedc24986c65ebd405d22d42c521b66695c5f5d68bec851e0586adfea591f26ffeeadf87475f5b4f333f48fefa36840c5837c02979884320b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13114280b3cc9cbfe7500cfebff147b5b3ad1aaa44dd6a1237ed8f4b16b383e739f7f5e489beb043486e7ac179ba3e71545273704b0ffdb13ac8b07d5f2dc88a08d18;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c9f5114c620b2e2a521cc90365af8ec3282953405bf9adf6f1e0b960c368135d3ddfc25c20d381953ec1886603b58ff924be9660a44d5a293d4eac7738aefe0f69a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15308effd6783346cd02acc957d0319e94c54759ba6371cd4bbd90b676466982c0ae722c9c46dea610baa1744d096cb9df2bb00ade065d13bac99c312157a3afa37df;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a48c76bb650d437c19eb7a696a339c9c795c3bd8ffa96f2dece7627315ff94d945cf443d31de954b518523cbeaa54c976d64d32a3e6aac4cb18e42f9adbdd581281;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h72903cf49eff5fb57dab3c1f4d13086b16fb8ad6fe9d4f0da45a41ecc08e288bf23e7dca1b121355e79bce77342125056a348ac392fe02445aef44d4e576a3e76d5a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc05ee13a49b401b32b06f9a7bf86823f704bc6779ce7f299d93e76768aad943c30f7a6ffde6692f933d2e8b0d96dc8013a73ec465e4f41436c61e24e1124a987d4dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ecfc640fd9802850a6341ca203be445689a60f6008d6def4acf45df2c031c1da1b33b6554167bd1cb42e1f222e0fa745f063c20094d78490ab175717d06b8279938;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1812679f02df18fb7215f20d023e312ce95dc1bab9d8fcb952d28280b1eb323809599c64ead7d61e1d95f238084f3a270df7782c1b40f78a39b1120922cac43cc9cde;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b35b21e78d4086166dd88558c8f5a5e2cec678a57c13cf80b4e43e355150da6f88bed59a14587427c5fb74d50dfda80b9b48d7acdd0935cdfba62e8ded17854c394;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9264e52249d1a8c7cfd04bf4680fe84f3bf5490f645e90c4c100c2f13ea9247fe8b66d14a1be238241ead9fa64693853ec8e75576c0db90800e7de8fcfa46635e7d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f0390130d6511e8b932774674c2aedb37d5191b55843c017e2b7d2004c41df2b0efd724ed1f1005816c701b22bd2b9b06315e45d18ee5976c96496f757d9c8d9c3e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcacdec49c3ee65ef34172132b7cf4d194740e4dc59183111c2ba6a38c36e855cdaa0237028a3c8698696cb5582901edb18977111ff387da07765090dabbabf7c3626;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf73f2d1dc02b08c7095033e464ab398ad7a7bb2c16b98173edc1c195d8c0ffda911f8505839ef7b85faef152039d6a614cc9ee2ac18459d77a3efeb73ecc82b489e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h125a31a4c3bdf7b394bc286d553e34f84d433bb28537d60421f11e29a49c338ee51d0054738d130d19dad26af8368e6fbe76409327aaa5fc4fddea2a98f8d7e9dd2bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89da6d681995e90cfa32a8c1fe6352c7615a4336d165e3b28fab616beed62fa7b915deaa7fe889f7d66b4fb5ac98f5e0161f4defc5cd36b655b63e92f528e1587ed7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc64eb40baebc7b65464a2182d01eb28b301883f2cc6c71a0f1a5c24156dce21631cef7e30e1be8b596ab93e499da35d3323a225f99003b98261eb5139bf05a50560;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde3cc7414abef1ca5b670dc899c2e2d55b1b97b03eebb5ae8f4478a83e5951ee1867785b9ac4400ec79abec14ea7890ac1ceb30e71ecefedcdcd2e792e0c0a6b08f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2a76107cdd6495c5c0213b6b7eb34e4356244b1a3a3e00a353640ea5dfe8bbc29b12e216563597eb79f287789ffd552dac2d838fc6d69e1d45351b4013776983ef67;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c33ae8d0de617919b48ad21de7b063013a80b848feca36dd5144edcbc3c6df8395e2d9bc02f506f6827a34c12a3c17e95c677f18681f1ff7aee3dd536ce08e61ceee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190577420c8032b838ab3cd2ac721680426a7087381159eae2bfdd45bbe2073b35d364f92e2c1ff9792412da0d63d211fdb2149c36bbf3cdfacef3c94f0367096bf44;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ea3279bb5a9abc34f52457abb68bacaa6d74f7aaf68de655ff4018abbdc3e57b51804dc1c7595868a623ad32415a97e50680d14c451561a7d73309bd671b67d45cc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a64ac7ed52baed20ffd236d8bdc462129c863279a68256724f4e1396cf6e2f41af17a16f718a8607055ae153746943f4d18813c48be51a825cc6f194d6fa8c8323d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c51f814d5f73e7e4a5213b379fcdca4d27a60f39e400db1ef5e881ac637a235063f5c0f7d7ad86dbbcb672365a6b5d3676027f753e12dcab8a84215c12ca93291cb9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121aa968f3e224ae1433511883fefedf04804e1247994e49048a1da7a7aeb440f0e786457aa594686b584d590cf08d87d5dc36fb9f722bd363656532dad4e25151d7d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9969a47427981770f6e3cde9f97db6f76165e483daa67513eb4d120eb852e02dac7df6a37fe53363eeb6a58fd7d773547a6531dd7d25f38bb6effa279b13265f4e67;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14f18bc7e19fecb0a4ae33e37c79891125aef466a7813beb3624881b5f9bb8315278ac2dec5fcbf345f5436e57959ea1ad5b9be6a97b8cf3cfa188a6a0ea4ee205f4f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hec09aef45c5adc4a13bf49d4c374f22dcf769dda1a724029abbf763e6b21b74464779f12a7c8ae852ea980531c31a1a3ae342fbb42da2f415c1df8a85c6e0ff85b89;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6bedb698d78d906289e28a6acdc75319d5806e3dab20aec6042383584ebf142e53239dfc44002530f31fde4b1b6a0b4302bdabb2ef0a312640448ae179f54a849d85;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9a9e267486b6d2d3320592af5edce787c7f44c1252c09353ecc73d0158b91d81d4c929805f6d87c7ea163e1170324d9343bd5a2a800c76d3c1b3a3eee51f33f261a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h111cc4a7699512130f1ae933d4f9c21e2212f4f5b9b4ef98ad4efdb03c25037c6799652e9e450230c35cf6c46dbd08ade3fdaf1c3d2cda51946cfb1241568493a95f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e6c279843c113beedd3518d89b342135395db7d3052ce98aeb6b8bc1c4b8a53c8c3ad6a037cc473cc83c3a518086c76bd404e6bb5c549930a6bb196475ac0fb8803;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac48b41c0578948ce487d90fbff8e99bc5b0436850ecad8df15c2f6f0052caa86b5c07cff0c672f94efa5232fff38b35952fbb851f897c510ce9a42efc87701985d3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17fac984ac08c6aa4707f5697f03b1f0e718a9f9f25e55ac1e37bf027c796f80fafc009697a400bf55ab473f07392712199cebeaae2055a242237a234028e1d55ca3f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d35fc7e0f479fa54f0a36ca69f65ca5722394aafaf1b1fdda1e57080e55180b3ac967ebdaf8e208312ba838243022b1c23a4f8aa8e4257558f68492a99d4e69858e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he14314ddee6522e8a9fee2322e0e4c6b42b0acfc73bf7efb17ab19fe0821c1d683de1e5c34c1be70f6cb14e64da0bb66aa811ef77b8f5d160ed19d2fb2645247b872;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haac32a57df26146106bf6d333261c0d1e6b259f375f04bd3983ae2a0593e8e95808bf699d924c6aa43e5b0282cfe25b037f909bd6ef45a4181fd8515843e84a4aebd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e896913ed09379ac6e473b77f65186d7969fb480cb6f3341aed6b2b8c573b37c03d32115f9404aac29ec79521bfca318194eb69f037f657f6bbe9571b8d030a6a108;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ccfeeeb7d38c2082d8ae70d55dada7b41adff0e7d13a45362c7e86f462e378593067507e5e95eb7863f6c117739c2c2627645778a7288383cc7ebe4713df38181696;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h131266f66fa559772eb422b2ecdb28eec8d591e2e20271e95c9ecaad9068483ef387b8c67831826365100a41e414437ba92ef47f6d9cd7085f65e9b085f1e789f08b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb691c58c5c54bfe3e437f4d0c1f079aec157cfce4398165e15ee88a071f3ccfaed02e751de72d21d456c74b730fd5ed364ce6f2aa552e61e5a6942d29f1dff911fa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8fb075d318f96b9385cb6e69a1722b17fd22f410bdea10cead2cdc71477102c5b1a66c9e826902d1aa226ec71fd6cea1e77a04e2cd1e6960a97ec1e1ea9556248fc1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9341f1157bd783ce7a24d82a4a06cca1ecdf71867d0c907938456eb62738a83b6c37e5dad7578a46922b8532c467ed03601cd99c098fd4e9fe2c2106f42e50439b9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbb73e627b4601c28b3f5113db4ebb5a16d9dd782d958931c92aaa13664dba50ed7cdbaa92e939a52575a9d5616ca30e35094b753ef545c0c514ff5a34d4ff12654d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff12a19e2248f16e16d381d6ff1987a387ed550ef79c038164888cdd60a59a4f698978c9fa6b20931d78d6ec2d69bc55e478e94e7b5c84825a1794e482f6bcceb3f9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc94d536c93706abe9c0de58aedee1ae4be7e9d4b9c1347c6b87e3885e3149cbd63b26d044402b7ffdee61491c7d71434f32dfda4483691458a942e64b16737fc614;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d45639db589627bff2d177b2ca0e87e252fade5eecc7d5d5ae18443f07ea480778d9749dd2c245d3f70ec70ad189054de72b6924ac9e60d08eb573213ecaae03e65a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d2ad9d86216869d32db7930c2d5277039bee96f98ea90eb49390b83281cc83ea93d9d2bdf7a2202da9e753465b3427467c3792af95444f2bacb3859972771878851;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a70d7935fd64612f402ddc04a5c1d23b641d9ae11afb515eeb9ca69276d879d3c140db4f13afacfc1a7903279c37a62cab11dc601b61d6b5bee16410892155c12c9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbdae10f6704c4c35cf768d8295ef897d5aab8ca9cea03d61f65995559f325eba741d43ed4489e65edd3a3d486f4ccd59fb9f20e6a3092d7672ed97dc66345ff239d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h130ae8e624345f1cd961f1b07c8d30dda3b83fa96920d9ae3b912bcabc8eaca5894b09643b4193d44312e8f765ceec1c778b2748cff58dcd87b511256f18e67ce09fb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17754857829aa58ce30c368e1878e5160e5d4a003570ab451e09fecc28ae137c7a6edc748eae5501f5e1a870abf1a637cdc86f05b69f5d331f74ef6c23894d497bb21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67649c7ef223f724e97095e9e271d69f57e6dbb4706150d8ff07de08c855087b82a3efdd11962abce24f679277b98adc00ff161a4111a2dad20e9c9f12ce1b687ed3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1defc023b03408d64939844a229109916ed0958a805a0b528037d12aeb6b4e1af7b809f30995b1b4628a8080e52b4c4dba51a46e51df7fb8392ef6b9f8efe21f869e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h795b206583de976a2cf051c3f180e06ee76919d5ee9fe04b290f64ee95a73f36bb20a7759708559356ea23c5c286938a7840ae7ef82a89a026adfd8055b672ab66cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h78f7160cdca7bf8cab5b2f121394e70ff03251b9386642bdbd7a366fcdbd27dfa600cd41d8532b8e9bbf7cb0db5d5900e266209ea33ca54e86ddf2993dc3e2249dac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96148aa47079bebfa28a3de4cb29c404c7bd583dfa0c6de2288f07002e00e61ffead8cdf8f5d59a42ff1402d938015f5dd4992438c1f9a252a57d712bb61f8d05cb8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9bc9e92b4c6228fe53e6c2f348c5df655babd0538c561d5187f315d1a9b57b6aa73afcd75bc9c096730624d2af8c31f5842a332fd6b2d58507f686293a6ba4e06435;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e8cdc834170bab5048032681d090bfe3b3f805cc0d5507217779b3a1e3b667c2217d8c7309a4e11f4dd9cbc70cb1b767a5fa8ee1d4e693026ea12314130ad6f57f2a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8be8ff26b80da4ffc3cf2f7655aa70bf0aa9b2f039ed638405fed66806a324e16847dba1d7b270f21f1fba9e68d1ed5e59542150df260aad9b67b64036c4617c17b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h307e69ee11c32d7f888f88e3436dc92c6fc42040763e0de0f66b22c13d90e02e4a9cae4e7723419d18b5b321a3c44d6efde179941fc7d9d8176c966db58e3f4f6228;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h142d9a8e909f065c45cbcca837f09e1d2d7737486c0f1d2f8cc028215932584f821577be6e1f7b73a602376d38ee6e69ed56405e3a8e210fe4ff89d2520e7e3182e45;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h154e5dd3720dacd6909bcf951df37d3f6d70b079074e436fd5791e826c88bc74b92b039a5adc64f9221f93774f97b0e9ba6fcdfe19bd9152a0c92a6db828288c5967f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea9f5e832e20696b85fbc27fc5e1fba69d2051edd64d6833d66709ab387c558c40cf4139cd6b38bb6c51f56c6b8460d0b21be755c6c22bde120cc4677beab110f248;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h908e07ef07aac1c4ba6628c7b8e0b5275d7c6dc043539d43a7b2eac965399abaccda2db4be4da1796cb57d4f43c1a75257c734e4b3fa3d96981ac68e5bd2f5503d9f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h809979b7655190356c7e772239ddfda94677390b6c3c3058786c000900fe2c0b967db65f72c35f2e240039f0fdaf953732c93c4eb08b189cf3c8b17c8251c664a836;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3ceef563b3a068dfc6172c7b5e78772c124dec2b405721eb2a98898f0a5016c9c6cbb484a8987aa6f98bb2c417911b93770e0991ed1bdea431f7d55dc7e38005510;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b33be9ec0cbbf74d826a97d09fb8c348f1f15f5ae5d5409c8ab9bb5315588c9b1605164d34da0a938128317a670178e8fa92d8f797dff7fa4891a778a6b16a77d9fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ba0f7baf94fc37c9d9d2bd620233d0318d160341be31124cef449ca3a9d157311020f7bd4b1e2a672421c74e4ce2f394fdab6670def5b00c8bfbee5b07299e1670e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h59598330db7953bcfa993bc2fc747159872b04b6a4a8615602c84d3a35d4773c3fd77be7d1ba12897dcd2e9856a4262bdbb78ad0f5d72f81b9edcec6e6acc9204a5e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b3c8630e2672a4467e939617f7cea6399962d1163fafb961da72c0132105cb422924113c0ea445108e9e0eec721d92ffa15475e8b2f9d6b64e31a4b57d2ab8ca87d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd78b083ab77f9ccdd689631ff4eb4e9d5ea11c041123cf24e153245f6d93750632008377b33beaffb766a0e6ee915970622e5f8622dd58240010b5affa963ed6bd12;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1124ff7a809e9eff2c173dc70ceaa9468e29148e518057e34af1f679021e66a5d5f5abab60b61900ca374f5817a8deb59f4d26cbbe8e481912efb726739b4c531f992;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd361395247d1a8354eec46d22f9f97796b1a95d09d308330a999cdde3d3740ecda0c929ab20dcfed957dd6d99862614da9063df3adfac6f0a0d1f1b1c578e344ec4f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1866d955ef654a5340c234c15893f2e72d404aee97b19ef1caef5edca4e8600a09daf63bcae15f453a804f342ffaf6f2b3b6a10706ef6cbd3938ae7c37ce07235d4d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1630ac93a0a263ca76b076a5ab37aff249581eb1c88c456d05770e5ce23e8438c4c1638023fc6f3062ac6dbf5cdf08251dd8641d79d73f168583489b5192be2d190bd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e800e0034009dd7fc64e831f2aded31d0f7396130ffd63fd23ea31bfa51624212b8524404de6de7d65463ab59a216a5ad0dbc6c37bf8a549ece30c70b12a3b82901;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165c1c9590be7855f349d4e5076a89d5426afa6d1a6f14fa4a2c6e207aa2296896c0612db87b351f8a70d4116c1708b502018238e46987f0221230eef8418d15a5e19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha9536c6e88f9d68892151709f296d42c966bf2dd8669356a2af9aa077ca541bb92a84565a7f835eba76d36e03abcc9093fc88af1a01803b1a4a5ef21f1de0b6c410;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ede4e9055d32e6b21c767745759b5559fde7b8ead5512a87956f43db19494d7895e1f5de3caf5232285b1c0bb8bdd00a441bc1b8e239f9c25326f37025c810bb45cc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he72ee51b24f66f4aa64da8637acf4fbdf4dd15da2d91300bc05a84dc68df1edae0dc9e6f9de34353d0211e23fa082d533a1e4cfd00f4bd248ccd279de977991bdf08;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae841c7147d7dab692e12cefa26c16292159add32890f96ef051f821216d82fa423ab98788cda2524595ad3bace822c99b94a92dad952631463070971d6a2be187fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1038683e33ceffe727a1558e5e5405c26d35ceafcbe1ba2c09e3fe897de41d9630d938b9257b1aee32bf3e8181e2dbf95d9c1a97ab053cf26c81e31c9caf7c835cb94;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a2d3511bfb3204c819347d79d3fd07b232d8ebbc492211747902b7a05ea749f192de169eec82aceb6c520134596997059916a8cfd16b53be404f496f4589f71ec93;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d10c9738677571c8687c8f1cb22d57731aef99ab381db4fa10a5623dc988efcaf9ae5e33a94e6226dd746a82565c2d76ff671afc4ee9593e6133b17160a170daf2d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hef67917bd1fdf1e00e6fdb15263b7aefd489c72caa504381dae088e7ee06f4745231e5c42fac2fe08adaa1d52ec8f50d7dc126d62c4145c1154eca58d334d481ea5c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ae0bcf2b5cc48e7460c29df1a5d1d871db00e527754f21a31695d8e5c021f81a2270a0f590efa317b43cc0ab20de9c01487d234ccf8dc4d74c737edfb52ec7e50fe5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h115604bb93bedcdc7d98fdcbce0d466cdbd115367a3f0d135f533fcc912d50517be9c555746e7c5ca8b4f2787e3d4521694fc035b81b040b7d44332a269b2379e9ad7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h47867c27c54b3c60af420b3ce0efe2186d9a6aeefe6eb69e3be52d5eb102a6861f4a38d5b0f0d751b21ee04d9348351b3944024b6617af4e561fa089fbff6841e4a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d9eb7dc87df56cbabdc53c552ff6bfed7e07e88f40e34c4d2a36dda03f0c99272167862b79a1ceae5d1c0a6a5ee6bb2d5a9244742c95e8505ff268261992b0049b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165449fa44b03bf18c8b57d2e7f73fdcb80d7dba0ed5c79fb53ddad061b8fc61b5e0d2e9861195873033422da1c3f97526fc12ea3c0b9eb6e9aeb29377be4f4fea9d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c2e839984ef2e395f17cf7868448dc844ece494dd863c5c65b913aa071490791e11135ed110acfdc1a5d59c639806b6017a45483c2e145c1531c2ca637db0baeefe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1994de91ed474c4cddf5a776a01bf49d06e9e3a589a45dc419e1b3a56fa1c81439ff9e1712141d4ae7a3a983017d575d084b3239a2f220cb3d233584ba01a77a06d34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf210b4583097cb1696e141ab912099eac21fb376174603b8a26a80f40fd254658df6bf3f738c93cfdf97db19934a0982d14734070dc97ff55bf74efc5185c0d8dad5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a32b9f0cb3fd9f815ac0876114d931e6e66f244259bfc2f6a1fc07597407308e90a28fd91df41d6a64ee519474fcbe85e2bced0c102cb6d3379d9d1123240bef90ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf20258d08ccf90a79caccc13e300276b81f8bccacd043cf9a3da1f45bd3ab3b5e77c9d78d06e187b97fbe466272a53f7444bcd60e333530dfcbc41e120516dc3bab5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h41ba1fbea5ac9a3d8e7dee43402b19b1ce1534ce8700ee8227b22b92c2be1aeeb70b09a61a93a1c4fdad1350b946d74cd8926f86a115de53548092b959e4116d25b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13cc7c7257837eac06b707697628889e1b9cae2b6ff9c8619e502d7a1f3ee87414960ddb242fb233b071b30f86bff19a55378ad6dacd9d6921a80d17f1537e1b4031e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0045eb4dd56d45786b8c86884f6a04a8b028bbe7928634be1812752a08d19aa42cec649300b0f862c458df6cd5803d592eee9ed2fc117144f6d2c8616cd79ec7540;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bfecefa5e5c465638a2413b9c2bb23d9c8c5ea3e30a666f7a2fdae05e50b7f4f8fa3b0923ec63c3a21304f0b4858ed09212cad3bb6c85016d4491b9b159422f532fc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h76f803b944d5d3eb60360916d9da8d47462abdf29e6d2ba07f5520a9cd3615d1cf64ae10f56e6f02d405ab83d9206f6a3d3b6a69b84d29f5e0f7032e7007cbdcaec6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11552301f1cd2f9f4f03662a8800f7157cb82491b76cafee60f710a8aa87317130d9617df62d17773f3251d254d363d9562965e22a044380b7d4aa103ee84496a0efb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h559dccad129836c9728d55f7a5d72922405414ff1e96898d3a1909e4e2cb292b7efa608895927f6bd73964503f212a778e956711f0e0d71d897dd1f36f787490a691;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h167176abf073ec158485955a85399710a0f42f8927a0fe9e1caf0ca6e82d23d65024cb45040f079aebd9435dd4c422ab8be33898403385c538275afa4542b9f73d877;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd0e71bd6a8c279c51f8891c82a124d3448dd10fe2effa614578216c74d9018f57c895ab6d2e888a5483007116f54656cc9453697c0e1a1c9426d3e237f5c288922b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b10654d886b8f59f3a2d14802a61be5738119a1826b0b328167a05b5de341d458f11f40b0b95797ffdf4d7b31dfef642392de0295937332c19040752e9e04e4c696d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1868c7936185a08278c7d53470ea47de9a951f3a0a00edd51649a611f6aa5b7b95b8de5e64423426d9239617610c5cd484ae591cb6b2467be185409b952bbfdb12505;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e6fa24a470d098b2d6458d4e028bbdc996eaf3ea3d765f807e73c70648da1207a623fbfaf476aa8f8a68e98e989d0c400fdd4ef2e01124c05d0235d416b31591be1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1815f3d9c936387ca8b448c9ace72fad0da2ec74af140d7eac05990a467a4b5b043926701e839335ceaa73c33c8f88e98dfe1c8c6f7c548d916e41c5e5a8ad7145f0f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb113098e20a394dd9564e1d60e1c6040a6a931152f8c92a90bc06ac8cccf04a59545de4acc3e8f9cacc6d4871b68c904948a43ab2a43f26684281449452b135bd836;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde52c8f3d6f7aae0be34dc396a6770a8c844e84cc01762419d9a5498091891b693cfbddf58a425099c23dfc58d3a67b061a87693f20a55f70c247523307dd8a6f1fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5a787e28b54ba8df0e5f400f2ebf66f277d9c12fafce3ed88263bc9f3afd2deee73d1e1545cdf2ffc3a5171ae3cc27b8fa6e3bb58a4c62c87c0d96aedb7d1bb4551b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dca4991b273d8b05708936b7caf25729fe3886949ba967bfeef9cf4c30e5a855e60d93b1f89f0b2ecb6a19793b563a2fa0137cb84f7bc55fe876e3f7a7d59135a591;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h188358e801e6bcdaf0bc2c67cab5f04c08b8941cea95b3ab2d2bcffa22b673e65141f9308962cb7ace43e85be355cb81ddc85ccbb9b297ca3a7fdc4671a1ac0c973cc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h137e9f2c7823a9d041046fa8ae9c6311d169fffa698777b968b8c5e39e96bbd207d530f220528d98506988db5978b46bb4a0890d3663024c8eca651269497ec329ab9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f91597b2b273b995a3737b86e3885593400252fb05661fb944dd16e81a1f0bfef72ca8febd96e6b78bda95e760567b5b8e1d10463ea23f800600884ea1661d4fb3e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b80cbfde21acd8087905e440f0839457c7f20596861608ae55becd0d034ab988a224df7138174b4a9958b5bdbe3ab4c797bbac320235043fd1621ea0643e131bdce3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h145e15ed2f94f7cdf35721f19d6e1a0de9660b05e9d0b2e2daf34764594bb4e179244a53760b3480ce7cf2cf6d09a01b2bca6137ec234641e6aaaa4de385917829d86;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha246406d007ffeaf8207f099ce8956cda03cbdcd8c75925cb5dd20bcfbbc08ff218c1facd1aee6aeb428285940c22ef3be58a1c7b01470f693a4ed27815af35c2f09;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h122c427b6971fc836201aa15f182c030a2a98379ad71194b5da54691e177cc8c662aa9c8b08ff0ab158af9942acbce8d3408d6906ca8dd54abe8b9afbe558eeed0923;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13087596f3b062e4f33c9db4825f5757ecf79a631e856c2714d46ded8cd802f391b8727a170ca5535d04d3678c23701795a2c80c45522def7e774ba04b3afe503d852;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b3a08c49e08d4d7022ea1bb170b1422c8322c16535bde966ccf5b6c478c8df615c886605c3c73a1f17e017c1354a480b479bd16e2aeb33186c2251ad4b497e7d34e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b13b52a5b017fa2d2ed97b74aa8574cdb55a1024eb06bba41b46fa4a34cda1751bb0805648845c524926302d355fbf7974278761ff9c481d833d3d0c698a865e4646;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h32069058d1dfd25d8817ea46340c491202816efdacb84f7d8804ad2977f0af598c188a21daba60c99e2bb0b19c8dc288a2c66c7f0d95e498a3b63afc771b9f3acbbd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9efde996c254af255823e4043ce282ed685d5e3c795cded41056dc4bd9be7411bd8c4f84656f6f10696021423ef77b7421de27fcdd14f6c8200170b760413b66e5f6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbb66008c027e3eb381b20e535713823b1e54f5f6c4ffe0536996ed24ba7387e51dd9da7f88c51b2db4c56013d54ab037a88370775874ef2cd886283be1cb106ef13c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h20b8e921beab7f5215d4bcaa1272b049cc32aca76111cd8c5beae33d68e481bf4d43a1992f5a03cbb3c55809b7df86375d31cc53419dca53fcddc8895218abc3d739;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c6b7ec3e6a3ffb3c422fec406b99c03fea63c3556fe57fb031c95e86b57f265f2de84bcf5b84833aee6b1fc6e15360965af715f0079a38e10814a763ffd823d1314;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1533df0faa96af70ddb326aaabd1704ef64d2c00feb82c9c1e0f871b123d23b0a2d76e1dd02f513e061f2dab86a981e8f1d1614598c16e8606c4c267b730ecfb6253b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d237392fec05dbf4224dac55c5c4b6e4077ba4bc44aa6632895f307959739ea81b55f868dcc4a8ca3b6f7e3faf7c0093db7367614f38d09a8fe230d847407fe337b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194d8be012e224cf8f71d1b3c0e4eeeccd6f051348055b43b80eaba9acb37eff8fd3ca64855c156560444fcfa7a109fe66089c71d49aa63da241f26aff4f3d36abeea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38a1cd8b725bfe11966813e8470db2cfc761546bc55a9d950586690009e16e1567b5a8e9801ad4105f687aea20212103370881def1a2589168845d0e686ed4e1e882;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2d6994687a438f0951c61fb33358dabcb3b311a66ee244a2772367065c56dcf12be83a3401ff49d322a371d34f5fcdf2730906d99f2bab43b6ede994000df86b286;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10424b0092fac8a8c2febcc9c181e0199218ced5d08a4d93939585867cf2047245ade23dc7193226ca49a13f90d4fd9100b8972d8b4d5f23e21af201553ab6a023b51;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c56cc3e31030d99d56dcd80a9203da0a0e16cd41f1c0111069be4df9e9f4fcc941130b000fa9615816379986d9b00ec3e9d9af5b4cdb5192abd6b39b1be31547bf65;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h44a39c07571b0745a8d37ff878defed80a6779071598c0afe091afeec9463e0b28fda50907c8f7b9949ad307172df3901a6837fb7a25e44790b9a37f280686ada6f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34efec011b2fc39347d180f020347eb65feee8260c9faf376af8c6bd0db9231683fad1ba39a1aadaeec83c509e2d7c4b305a26bd61ed8fc1414d2706d446814119c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d03dd70fe12c5a08b918d48997b5d31865dfb0d0ba086ff85bc6950cd0eb9d1dbeccd1b3fc3700a74c0129a32cdf89126b23d55dbf9393907971a3fed1bd90595c90;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b614962cc83fb9b66635869266426efe542cca04963ae6816d2d1470d7dfa9aa657f983ff6e134e0085490fda151d3923402f272c71c2dde29c386622db96585449a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74ce4ebc2ae43beb95ccfbceceb7547d74ec98ba55ec417819e4e859c4d7d78c0efd2452ef7a7624cbac2981841b7d390e24bdd04373920d578d3f4986ad64af738d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h56e8479dfccf6cfd48f3bc280979fe8929be4bca80b3aeb527e48579ca26ee94facea2faa2f7d358cbc706009e1d25162aac8bcb980908fd89a917fef623827feac5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf3ef0866ca34ff0ca2155025a307607619fd549039d50d2177e66bccb444e11fa1e1ae2f78228e9ed467a2a71585ddcb8d30da0dd0dff9ae1603fbaff41b47dd826;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h128cb4b459b6b3bbc5ee722c520349b2fac4bcfbff86c3a3c3917999601e6ad2296dc6e1d416f652fd6ada4a4ed38717ea2ef95a44ecd058d806fc936c5570c7f0494;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f7216ab3e496c509c44002fc089ee7ba342d38ca4a842c7e859cde62080d980f337fef68dc790dab374b5323ee4950ed31ceef487f97dd62e6ae902fa035cbf34ec0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1428705daa6f4dae9c743c295da1d59c9163dad5d5834c42069f63d34bb3e3e65990014fbe6061c1d9c187b89c03623eb79dfa5ace2e4c2827ea3af09c29d2605c301;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f8e06a1553b309bc9694876f0164ef260b8add55e0b8bf4f12a47924a77831bc27bbab8c81dde2b41c7a2061fa0dd9dfee7162a2d602b81df49c63b4b78061aadff3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he0b4685cc95f9d5647d125142c3e4a384006b4c1f3ad28d547d93df9aa905b8aa4431b6c4bbdeb68afe3574423541ae89dce3fc761db6878e4cdfbd1de5a6f3e466a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13b2acb00fef8ace19795aa71737815b7fcc3b4647a8980f27b0a8cf7cbbc0e70f2f0c07158b72cc6225afee4a73aa165045deef9b4c95a7dfb8eac96699f811a1fb1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c3ec566bc2bd9a70e8bd95a6a8a7b51aed7debfbaa64ab6fae476dc0e01a90da463b36f77f7bf692807c0f38e39562ea4cf6e03963fe334619a987f3e5721add627;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e08f180dcb3cb745c7e3329b8e559e7ba6e162e877ea4997f6f34498aff9902bd6a90499b41c2f8930ae6848a21a4c30f78ca6554194f7968ba35d2585473a75e8b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d1e19a645f275c69a03b052bd9535a2a800afcdfc799deb142b38ac5f3f7595068a8f39314cd7f9d1372ac36475a9684620f7180a20b3d32a4753cee1b07557c2d52;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1efea31c58fe4bd42fdd9d2b3f1200b3c600344b6cf54b28ec4932e0527d5df846425a8a59990280148b30a7ba4997deb9da7c52743bceb16f90e52d00af161be8278;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha637c27091900990fb76b893b643297f0103346d2f14b57c6805b3cf8283432e69e13caf144e93875722f79f02742ce115324e9020522dd34a8930baca8adb96ad61;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h25e1639f5a0609148a803c4a2be94ce4c765bc378f26187ecd1a1b86c8af0ec241fe67f35e5bdd8c538c4e94c34c86f322f7c99dae10c8965083c0bc7e988e7c1e4b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1126a2b7214ef6885f5d5780d44c636d8c5c03ca00480c9a47eec92421e9196300553cce2b5cf8b1d6805459707f53258ce4aeea3f27ba35b369b82c6c5fc16a587c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13eb85c0ac5f68afcb26e835c98bb93b28990e7d8b2d77a979228469dc56ddfc8f48e90d2453da394d9502b60bbe9e593f0f169b03c67896c7f6b59bf96e73844ae3c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9e8b7a73ca8ed69eca6f572527b230aef1bc17fa967a0697ce3fb654d93114b1f68139cc92ab1b619cb3a56b78ae1cd33da98f51e8a6cb18fc2c2315e2adf6bab2ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2b74b0bc85cc7288bcb86212018b3fda36acd5cc85d4321302cc9a33876aaa2525f9a3da6e2afa3ac224c7e715b99efb39aca2944aa6d266fca53f026913eb82851;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h140c487621c24a17c9e2aeac12ec315a9f2e6cb1d79e448ce375554d658e92c60936ccee7f30e756bbcd2e65887c1bbf7377bd5659c67b67ac0fdabd8560cfb70c774;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e0e1baa5ea438d1133597b5955fba3acdeac13df495f3509561b2436602296c4031f81efb104a23fd1910d363f7b2a15d83df296276ca471b3cfa26bbaa467396f9f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f902eac8874f3c4fa99403627b4bc86922919c7a9c12e8a425f071511bbde38f1c853306816388a484828a5bb121227b5fc2cfa1b41153c25de0ff48c5bd4f63c88;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a6f079986de3eb84d4217d2668758ec4400292a173b0e2fcee08ec5e808eee9a8a7a030e8d4e9179ce7e3ad08e8c6184e4c579d053e12d9b8ef8f9d3935e56c65d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c0b7d2fcdc6707dc94f1062ba78e1476ad53b045a848c891ee087d21461a5d0038d563e7f027f1003e01b78c96dc47d1d8b86bbff5a1e98f62388d95b23f2acf472;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b77211d688ee0a411750893b27612c0b70c9bfa726c1f9552096d498b50f1b7d68c58ff24717dae7d41e34afece9d55be21226deafe5cf5c96fb38ae21c6f568c719;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b63c0fad460018dd296f42a1450e078b03b6018da92c32863cdfaafb7295e784a0fa5665298d63df0d7df7b1285c70d4db61e4e231e9e3635f68167b515e251ed542;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9e7dd5385d11ee332510831ce6e685e37a9ad0d4f290e3bee6b48ca962d593717fd4693cfa095237479fb8dfb24fe9461f31f49eb58035d5055fb565c751bdbb7696;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f10238b6521edff8ed3d9b98ca499725f13288b81fc3dcad26894c891f52a9d3cee9f8757ae09a06546f2e23ca3be22c7ec3c37d4c993443be0f0c07d18226336c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6734a0020d2eb2adc05abdfeb3f1165aea1e124967eea69ddfb3c5e9d3896edccd1b9771510680bc81f2be8af0800354ed7b6003f1ec11668a9abcf31f1b0be5f955;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c1c6dbef9c5528fb1aadf20a335c94ee2a494e19c922d7e5658266ac8676b6da11bb85da11881bbe6f7ab72d41ce5c1154bf02846cdad2ff7333fcfb08798d2e376;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17e645ed299b42f5802170bd59df94ce4c61e97edc5f22e9647aeba1510279d2e148a8d8a198795e9b3bff756526b5650367a6045e242cb455847dcbf304023e2bffc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1be6a5a57d9c02e13dce01b47e4b0e41f6dc6b22aa6a5743f5c9e834a46302e6f425de9d9626ba8c5be345c9de165ea5c257acd77890321094e1c70061968ef651950;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e9eace40da84b9ee2a75020341e4639e8d753d2318707d5501a9edbb655ec07c0f00ca1e8c3410e8a00ac682f5ea1cd4fffc655c55dabb03b37e4afde2fa064361e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h827fa9a108eb280835978d805903e432377c61d4aafcbe5d24c0005b1e47f1dfb68f0635e5aad46da93e5a60247cc6b67a28a59f274d8bba32c1ef95aa870657b3a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1986c07d01237aebb7f6d6a29e6d3a4c6e392ed2127c4d962d650ce9a855d7c12f1dd896048c6e22df2ff5255b573eea4bef7d633227ca12575090b3a7e6898d7d89b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc9f847e3fce3a4edf9dc34ecf25ca0117280c46fa6eae01ff5b37a7cafe01316f57e7fccfbcef5ce329b8e9f12f6382ec449f4e1151c573d596a226d220de7c6140;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e2b3971a1a08178465b4e2fa6cda28cdc7116367b173a706ec41a2b5ce1aad2028c2f4cf024894aecd6b3f7a89b301dd1610481f8a553a4868baa0eb759c69b86fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc14bbf8229484af3b862cdcad2af6afc5bcecc7b9d3d6a40e997c707035d65e30eae9704132f9a1b130804d30da2e088a6b38e06d34ef3195cc936f6f175c477ee9b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bd2eadb4c419211e5aff2a7bd1dd282b173c7929d87a75ed3ca16ee0952248a29061b32b55c722f718d8e55d05f31eb1c00040b8e6486caef8404ddecc206c0517d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d2d30cfb891258c72993252cda730d005cf801cc90276dda83cd985161c1c7fe04cbb32770fc045d732d40b14a3edd190e47cb9bc1de5cef219c15c6bbe255defc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1382a17ee538cb799a29aa0dcb6fa2e7f4c82b54a6af8b16ff2031a2512a9e375546e669f7bd289d84d6bbf726bf2c09008bc5b39672181e6162ec674334b81f1ef7d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e4dd4a4de573e2dd113c6bf4c89410fa92fee6b7988cde9b138ba6b552f90352dc308b8a889f8c5e38cdb70b2ae1616ff980fc43ed088d89277170aa370d1562cd96;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he1a0c379c85c736986fa937d4590d8bbb273c6b57ca43d9ff363583948568fa34f19c05509bfc056efcf609127cd867d93d0eaec4f6174c7648347188b197e5ae7f6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h137cadba707e2b2c3b27e2a92ec7c2b6d6ba5af20e073da7a68da153bfc25c05e39fc3c4cd1c4fb874a7c1a36f9f01a0c2d14e7bb1407c9f3ad036f460e7271a224cc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b9fa8c9b2593f21784d1ebb4924e067cb5be82416baebc841ed59443718ddda058bd6b369e00914e6d4267c885b021fe499d4420e050e151f5a19e18f967289bcdff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a3703bbd69a5ef265b5a7a032f1ca759739b81e5850d99fa97d9751299e7d92c1f016ec3cf205a08027fbeea146f5e9b477dd8ba10591bc79d63a1d271a7a293315;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9bb435b45594a12d9f25f9a17dadf0b8e8733df9497d86bb1261fb1a065419de408511fdcfe03b4700068e9f7a912181dff89eb1639f5c3706d17b03d829373f460b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cb8a8f940baa522b7d1444f85ff6c8914e56c7515ea8dde08468f629ab6a43454d427c8aea589fadf7ff4ea9690e3f9a145768d23422b29d96e71eb2f2e37d28d701;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf934b5bf3949e4cf303c2823e3a92505820f58234982ca7f4d53df1ecba54ec40d4b90274af97b511dcfa65a2c32281ee25fe1b5469952f6b41b018854acfeed3437;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6392d4881057baa1b5642bea337e5fa32d2e41e00e7a9c10ad54f2502c8d9e31a5fbe91ad7075f17cf7ffec0c2fe7ccf76ce713f240d48bc7ba82b8fda9c7ff1787f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d4f7208ebc202ecbddaca94788ba63a1fc5cb87822ae0b1c513791809ed5a832355dddeb72f70015d7289873f3b064115b957efe5142774c3304d817c8429baf3ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e5215394c6635bff42eb5c4f513b3350e5986c146ca12dea1cc9573768fd7efc68ebb9223ac5a8228040d10d92b6506f074e58c4b97221bbd1faa05b15f5d841a5ad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9980f630f6e1a050b5be1a60e94aba2e08a10b3c9b49c9b18bdff28a970d443151448095fba88735f3f2b125477d96c7dda924b6e27b51626fb674eae2fa5237db05;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1946a0fbb6dde6a5eacc8b25e446fab7191fe7f070fd0c84f84101d3a579ff758ad3c404a1d12c58337b5258fbac19ab1a744999cebf806fb128f35af69839e3dec9b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a208c987e57552340264781881e7afd4505bac67bdd264bce6431e34d786abaca50df75d387fe752ad6713c7b2b6262dfbcbb132e496ad045cc6a05a1cca04199cda;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h46795b8bdbc1f8d0e97f17469443bb65d0490c8759e120d477187dc2d678ea3a64c4712a8a328f49ced996d1e6a5a9038f08d0f643971e3c5055430384333a0a43b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a222a768edf44421eec54109505957162235fd1f686a9b38454809de9eefd6106c748a4cd694aa9b7fec2475ebfb1d88ce2af0283683c24a51a7d9b5b48fbfe0c191;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c2a69ab271fdafb78a95ddceb0b7e619ea5ca6ce0be284c1bc2cdeeb9bae5a70e339c2009edbbb9aeccbeb7d7082b6e2385105bf1b25b5bceea39b049b417d216bc4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h123b6e19ce8c0abaa74408046e9329a03cc0168fc500134bf8a60f30212cb156c924709576c73d80ab34e54c9940ee31cb943cc59ec72125bdc6969258c2076c818f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6e2f8594a98f4eff1b7a5666fd86e1365fca1fd7da1b481bc3095390c1072a2dd139ae3d91db8e390a045f460f96b0c13d6f85509c86280d52ea2e242cfb7f0eb83;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha00902502da22354f91915ebacaa99048a2884e2bab0af0b56e5ac4906f776a8ace568d475c9ae83cc3d451091353280c4acdd955159745f30b27a243663bb0d679;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b5e060f9478378dcd7e72a9ea29f24a556409814a7b83db2460ad9a8f772442c8dc0e8635e73c5eca7abbc8821b40780b14234622e1e7f8363a2ad261f69178b822f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h697efe8b174e0158eb29bf177a346cdba47b344c73c8a179fb4605be6368468034693097fc579472605697f7d015a5b28328f4819def15391ec9c6193bd3c879b553;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h70a203f5ed4360fe04ca0af199fbd78f1f11e4abfc64901f7f4237b377ce85275e64b572a904f0068a404a0b92c0fda86a984b0024b460b1a5339862b6856106af14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c834371149baf7367b41bab3a8406c02f399a864f37b1a864fd04c5a3901f675fac780d23750a69e4a6e5cff459aadf5b0929dc82e77ee957ad05424b56127b9b0e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0e7862b45497ed68921166ddb5cf1105c3e2733cd7bebcfadd2a6f2cd08ec18fa94746be868b1197168eecd7f0afa20bbbf51943a957eed538adb22c93daaa618d1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h534e78bac0312862bd03c3f95d37fdf167cbfc9d00914e39e3405b948cff4e8f21cb6fe41b23ea79da42837da3f1f577e75f4fce41cf0efa2a8166ca306611386cd0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18e825f8e3fdbd27bf8b891903a0c5274ad23c493845c05fe4b3609b4e3b7530026732ef3720e38e6d86f5f057f5756dbb34d2fd9216c413074fcec220d1f20dc172a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5b46d8f7c0aca3464b7c3a6063133d4058a9c16697be359de1f454019f9d204fdac9ab6d10b44530388cf1c10a89b0b8a801b315290c713a78f3b3bbb7393ee3696;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13bb702e2c09e4a0956ae06b0a659256669ab0e894fdfb0265ec0b2d04a6abde2d94771fd8da3a2bdef8073e58523d21157ea3098f21f5a2624263a786674f4144ac8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h31d1578495aa7f0e4f0c4e6bd33d80f73109afe8c61df59a932bdcd32925afad4b830d465880aed11e48e7ae00824d115f99c3ae9821551e65f9453356d16cfb4139;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17e74227a25fde6df847fc65190ea999ed04c99f6300a0dff5bd8963e2f3899a0b6d9f8fd2a00a2635d991e7a5999ce828881bf6b8af0546c9a9b55870c0903d0dfc9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e90c57357bfa2bae7ecf6dd47edd998cc409de256ececd74e9aaa5c0b0abeda5a659ba3b1abba22032aebf4219ca073a9d84e73afff8f023cc0c415a04ece3245b5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13a691d7371f90cc1e795fde5f89841aa0fdd7215eba5cda6b53fa52394d49c73aaad8b106b9c3c66d305361e8ce46679ebda78218797d9ec2058c1abcc8a59a172a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7a7eeb458e4d992bf1a3a233e55c289534c25e303cea7a8041294ad27863117f32534bf1a20a14b81946cbfb337b51dc50f1ed2b505589e937978c922be139bf4fb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17ca6bd91bff7596d40ceda5f52e9b77b5169a7835eec79e9a700d5be8ee64d4192feba0decc892f5072672c2d2a0f064d3544c04569f7dd327689666260e11c85dda;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3ff939b99cec0600690893f6521433e58d1e9ce45c5be85ff6231abb13a1031430b55c0897afaa2c6dc0161304751bf953a8555230a550be0a0f24576bbc570458fc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hebfc7d1d79090334f4035c37e7b6cdbde38ebb90c0b4bdb6b048e4ada24b7f5b380bbbb008435bc0fd9f7e9ecd9e0b989b6dfff21bdb9cd2ba5ebcba472065f24aee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fe1a57c3b0505b31eea0cd47209b34f74841db743063e60ad7a89869de4fcd1871584c8cb0c16671fd8f1ea97febca5930f97db1b22a6c9859c55bfe195c68e6ac7c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h179d02e7e5bfcbc61659c2f5d22729468f2d2a19f4978820aa0660d2117a9661b381a02ac4859948def8b553b2043feaf8c19c692646a1a0a749f805d505aac1c9b95;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a45130f3057c7fa3db1cc02dac75562fea081ec34f04f981c90ff84eb1e29ea1bc24a023034b9771b1c0125cf5de1a12c6cd88d67bf70f230c9c53f834c71dd38e6c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9eeea61510cae1b083ed0fee5cbb391e4dcbb04391a2308fb0f2341fb33147dd1dd89dcbb3924c0c284b35b26e8fc7f52de6092140bb86da69d5c399fac30dfb5a77;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7de34f4d09c45b4515bfc9d032131ca7b60f725c2a2d8dfef6805387289ba2c24cfc0c093a8852e618d17b68086fd06a10f33d30dd60ec5710981e4d04342fc5ad4e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10d3e054d3179cafda1d74d7eeee8d01ae3449f91d613502328ddc0b82bf6e2da599140c10957d52d2c20f22a159723477193e3a5a05d7657d8898b7de4c61a50be03;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e34af34a392ac988f79b21c1beb7d3c97ab62544e50a4d553222f1ce33d508729b7a922dbbc990172a3e4e0f57e95edba3da2a75fa844886bfb0fd35e5e615c0c0e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde85c48c6b8141de531a86df8bbea2effae4fe3ca6d4baed06894c73a76abf148a2806ac2dda33d1ba0fc6d4e3ad56faf837e508d423bf1f5b2dc7eb4d944e43ce88;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c2f92777264f364fd6f11eef109d76fe8649ac0e0dc0ddbb0305e3ee2782c491f53a2410c8de973767649fe540fab74b887b21b1cc04b20524f4e43bc6eae893ecc5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb2d4dcb402cd6806ca889d722cce6d79d74964ad07d162d0cbba9562b74e4dddcae5acba74476495cd1e6031d26fecd26696e03d0742f2bba99e49223808847f7dcd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d52b810843eee8e693c1a55853b27c87db5b020c700442f5fe6f9d51df91a35b83c27a79786b2e812b11ec90fc2e04ae6e409f29b8a0e7f5f2ab971f5d7cab96b8c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h110c9ebfd5d2641ec279060caad4d21982fdf028d43265ee8c7f99ccd5eff05aeb9f70f5ff297b0f1ec1a439eee0fabfc8c0f8eec60e7b89b4aeafe96e664920aa16c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e1ffb8d78c6dd2a46824317735fd9a3692c814934d9517b5982af138a332d69d301305a92165e29ddba4accbbb4a01562ff8ec9654a09615d86c5aecaa2b77dd1993;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1568a6d9880b0492bcb0f146a69aee36abf1ddddf78603d65a2610f4c8dc16d0b36da14f92798c0d095c6f2698b98e06ec0b8c79cb5d192f555e950bfee5eeecc45b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb6df9b906825b59f195e2cefe05e2a1a32782f136a348ebca37076992070c5b415c441ceb5d7d735585b806d9c553ff9fb37c37e6ea0fbfa2c0ca1a43f345f8f09;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1447bea1bf7e0e71f99dd3689bfde8644c273a13729d7cb776763feaa3530c37519b5b1c5dd8fa0bb664acedc4d3c1221b1f6fe2624c6be220dca7e07be04c5276a2d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d606873b3f6cc03f2294b474634d1bc6956d772785e590e201f7827d8a0887bd17834126fd1e8392cdf9a16cb8078f6a46296813c49c50c00465428b3d88b96b2658;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9ad984e777ca6a264260b79f4fe5008acaad7518900843be4b2117286e1c5281bb8c6e7e9777652a3e5e67cb889b7d8207931a8b7671fe74f96d7e3560226283f6b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f03d9128a471a1a59fff92ec9fd47dc390ad17a1556e5ccf36feba62595e6d3cf490e107b11fdf3b9df2da6ba94c5a8a67ccd0c89548c7834c84f43c98875b9318d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc565c35ee2ec77bdc2f5be21ad99f6f663fc3efe07c9c7cd297ac787c8250e6496d27d2f81a52e83d05ec4013b74d3967c79e4f34746c320c1811be7f7a1c4327c8a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h714921dcbbebcbc7374882b25a6fccf9de42fd3033685c572515982ecd75fc8fee2a69ceafc79921f7eacd044229122c49418918c5d20b1999a88b39ec60d3038685;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e62f39b934d9132684dc34f57031d3ac3e69a1fcd9115f1f086d0a02f02e329ad1607494442a579f53821ee32e15dcfc05cbe3d314a6047bfad1460b903a62afedb2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a6eacf59090e01e8e44f87b026f13220e973d984d32e72821d8608d7538f7a11b36ad4bc04c6fd75a41e1f0fa36644fcc0ee6f9ecdd415f3cb34b21b48aad00d559;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16b9773ba2632cb99697de54c1a656c2527492e9353c11449cc826e6e05b2ead48aa16d851e1d475d7ccbce654bebc121ea6795f0146cc35319a99f14e49300d04ee3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b1578832ea45e46cd297c7eefcd73419aa5c5ea1ae3c8c63a7d86967d1db1138adc3abdf714e5c7bf1bd314b1ab03070a753480ca9a6bcfea32fcf64719de4c5d99;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h59152dbb952e85922da57e1237988848335b06fc60f48825c39bf3939c43a46c5d524c271500173409cb6fd9e0e768c5ad9660b671ed98e4f9c1ca96b257a3a704be;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd9b6805e5a24812e4a61132f15114741109507f7f26bef2e32c7dc85bf779105ad7ee6ecaabf2dad85536b9372b10705f726122fbbdbc096d882f479a636a37be22;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c21126e1f09d62c7540db27ff48fd14be2ef01ae6e2fdaab364b55ba53463b1021861c6a429cd6c5c9d9f3908f13c5d72762b3737198d8226e37da25c5d3a06a260a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1227f3f8437db57a4570b99862bbbf70e8da664c0c1596fa52aa8499a053ca9c8f9ad520023e3472ee701650dc2e7b41a327b4d5764acae7cf92e338cf046f4221480;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ce129c4e1b2038d54aea2172814b507a8b7bcc048438431a7e0bcfe5b06d31c43f278e957cc30e5a2df05d6eb9a307cf8ca29fdcbac9d3cf910b63f07a5ab7a3aae3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e927d9e2a9f9c25e79d014000c10967602967b70fa5bf998da99e13db996c038df54d73a78cdadb10c2bf014e30b72c9cb11b48c093032f0328657f19204837eac05;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d06b212a267d99df56353beded36c2c7799589f2ae2dcd39546c51d203ce15464b2635b607254b71167ed180cddcb395d339bacad85d4dba88bf92b4969e16eb308;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h102eeba2babb88b09dd291896087ea35a16fea58d0fc8302103571a56b1d11fdd1ed6146186966fc0f4dcb597c8c027694dfabaa3e19f4e77adc145453655acde541c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f4fd6bee5bc47bde0eab837056c182f918a370a2faa75bd43bc2b86b34af3112f6065dcfd413ffef1342e170656cad768693d87fa0a6f45142ac9a4119365e4c168f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180f660fdf126f113bcbbe615aa9292e40c00074251df823a3726d0d9aa9249abad509ce54e0903b93649cf93142030b8785dd6d38a20e9f66a2a2e748c22f68fb0d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ae4252252f88715d948a8aea6271ea9e0ca208d5c0f6796251d9c8422ff2fd9cc95650992b485872d36dfada7185793fbdf50b2f1a6e11a9f115f96e30352d13ff1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6b170834bf23fd52930ebcb6232e7a1f2047040ec6c4180fbec661b9628c0381d776958840af46e150582991048b28956bc8aafdbbfb2840e8af642e6ba9bec338ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1074db6933ac529bc12883e9952240bae8ad1c4c64534b3397d908edac53a65eea296cb197db68a10d17cda4a682aeacbf06d84e263e1d1711289a24b15a21083cbc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1160938ecaf84a4483f094c58f1c54ee659558df20c35d5164ecf0c77104e47a2d23d9be74582b0171e883e83cc533e0e5a0a25da8c3657e648cbac8edb7677d6de39;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18fd8a188495274adbf7e4d9d5b1707dbf5edffdc5289bba8dc11a6c4067e2436c48fe6e1ee7051fd320910615a9512bc916ccd6a95b1d6254aa4962ca985a857d9b9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e6dc35e6d8d5693fcf694cf2572f60482873b20f29b3d0e7a14365222fde82499a6ac123e52292a8683bd48e90a532b901acdd044d78694389e80dc3442e8ad40ec5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h51bbe0c7f813867ceb119a7bde79d92ab43b35933a47716e63834ab4c1326bccdeb1878feab5131a77cdb36c2ca252064098bb3b3cce7ef24ba4cc6e6e52a236c0fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11eedede03692a34cd43ca00f542671d1262295904ba22d290d996f33ecd08ca42c8c834c23d39d07f519ea2a01fcd9f55114d8770bfbf17959a5ad05ad5b8dc3250b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e96b86051c399778b6a8d86b9562c4e1d9687e95b2a1feeac210834c49dc0bfbeb8df5bfd5220d2467f43cf48470f58141f6725ada089be20c7ee8e83fa6cb7e9c7d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d89544f936977d262aecc31cfb63ba2e10f1adf5a225e98a780f66580b67cad5a8655264c4352355c8eb6d51bebe09193bc99f0d1acc8e0d5338f2323523e3aaf197;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1188d3b870862cc9833fbd9e4a5cfbe2d0325625c4cb93b15cee3b10b35e203a920e0d47905ee67c46c9100258ad903b0c8e9f09b404c8e05b6e5266e6340d402192;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h167d76165400903abcb479256943d9b25be67985ff86f42a8a58eedbccfa2db4bb81545d6d034d48f4e53b962adae5bb3fee9623e928459dcbb02d387b2b8ebcfa16f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c792115c1ee1056095528948cb5649a4c54926c4b76b9b2c93b2cb22318be60bf053508415d1ed1a5c1b336c769bbc9e648e122389c7a805b01d111c66e3ff1c704;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e104d617bb1497edd0c3e94748094ec7409367ceb59f6e304d8d0436f51b6e95fc9ce7260ffe719578dce5779dfe8d8388b62d72348041d9203bf99f0baeed96bae7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h181d9a19468b8a78684777c83fefedd2b18c7e6df3c1d0bd2ec30682054f9b01b7409ff7888b7842fb3419e52794687b76fef0a74b3dee6cc0be1ab5eb9786e47fcbb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91a85f643adf14f75693d88665139b97e0c31b87472b35f6901e069101e0d09ebb4efa430e473585134ec0bcce7ed85ad2b6b09763f76d06f2dc2823c45cd0141546;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf76a9e102dc337caeacd379e3dfd0431bd56b00224e5efd9ac5e91c46686d80f606921a8c55ac2e7febe705e0da404e33e618d6b37cbebcdc6e4aabf54ce8b663924;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186bfd085b5bdd117b23123ff0e661da62915f717645daeb985ed7997dc5d291bf7af1575041a3af0e21663387f384a908925c630a0819f27af7b88b8ed8598250a5f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h107c72e7530df21eb4d233de996dbcb87362b1b6e007ca7d9000e106cf246ddacbb33a850f7a53b4007ece4b72f66f7671b21a3e439814d2741cdfa0dd8c28a75e90;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h132c6f446593dfaa1204c849c3c1d43bb3f171bea321815fe4ec07edc2504d6ef8ab1674d8f7ee05702cbe214aa9d2c20fb8cc935abc82676083c7aca88500f943862;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d8c829e833d3c4b6257b25cded383e0653cdbafe9792bb51a1a86b0439d7ce9cb758b66f0224a96e2810b6e4baf2323fb0f70753f0c619004a64a6b71cc754eb297;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0ef3428e33db37f551a313fecae437fe6a889dd160227debec6d28a2b12b92a938138b22f624f082a0be879a080befcdde228a2ac19789f804319a2d306f301f15e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a2835717153d8ab7526a15553084ac87632a1bd944bdb00805c60a4d5f2e7383abf6919e498e6460076a0f040fc0e9fe88b65e4aa669b9e52fe02bfc869a2e2df26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6bfdc218238ae51aa7736d7e8e54662624c0d5d0c11d3a1869848f1fca023536a204c562583b144376ac2144704558faa8cbd61b131f0f598f7b04ed7517b4d29f51;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d8887974b28d28cca96eb1c58660da9f246a03eba82cf82bc991d588908b9e8aebfcdad2c979b0a841e12fcafa59726be069c0647d2a300889f04d9aa8e69fd4572;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f02370b3d48e436cf80f8358c9358a561ac3e5e02c1da1a8e62a65ba6c31a060ddcf63d88f12c9a5959088ad52346214cbef9308a555cd13ae56461e89e273e0f03e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h628e2fc3f5444a8b92584d7fc7cabb9ec54782a04f5f2c743e4fdb47f3bfce1854f423af8d6e1b5ce20d27c1ad672ab5b3752225c5c2bce1547a9cc0e274a2419d92;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ce840990579856bc3e9782d64abf7a86d7358171b01a9ad3b92d1291f982af5025e05f126f9c87494b90db2f7eefaa99d5956a1372409050c9876cf69a8e5c6985;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13901affeeb3359258362d684c3f608db9bafb919ae907f987d097f6839372f8ede571fe85f17fe024119d1af76de276365ae07fddb36b2cadba30400ed2d13739649;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6b7c8b2d7d013b8df6ef2e4669ab7e62a7a23bf94b876ec838035d69bfb6ffadf21d5827cfb5d54f2e39c7503ae9e49e073b30e16d61a3793b4353b497d5edafe9ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb127c740b75c9e1affee94bfd97b644211227f4b32046cbab6f390f38f1d16ebef50eb781304fdbad34fd974f73a5ecb4a34f137ba87ba9ea1f480d273103dc677c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h30d61cb85aabb87cec7c064509d95b76c03e63944110ea427276913440ecb3175e2c76f3db7941da983e9bb0695dadbd49c84218fe16b258159330c1cba7d96494cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc7b2e72422a6c5333ad433b72722403dc0a254929d7359181d69db2895a2460718c3c1f0360d4a9df0193f7fe804fbb274ccf44d7a5f9468e1837b023c9eeedb82d1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8c3d8b36b7434eab564ac2945e05a0c91cb707b191a665487b25a37b02c1a9313d362f9b8df1bce5fb0326c36dede7b5d2e84b92603e198443cc7638c5ddaa36f4bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h84920cebbfd3c1111a20e2c6f548f82f13a1844585b79272fe17dd4090cf7fc4f9eed19c8b043ebaa870fd7edc52d0a2565f7d17493d77207625f1b196aa2ed49b1f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9a756471ca7834c22f2e70e07c19baa890a1551c545a280d62c5d752ca82fecee7e4cf3aea29e5837c7afafe6d201c83aacd58297e748de0cfa9e4d45ab13a18334;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13652d519a30f452b87fd5939c170529288be2d4450d2cd215be4a7181f9c99ebf5b0cc2bd52bf39d04f2d1fc789c77603e2c56641190d771fc7f0b80c39be6881fa3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11770fc264ce1e8552c70b03ded0ce72b2fb729be9dea1dc40546f3648ef08e96b2a9d5d97adf41277719e7e2cac7dbd1caea508d05dd1899d7a967175e2ee4fe6fcc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f7562e026542c06288b0385c5cf23a4945ef0f48f5a7bfccdf6338fb708f3ee40d3e94f8110fc694b37f18302c1cb546e9683c1352896ae8188fc503dda5f2240b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h169f763922639d0a8e9388292bd363d52dd5c2e2f9c14cefa176dcb8f1d9de8901cea274601756f28253736a597607ddbcb253bfd0294900c54113cd07f575ac707c3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11116efa0e308c226f508d7ea9c675d64ce2b5720384b394e02829a13b556842e612cc9b5a719c2b790b4ee0f31a6cf6dcd8e0125b6478e501f778028fed7a3d58ae1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165341d1e556de563e09265276fd251ccd1c1c31be3b04436f61094f1dd60e1dacb19034a8ada73fb5dd934df0db0e2b8b39f1de24ec434061b9481b74ce0e9740716;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h551534f0a0e16977490b64b46a30cf2ac4cf3f9931d750a294a5a9ea4f211541d24b0922415f92773119de0bfb111c4da522a2d7cdf08019b6b5a9614f57c299b584;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f547d8f02bdfec5d688279e4ff52792e38977612dfaba3021b89166949156443b2e949c7f94f720954672620627b2899059a42a8669c834abb1cf4dffdf513e627ba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h179feafaa84c86abff89ba6f5e32f011308d320488b0453bf9b104a8256bbad56f6a66b17da843b03191c45426fb9335944c2be9e6b6d985f637ffccadbb10b31246e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcfe056f0d70402831e84ea67cff0f65fb2d54366c4fae37a21d97c5ac61f598026600cae2dd48ac67c669180338feaa225de4edd697ab16fb5211c5304d519896073;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h21f28a29bb94c29a95415b73e1e37cb6eb1779d40e2ced8136eb3d49de80a5617c28b95c67bd6988a6204cd70ad7e7bba236965a93593c2d65b1b0c574973cdcd81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dc955fb61abd79e80f714192e526dfc27f39e5eb92400d8df4525bb55519a62de5aa6da08ec96b5350e482e08f92815e9a50c2b9743bc3601dfb46bfec3822f9f6b9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1154ac8e234d16dc676bff41fe0f2e906e2501ca351d3b7334c64b6b97d0d6bd2e6d5ddc02cf0e67dc4bc30037025aff028b6254d4bae76f0edc30abe8f0d611f7d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161d2054cc1be6c9a2baa902a991513cd925831896d79fc295a119758e92bd61cf7b86eff4f59591293ffb027c5d264ad7c4caadd43f13d8fdd4a5255c4fbc1de5a62;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h98919447d9a6ed2516d53f63feebebe3dc7b82844131a4e648c4ab75530209e9e3af1e6be819fda95cbb07a59646086664605b8ad532aa16f5634063fdce34a0f4d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1092f9e5e9bd547feebe30aa871ae854f32207b4310038f7400a491236c1f99e6f4c6f2a3b22a76e6a0099c7d65a9c958e2652575190cac428d961363cea24748908f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h88e8a283642333f6dd921f76ba80b181027712014cf61aee83ba14140bbf214070e60efc1110ff86b8e63bc9f79a6775daa8e60bd20257abde10fdff0890b1d4a6f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1712a6114ba8422cd07c5654cb2c6e6f916f732530cde53515d3d634bab38fb0799c8c58dafca1499f5785d769278b9c80bbdc7df1d95bad4ac92fa08a9f47fe2bed7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69470f06c01669fe5696f6bb891b1a34e87de0d287a17e47e3e54cd00c0049246e49f47e9c3936d5a85a869f7a0de623435470e8bc4c0f07f8d555d3688e490d99eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h447cb54b75dde3431f58cb4896132e4da2cd9704bc995260350e63e05bde0fcac8ef8e880b66cf47942a36f2a3f293c3855a5ff5509c333e2236e49d007367063139;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d3e01ca9b4fe208b622463a925e51d66cd077b2689915a605d8c1dfc27a6207401585cd0b8b4fdee7fba1bf511906f24afb5c682a250a48476af51df31bac6c349d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e9ba8b7029cddda9af9739f385685ae9716d0c7bc02d243727e69f860e584b99b25f758e7caaf1b5be1aa83107851d4cefd0826f5f0c420ac1d765d9c16e12146b20;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16971af58e52339952b582c140ab4d9883331f48cb248ff4b6ce1c81b17e8a93cf61aeb781f4020fbe62f66bbed42af57e558da8c92341319b421334217b8d90b157e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f74022f07debac0126352cfefcdea438fcca023b76dc418c32f075406950a616d4dff871a035346dfd4fdefbcb1e99d26ed67c3222194dcd0f4cc903ec2f396b744;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3828e2574fd97152dfdb0e1a40bc272224b682d59fec3faebf2be8ce095cdff6ab9e7f4d9ce20ce352343f6d672cd411c0715b23786a4c52facc0642e81dba0800f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bb90572ed743cab80a8cabf9b6139014b7786ab1627db35ced1b1664165f483ff6d10f27b2f3a37d60a2f251ad5958a28fa4fa23e93077d3eb9a51f635131a106520;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcfaa01fb0986f4f905157010e266149fe1513ce9df5b00773f4e4232496c810a865a2356f302e9b50363dcd64ca98510397bfc968206db5c22e358617a5dc2684ec1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc1ecce9ce7467f533c8fa5ce8f238c4c7223ed1d9cdf19c930631e38598c74ee85425bbe717a89be4393ba3f0d3e27eb5140684f7d9d113e87e846d92c17ee868787;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69d094c2b9beda7a208f1f1c3f0f652ff5caebb6f46425ea204c027c2d33981afe56bc944352c1795532c78e547038deb1689ad8c3e83407ee7f81644af3bdb78aa3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffe414a380c9f3f330c5495256bb77b7bdf12dfbac8147b509f2868bb401376a8e9bacd0d36706a8dec6c193a63df6eb8c359df016d40ace4ed02d217de0bee7bfff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f50689a6a8f0c1dec7b9119ea82d1011d5bb3cf48816122faabcbd417cd62424b38713606efccd2a56f674d64639a5ca07a643d5fde3cb3eccbc867a5495daba3c9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he44b4701fcd78807562693a75bc86d64e4f91884acdb040797cc729078060efffc08ea321bb88ad30d6b80deefe4008490549c3b4869e33c3bccde45b53b7d8b8123;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b3d65d8b4f0f3d9aee3fa17ed119000c297dda621a3ae76e87d62ed5ddd9e16581df968969ba26da27a7ee23fdf097f84c6be2c5a39eb4b0f77a36fe6d901d76066c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc735e4a2fc8f31d1bd30d4b76c72de3c404ba43f84bc74af1eb762388b5d26ec62b7360fac390fa8e2c59ef877d4300986c4e9013bedbb0af92eccfcbfcbc68829f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b0c287b915d28e268251c1e855c409c72b5125d791bec0cce81154f82740c2f2eca6e3a2ad5e3b5291b80086fc62c339a6255ee5fb35c261726f365b5ca918b512ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fef97df4720e62b984b7b220ac933ce6c724a2e53ea59c2c1c85ae429388ec29708c72716464d55464e03b1fe969670ef0db955aaf4491e19fcd1252aa8cecbe46ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c97dfd7212fe98b10e8271601b67186e5e2a6b9c4939791377eedadef3fcaaced41b9597bdfdcf4f3d4f2a19bcea3827408e06a9f5bddeb9cd56a747c2520c20c13;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c30392a2c6961bffb3b0c2f5c41df72043dbf8681e9b5900d9e9bc559dc3cd0ccd03b9cb6d0554d4b987cc36df1aebaa7c02199ce9392cafb26b75dc1f3ac1c29e92;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a49668ed2a511166ea54894caff807f17a59ad2b31ace9750b2e0549ac1f527c2df6a0d40b35014187993a961a5ce086c03e8dd12a1430a3aabc65a0a2150698b2c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14db597971e1dc4290a1232c915c189c1f711a83163d3cd63f59f82235aa851f8a797cfe18fafc66f3f3ebfc9bedc02e29d8c56f1cadbefc799dddccd69023d2625ea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f8ed509b7d22f2353434dc18a73036cc8d793d43a35a2679f282bc96752e2f720b1018813279fd8b2fb8c1bb5346dc208130387b7b3854ace0a9f084f368634e2b46;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h104dada20c0958b09ac1bd805ed49011314daff2c4564aec52dd6efaa8c881fa30dea547fa5ddf0789196c72764bacc88cdfa8c062be7dfdf6a5fa4bb672717b6418b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc9df36fc549aaa6a7d679de7c00385956816b1f303a78c9d7d8db77c80d673e11fa4172d940ab0b5382d7d2cd745a9bd11f6c98e90659b8305c7055848a8e8c9285;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcead3f20d8c98f515bc6eb915035755c3bb3d0f9382dde9e9dd6f0aea4ccce6e947364b9d6b993baee7e45d4aba3f87039208dc071997d5305811cf16aa2429fb1ad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha73d3798e0f7a0eb5f84aab68bc1509370799a326aff6a9ecc6dc9bfcf1766eecbdd9ab0f5580cce903e7e615dfd62c50147a06d05bd9d059f1d4c0505b4487a98d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e4a00e519bfb93dc1da357e7a9aab44d3e9a50982d5c25e20ec1e39dc5f2c367f68e15f25cedf723593c3b12500f09a0997da5ee11f02befd03969ed127ba43a8319;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f48941a1d1be48984082cff13ce1770e2b5f73aba2c13ab8fc6c67b8ee54656cc360a7b1dc6fe7579071261ebbaa3cca3b68ae31e48972ab4a50c26a95c86c6ab06;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfec3f769452a183d388be4eefd6258ebed80c9776b6dc5d10bde976de7ef961e7c4273da520bc85a737d2592e09a686185b46c781e12988cbcbfed7a0a11c4b9346c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa8eec6b169e07eb340099f33e1a5af8645232529c8d2367f16ce97d5be4b7509d8fd4e1604ce56a246389418ec2c5e5d0d0ec865c13aa331e4344c00e777bf98dfb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h199038bc609a228b87e7fb63f7bbabf4fd291db1d2c6a880cdf041b8e317199f867e87618b00b41ccde09dcca80329174cfe39ae0ef64f9a370af5a95dfd3703ab050;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c73c01f92ec2b118e97da179b61937db2fb587e2bf57333aec397ddd9f33f9a9dd78f1e267bf5fe7e8c091f195f826305e63c00712f0781602db8f4f27674d44ef8d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e92ac61d18dc032ac1aacead575484da9c8256d1709b135753036df6e6ac54cefb5322fb3bc1a96ce42d7b62d398122ee7a1b28e58088509c9abc783b844028d362;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd9b660bed0f47731f346adf865fb455319f762bcfeef9509f6fe6ebca11712154d7c139c4d0df2136add6dd629a3fd74b6f4b963bbe7830a613b6fe50e6533088bf2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11db10df303e195d1f2e5f3a78a6483ceed859d4bed0ba5e56ddb36b0c449998950b881f744e2343092eca2e0163b89f2715308281ef3519a95b65e3050a167d80e24;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h104ce43ffa6a1d1d95fefc202d0a4908e896e85f64d5e42cc9a75c5e05d9ab64055d6f893af98e96e978fbf1b1771de69075d727e61775bc2e69cc2cd9ae657dbee11;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f8f722272d5e41aa4200e4b8d1c9523cbccc76972e24a84771c0e4cb6d084a5c48962ef039d12e4b32e542a29926d7539598032a63eb162485bcf0ab79ffc6b366c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h131108b88cf461a6e69386e159d6773735d614d43a84582177353369c2fcd847c8ab33c5f04d615d5b597cc9708b041a1aa7c18b241240e064c61e50bef50bc32c215;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h146a12d6f17abf613fb9c0522da91d3597523e859e84d8fff90de087e9c574fa5f7075de5ddaae36fe722533cbf6f78a7d719fbd7e59801d60dcf5463365e493c46d9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc404bc8562d8a8bed0b96486f8be60c3e07a9936e97fb27442fe785daba3e6afc7b169f001c02125c7535cc0163d60aa90dfd9e642e9feb8a7d1495623f5447b02f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7934345826f62340da8e79a35ebb33b96fc5defffc6dff3720a10fcd2ac18438e77cb2a4b7807199f180878c35413c1bb1cbf5014518ae2d33bf25b21ecad91b5596;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a292e1fc0a0895aa6e856d67df3f35c995c065519c87bbaa6f53fa0c5f4ea854801728400a4be77ce3c4ea49a5c9b5eeb68420138e3df29d23783593ae82cef132ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc34993d84c6054c239d2d1da14eb2628814ad38d3c4342bae292df4193d74a688e2008010c3a9ad830cea10d324d125f5f30a8431de4222bf7577ab894f951c49792;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48b5c8fd3082d953f2e3ebfb367415b04a0bca7307472d14fbd34b06b79e5cca7af013e4fb8ef55f479258e4a79080d7c949d0706416d0faeabca4b04565969b059c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfef7ebc6ab800277cf2717dd02b667cb287ffa955719ef73076881b89cc00108f62540d88998cf9928d7247070f1f4b8fa3cea1a58c6cfc56dd0161bae553087fe40;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5798d9ceadb63f2103a94cec1c13949dafbbf56dc681b134b3b0135abb491e7cf21f12522b3562a285193b7089b5d5c368156fa9566c4c3c97f256c2e79c3dd5efa7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2bb7930c3be8e1fe7b8fb4105bc71f397389649750eea6b8e02aad9d5fa14589beafa562bd8dada3ce3e12ad3a0095aca8ce8cbc9753d8f17c1e1ecd16628e6efbb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d2a205389571fb949c178f65221beb86baabc5b7bb6484333d041689c3ec83971e13a4c0fec1e3db2c897794897758d62d55654a0abb0d57732e1ddb455f390ba9f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e146be1e258e0573f23e7196d3c4bcbc5a8c6eec5e84e3b42d7d92107e570824fc4070809e35a7464a77bfd8cb161e7faab4d4c2971ecb6af6e4fcce5899b85d3969;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15fe2b16e808061b476c823f56b4c48d6a45cac2c22b6603bfe1074bde33a2a0db470c74165837d28eee62c7c4bd8309910991388524d39179d29528a7a2fc82e8ac5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h64aa5ed23aa031a23be0ad7eb1e24a6511bcd7d8f6442d9573b49a4d1d93a68517d36916cc4940eb8d7c9bb23df33dfeadac3033d3b4b8eeb0626b3ce4a97e122000;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h109de92ae07e5b3058a85e56c0600d5f9da81d8e7f99cdd30393a7aac8875e198ccfdd323ad1b5f24d626884d40e24fd8db1d010164eac4eeda821cf0d55a87fe1f10;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h152632191b33a6ef0ead6d330725ead8f78e86d8e829faac9ad3e9a056bc82dcd6993ad323cd323d297dc8eff4d8f6bbcb14c4e7e3b4569edf87909f70749405ba38a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha9c4f6f386c3ef6f347cfd03717e29e11d93bbe5e992850c767a09514bfbbbcc63734a02bc66f872b9f4dad841afab51a972978abbef2fa870de66aaf8d146a0d56f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175c776558a9ca96d893c93bb4b63579e8122be6af2888a3d3f82d1a9c5081ac0e165078ce86bf569ae745f3deb201d6c72fef2f5dc814c16ae19b109881f0698c577;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ca296572c78d173b2612593c9a40e791f237f016c88b4e8f929e3840b0d36a42f4f6417a4b14f6c4abe25106ee0e64484c32f846975aef5f4e74895634b61a1f1663;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc470eb58e1c3591849a7aadd32b43936611bef35decedfacb8a1a02e032e3d89f3b72725b1a067bbcd46d9b37a780394288ab29f06d523c43253f7ad9a498224602;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61a0464805492263ea6a2fdce360c83272afe5e354b952c67d338aa3c56e852bba1d5285a1c6862581e1eb59f0473e212f394aad6cf679045ea32d91c14f8168608c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h176c80308a33dec77569d1d02352431fc2381e5866b19094bc286bc65dcaa16db4df89f10d291340d9461a58cdec69476a6ccf24188644fc9eaecce7e742b8b3b7b93;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hffd35062a1e70c98c3ab86162ea63a1c42f85c455dc03984698206b2c3cb6aba385517b3d4e3856b6acb2fb7e510012872433e0012fa3cb90346cb5c5fc77ee133f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h230b54257f490e504054744d5895e786f2a9b98b546b4178f94f16ba74236b0ec213446767a135c0e09fa10b62646682971b81cfbfa1815f851539828fd70df2ef8d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61626899959f2f2b39148492006dcc67342712ff7b657c0bb6291dbd77537a526ca8fb94bf7fd65ffba744fd14b3e700e48d30778aa07b4acffad12f97deeb5c42f3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7988f75d49110e4c6c258fb96eb7d22763203286e20f3692901cf299c038589c154b2675e254ddc113ef9d1e4ce52ff97776cc0d26abcb356633cb6a7aa1c7ad2151;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14347565166fb9363b32b11145e0f3690d87bf7cfea9bdaf7ae820c3bbcf3d42e2310e578dcb71130066a45704df68cf44a785c3a1acf2f1fc37d542cfa28f4070530;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12d7376613f54beb7293db0dc7a96650b54684a416b12b2ff47267a96caff72053981a84a343f3f5ffc25d09c69cd8d27d4bd92bd5202c8c9a401de392094ec31e53b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bea701b026fb79c2637a18dc4f19874c9a81baee0471e1716ce3e118e816d02c1287e8ffd9d345da4681fd31bb20e7d6549781737fe0f3bb16e91e89aecb8b8a4681;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h945a7c17ae154b9eab2762af3d7a1b4c45f49e9580d3ad11b12152384f9725da3dec8d5f13a5704e2ed4a22a9e3bf0cc0a030f7066c2e99db8834379d72816b12faf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1145d2131f52c3e816ed9e756e556a7bdf5ba64930836c4a4a940ab38dc97cfbf21aad827596cbbe814d347ce91b7eba0d8bc461a293ed40bcb65a7def7bdcee19ae6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2f9bff704324a94ec9e59d9bd9a391220d68670ca82d957d5a609aa05cca40aaf403601c6ff46c6a2342d18e304e8256811e709ec54dd64d2889940e6216e5bc8d76;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af0aab6a423638b1f85409122a2d2ddbd5077210a53ba92e6847f65fee42642456b12736be464b69542f15bc6d9248b3d54a1595bf262b3237edb503cf472b525428;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5982fcb799b17765be5334453c96ed020a3d0b022ce43c6d36600ad26ca8829b8a04dc5b2d138e67247134de56a2652c1c123206a14d08db842eca6f5c7f7ae46b14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdfe72d9f247aeab1af6b5c2e5cc70c42b2cc45ca331af5e91ea46aefc7e560ed8f07733d9e4679010e6c50d86b6f10edf5608fe45dcfd00b70aa4537eee082e7ad0b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h249538c21983bfdbbed1277e4d3be3852838068e765f7c9152e5c25315b355372df38d017444fe120961c971f15aba3a2080264f43e0be87231bd4a28af16e5953dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heda94f65f2b851aa3a9df28873f1f587c2fe19ea804bd36c53cd183826f4a68be06045209b9d395ff5176d98214cfc13ad086d4f5d2b87279d54a4f2689f700d390c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b4baeb076ebfbb17c66fda785c470e7ffa44f9a0dd275b497fa32eb0c775d7db6ac51dc00eca70ef53c9024079a7af6990b1d18aad961af966e521e717c53b3e925;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193c061338b0dbd8cee5d084e16297fa737fdad92211babab31b2bd0165021529cc547c0d8e0922c008b1308e5747d18f5c9e188a12516a13dc7d72abf8a0f011c737;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb50d81818149cd59c837ead5f749c24d383639fc7f9009a91c44e4cb3c2cd0b441226ada82dce0e6d1ebd0fd310fae40375a61488252fdeb71c68241ccce51cdeead;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1fc854c3bb95104a967e111ec31c579b558e519e392e770965a8ac861f944836ac55c7ca3a3c84173bd368cb8ad327ec7826a58a22cf7d50bf6c837dff4d08872cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h41a9a019fc908587865fb5d5eb170ecc0ea967e128a42bace5a22de9cd7faf4e8c2c9772ae877650fd5862c64c39510222369c96e815df1680d53240b303fc99c09a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1565d93cda08b56c7d11eb4aaf24dbdb9ba5a75490387bf0733c32b4fb1b110b7bcc0e36726afbfda3977d93233474e70acfd9e75df36633da4c0c43a8e1ce6a2161e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86fdd8c746723ba818472c3ddb62a7d1fb2827943d83e54d7f0c88d2ff9e0f265751bec537e888f92d4bedfc155a909073f61cf7bb1dd64a14680e67d2efc1f66c6e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h212baad59a409e5197dcfc25557fb7094e597c0b570b2021e151f431a167ae09e6e985d769bce2d15ef5ade1b380ee1a45bc12fc1eb3dbea8badf5b2ed2c8152a6c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18bbbf55793e13035b7d125e9a5b2e313f88cacf4e580480e08bc333920df6a76b4c2c989956599df7e84d951640625f40d6be0cf72e157c40816554f97f597a37a35;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf06375f27653d83d5497dcd41b9c4b9857c0ff67e551731d3f9351997c3e2db9e64bbc0d18c75b5d9613b19488a6937f72b82e8a2aefd1fb46b8644b4c7a5dfba46c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h189c2790203a63bfab2d17edfcaf5e09a955422914d49866e1de4e006e016e9de8f804127ba2c3a51baabf8eb7b77388234c128e20c535fe2d71a86c19b41e587604b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6609c75ceabb9616f6052a5e2720cf17107f7ea259ad2cb32dbe7d286a5b3cf1bc5c23b73c520cb924a08fecb7676626a69425b3b11b592c95c10d8a3466b57fae8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5fdff8ad5ac7a88346d0447ebedbd3b8e5929540f54bc0ef6345d16e090527edeaba51c45fcc5ee80b993c3e968268708e73e5998dfb586248e9f75546bdabf32925;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16368b34950e4e3f672e32f71f657caafd7edd357a76aa1d3bc510f9f1be2f07497564789951aa11d5e22622f5955488ed9f5f431eb73fa77ee663bc4c7bfe16a60c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb51d4f4ade9674f8d9a0cb94da9c18a1a6587e14b46244b7e87f60e178bfb82385668523b27460fd3b46a9ba8cbae61fcd17fbaaf03762e19506a3973efa62f74292;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h43ccf315914c8d2ca0bab4dcebfafb93f28df88359694644ccf8c8921673ac0135c810bd5cbb8daa4842d0fdf24db7d2cf1d8086d17daae3cd5ecb85931a7b2f46a6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79de51705bf94d7f92840f62e1cc4699a902aa10f3d08b456d9aadacc3a954f33348f40eb9a5e2e693c62845b991434e84ff2528a4c8d6f9b6040c4f10cb9e1592f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcbd64e3d47bf6b726833af2d2cda6db79f034a025bc3d14eccf7555607a798caecdfac7ed94de5e7b6bb222fa420bc093e888ceb3a1f88c320cf866ff8a75348a0df;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce924a16d1bf4e088f6f79898339424e113654c5b489f50f274c22ed4f955d21de6ffaa44a0d2494ad5be99ba3b4428017c351585fac6c5904ecf915b693068df2c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7aec1982929d3451fc82813d1e26c73ed61312a6c6ec09c7a7b301953926568fb2af11f2c3ac43a1dc218baa071f9c3d25ca6c4400b286fec3545d8320f0e77df2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a5f97f321a674c4d5d79a8f4c0d2d5d96bfe1fb1d5655702ae0bd21a7f859d231cf02b420d0130a74d808cc474a723189462f4e073d65f90ba8567a7c02008ffb543;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c1a22d205b1b93d376f3feb2defc1578c51f40244716a78b91250f4818110f3ac4545d9e97c03852def90bd8bcb50c74085c94959e7e34a3fb74b00ea4f1108c8a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbaccdf8e03bd4a9da3247ddfb695de5bde6428d6c28646ddd3dd22ed7e747f5d22ecc4a0f64134ef0bb9aa60b2cd5ccc983692534445b621427e00ea704c110b3a15;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h51ad40ca9a8c9271302b1d3a2c046f46a18a81fd5854ef9f5232044fb65868e614899b257b5c1024a3e5e251e0f40dc8dd49bd934d6f8d0ce5b1a9802179fe8f4a95;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fb082ce3958e1dae5743a69239e18a524f9260acb50d18debdfe8a97bf30ebe7985fd41d9c90049dc34b054b50f361facd03b059870cc348974251ca68b3496d74;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d98a4c2978313040ce976c989512c73d53d0f872b39ed71d5b7d62947e4d9011eb0b4087fbe4021fb44134b4f0a028309141a35cebe42e4bbb77341d7e1042a0208d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf972c51fa1155ff5187411f747c2badc28edae11a9cf3a8dd55aa58f77cb64209bdb55b26b9d2c0edfefb17751058aadd9189dd1779f1456f572a37778ab3657833b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1050812546f97e463a41f7b129ff5c5638d9f1d5d367ea338d104789a8b78fc675e80e32e73c69cf5909c617f6ca469b30f4495eddfd7cd011b424786908dee6700b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1313b6cb041a56bb4219eeb5d8ad770f5a5aa2c61d05b818929e6f465de00ec13485fdc8acd50843a973c0fbedea3dfa78a14490c9b4526035d754e4aa15a37c62a1c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h123c140297a6cc2873ee310314a5d83e1b4f269a36e384d62b795fcd792941aaff72a4786c3b53ef7caca5b34e3b0749684d7b70c78ff005c73942efb9abef55e19ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c90d29a8569b79e42b6dfac59da3c24ed655f52e86c60fcf58373a442d6cdd46d9df03f635cb0ebeb3b73df3251134a025eea8f7f1326474313a591d18fbe4d3dc47;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbc3c1cbd9659df52fa58c4f92641d2a161078222fbeea9a926cef802a31799dca6b4886c71b9c134c811c64b9c9918d75fde763fa76107a8f2eeb8d1f08006fc7c41;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1efd6fb88813f75a55e9fa06cf7ade6631a4760acd8fa0596ca26bf3302fe2788820094a48492bd56571dddafd730b37f68fff8b0b2a533d454621ef80ef7a2707463;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d3e83a270736603306c3861b2cc865ca876e76f84f89ff03ec8d03f8908bfd2845cdecb1fe08cf6631ae2eacc807d6f5a0055f7a000ae974bf5daf387c660682633e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h158d5e290a0709c15366be2e75cf9264095671fbb4814ceeca1e433fab1ac15786146764dd464ab94ef76201dbc259e582b18e0593c98521ed387b98f82efaec4cdde;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da69a88caf9c62adaf445084f18176fc7093eeca1ce6aca0662ed7987e842cf66ae6ce6d62ea96c5094ca4de6dc8a02d197ecefd9ba22fbc92756b92a82102975afa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h94dc6d474c8661563d79e75d02d6a9fd14c8332519748dea0872aee97da6321044df754f5b8f659ca878bcc557c2cadea8ba84482650f5684c022a926b31d95d56ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f2afae7894e7277c01492d2feb8a2f0b4b8ff01e05e5972c96d0fb52939b930ed58766dfb20142c4ab7bc08624e5cb6cb03e317b726c5b725700356f362d968a1675;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d4bc43113a3f813429564ebabb08efbb5657a074779adcc6b1832920b68f6dc5da0e218f3cafdf494ce371792bcb1264150ed60437c2702ae948b929019732a26e96;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff2969633aed8a5e0c3430a44d30c7cfcd672bd14057d165b32132926520a07f11e1de758d6b1adb3cc7c57f1a371a045c21c8e01ba432617ffcad7f43d07bb568f3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa7504c20fe2eb1b49cc498407895a973487e79e99388d8587ac98394e1514ac2e59ef4229342ad14cbdf3a9cccdf6dd42176bef7adbfdc713292c277fc321eb6be1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bd58f8a1312ed89785d8157ef3904108ac534212ee1c81dabe0bddca09a96e63f9e101d494af38f899989c946979529f385ac1faee19058c4148915678f7cadc2f3c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haeced96f7c71043f265270ac8809ac3bfda36e05945d3d84fb8d25bb6c1aa2e878dff10d354a5f6feedd97c7b3f237999a7416fd8dfbb1c83ed5f4617e80d539f3d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d75a235d04bfe55b296864088b16eb0783708ed5fcaeec14829ffd084777b2ea815e8220a67485d87ea32cfe45eaf05f62ea790a9f67b5f0952e8177ce1c59f1d39;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h135bd7c4a73824a25594e38fa0e80ac5234767b700907a3149d8b7a84341654c1c9c10196f05389493c0dd15e21fd663664b7b996ac9e27a40906a51c0f8616dd8a56;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1de04c7f2070acf1bf3d0d954da073992969a7707f9f2401d3118bbd62a8dcc5abe929201a21e50df2dfd5b2d7fd923ac4cab9f3b8e3958f0028c10370ee84dc0dfec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h214c70ed1008d0ae1bacbae2f2d8ff4fbd73f4444a78bf1a426ff65bb522427e4d217c0cf0a278d3346a9642c752a5cb87ea03064d4e8b1a360df2e31d0b8808d7f9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf12787f98944cf010d900d64d2e779f31a33f9dfe3151ab4be43a32b53c5148ca21e57da642848579c618662ead3df8e3abde20a0a41efcaef519cbb8e52929c0b13;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hff07dc839f306848d98ac4ae4e5c35927f2e0cacb11e9cfd7ffb52bfd8b409ed4cbc99bc23f32f74fb1ae85f8869e315f4d7a0263ed390688d7cf01e31952c2347ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h35f93afa305228d6f10db6fe88610c6c2c76307463c5e9efaceeea986a91659d8d158e071bad1472d7ad64e14d2c3daa6703c6caa50c383aa5252595e6811817401d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha91f0c17c060a60a6cd6025baf7429a39e0eb88fc15cfaa5c9fd0f0f25e9d20015d2874f70381ae9823abd5818e2b33dc7dfbf0dc90534de00fb5fbb813ca96fdd1d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h72b0e1266d444d7b24a532c4a9f0c62595469f5a7392074c7ae4d6743b17c22220e98fd63eace1e3aa3353fa85e3f5195e6430aedf8c6af38a6d0f9dac84f938933a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b11a4da3e0f6343df0d42ea4b9f6afbb9c0d6d508c7de33a10d532a917b6937fec5202289b00db67634a0ffe37f6c0c0ec7550d6adf8146329ba5245be1618931683;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14aa0e960f858527f35cab0e5e402f7a3c6167ce1590d21918f1c84011cdc2cdd5da3a16e4ebe00f1501e07b82fd73e255a7794b10e75b8e5ecaaeb97a1103f1ac715;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b0977e08d7cbd76f4bfbfb07a8ff2f73c0ed11bb7c69b5f7adb2f85a0756ba92e25e2c10c8c393641d8116478b27adc3750edcff28de1d7d3008a7271f342880480;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d03fbf8131aca7af45e1c1969e14922bc49eae71a11afd804bfa5faff2d237af4104e8c3ed647b6f21a97ee557e1ce990972f03f911eec4b032cf8cce4d3a367780c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6e84d35291f2b9e49e5e5ac2e05d4b2b53939783d54ae538b89ea8f5e6486a888626006f47244b369426aad4371f67a2a08384df892ea5f3af157c419d418b34c1d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d548f3a79529e64148cafc2e77fe2747c5d4502260921da78ba561f3788349bef29d7ac70fe4f8c32fbc3ecc56a7e8c5c134f7f1e4bafa4f0f3d65b0eeeee1b365a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8941df89d6a0ab9b2e01b20b990f3a30e5ac96aa70e2f4e9054995ecada4ab386c9e589cac9834bd66b967b75abbd2ea2d24e0acf8d7c265ada265e33128640092fb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h20fedab0abc2109287b1ef1875812e4556e11fcec7ab608b4026a4dadc12303f18c7a24ac79a445a203511c1bae7d097ddf063fe2136304b4cce6d10f015037e04a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120bbc9abccf9eb46fe32cacd2f25c5d01469ffddcfd016547fbe21221cccb81f2468da6c882a5f82216f9f248064d25b4bbb98e54302dc7e8e1f2bdb05428372457e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1814242e05700b588dff9a52fd98a3da614f802b80760bfea93fb027b56c394ec60d6bf00020f3049433ebf276cd28fa546de3a7c2467827825d97b159bd602c464d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17ace38b1823ca17c946387593cd1ef5b48b2fa0c87ce6ebfd71800a26443fdc2e7a2714c0dadd304c2f519f608747f2416b5fef5db20043a168c0f9bee54c7d29e25;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h39cd79c2e82db02d75352356cb0d467793cf72decfee4163dfa6b3d99997ff4028103b8d1d41b2bf03054e49d7c03195ec2ad9886eb757ac07a29769194b9726309e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h55599b61a49e43aa29049721733c4e05f9fa87d61654779a8c1a02967a3c4fa2e6a04c0103ed5804745f0388eb25a9e4a9ed53c19b3ac4868e82bbce9ef6f64404f9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e8ccb2f328b6aa7c7ade0bc15d40a486016966bcca030daa7ff02a7b21f15cd429a43c8756f0ac05572207512b16a19ead47861c5ad525e30d1e6fe96925a081e1a6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc5e237f678987e42394fe7918c94b479377d967813449e677ee59df149653c59cf5462101b9293638fb1fec0dc09494d202fad3f24a0098568bb761fc357553d4dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haca5f1c031ccef070f6e37eaba6ee3edf386b9c15b6f2a7fddd399cae9c97205f2e70124cc0f43b99c6879da44ebe5698fe213ff02d1d0409f2503a4977341a15ca5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86aa00a7af65af624e2678623ab613fde4a25e0b8a6a54348e0af9495911e9e84897657de6749efc906a65fbf31e8819ef07b213623f863bdede65e7bfbf08d8804a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2a3f46f05abe670590db3b1ab9ae46b7ac93bea0c2c7d94aa2c028031bd3547378313ad98b81723b8ae89923813841f2aca164b8b8d51d75ff5c5a1548a4d8dcb43a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2ed27d63da6bfdf199b759f8baed203773bf9aa40e61b09085c591d869facff95c81f8e2ad0cc5c27c1612dc7e747880e49731b8e89173d8c7d411a6d0fb1554512;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4cf39a084c055257edf691da25f9bff5d64144a3fbd0d4c210099b9994b9260ab06f6f4b95d251ce81a2ad80a8e9e8adabbad533c132a1dad43efc1c11d865cc884;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f1f3cf480418fe83d7ce1a36ecd979e677a5c57012b3c1edbe521fced1ba9a24d7917eb9e55383131e60e67bec445ed239d6010cfa127d963a1908227326989b5d53;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hee38b7ce37a5a3345504bff1b6ed910ed368b7344e75ef57b5a72df9e03e0a8a503badf35450b06b6500cfdc6d136f6bac2669703e9e6e6bb0e3fe5419d31ee5d1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e7583373a2259151047e7a4ed558fb9e09f2d9c92350a4bae85c73dbf76dad566b6f11ce09f83a5c948a8bb2349ea5a9c59463edee7cfcabe9b0adaeb9c45807a794;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4f347b202b6e31354465739862a55227778766858b5dd72c32014be4f86d2bef91367e602ac10974755a5924d130d84513d5ddc6a99062a30830d4267c5d8c2f6fa8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ea7e34744cedf732045610ba3e8796d8c5b34f3f783fdbf961b68690513183add00acfbb654ee46c0e2d735d975229a3593a09e7bc58ea4b0eef647eca97268369a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h169bb37a2948d8e73ab1ee54a2c4aee0996cd584548dc6a0ec46605b99b44127a1c8dcf9345211e9d1d67fd05a49ca0849be9c4e2c9ab6f50888f2b1fd87e0b11d6d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he0d606a856940dcef5e5f81a8e1554b4421b559d6392a08db4f1473e43e72790b916134f982ac5e5158b81a044dda1dbd8942c1e1ec50f098b81a54ac7d449d87280;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcdcb33dbed7fcdc98f7daaa35440de3dde92f716d54d6949636301b95ab538e72efda238ce94c153f9d580b8b09d3c5874e21ba334b4831ab26e470b98a4408113a0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c7035ee34769026239857dc01966ad69a93d56c2f8ea20d03a55e7da18263450aa8bc50db1bf95cea2fbd0342d6633a2783fb1ef21b0b91d1028c3bf11e8f774732;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a1f3317b19bc73986a470661b7dff5757efe157a24ab28f2dd28598d71c5697cbe7557df27a43244ef1b20efd2d05f1ad2cb8c5fd4eb6617fb653b9eefe688e88c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120c4c8056f318d4335f5c8ee66e8c2a34e97cdb1f93c6d3409cf4ac242c4a7cbafd9c20568e18ad1b1733b950b8f5a74fb0db29178f22f091e07bd72ac509bee5322;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a580345d8db9fde44e74170aa75afd15b8351dda82e59ff18d506bd1b63b3eb0715955a7d2224a56eed324f7991d072dd016cd7479d5e42fe014f6b7a15bec6d196;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c78c1b877f866b088e1587ecfc8acd2e497f52fe8d9063b2d800e101d1bfe282be3c2988c484716e5fd37f30ac62e5aa79f26f65d403ec3121773a44a10e48e49ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdabbd5a15928e17faa3490bd148a2bf2cd87a6da7fa1b37b0b495676ddaef3abcd07ed49853158c747d9968cda6aba82ff06ab0306986eff5be79321cb58fbdd95c6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h159567dbee64d1cd20e3a9e36ae70742fcdc8852a6e4dd9ebdc7e075765bb5d93710136ce4fd62697c8f4e5e169b5fbb1a16f30aa7e212857932676adaedc5e5d0cd6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f69631ab6127bb8d14377e6eb7c74212c276ad87e590e561b9e0494bc0141d43766f0e3813b2cd77cdb89f57843e2b992089d8650edba3b8bb7ca5cfaf33f59d318;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4dffe37fd289fe9291d45059a5f46eaae6a7aac9d7fb7629816edf0a0e9847fc5b2d13f883de6aae41d3fc8e9b02874e2493f17461245d611b7dff23f768d9b8219a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf5b4faeeac5918a58bd4f2032b98ab6e18ace3d3d556924fee76c6eb28fa81280c33fde0d5796874928634bc78e392fd8f4e2b2d769bd1d031aae5c86e1ff9b41c1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1615c759d27e776296eaa160c6bd9c303ecbf6e68f63293671e1b094bbff27ae4a54fd93875b79fd7a0b7e3d8c2bd64dcd5327a2f0d32bcc6c4df8f80acaab8fab928;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf10361668eccfd0bd673f23dfe16e8526387391291e9eb62700c056c131a3a33813b5faf58fb2968475a605cd07f9e8bdb11e8ef5fd1c7f419627c4fb85d1019ef81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb1f4bdb844d25a15283ddb2041b69efa6776c9ccbc9a439fed147f495898c6aa5a7f9eaab8aca386ca1cb3eed5ec24adea274b9142dabbe72a677bebb830a0cc760f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3d8a90186f40ec2ff270fe88d728174e3f72420208c058c6991598479e64b9f08bc698d8b75608535c93a815d39c87eaf165463a0aec44061a98cd216abd4226e806;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b022c3d0c12ebe82fbd8768b7fdcc6328586d2a5aa3da7bafe2c062ae4c6eb37252a38675a477ac78e5088dd691159fde3c4af129751cdf53dae187f70ba1eb9e439;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12607cd897a9159e953312081a754c17e19fbd47de53bfa4f8aa756ac31c380519ca10a9c660dc36c35122306b6dab5b79363dc582d89da47177c0c13ec87611f44a2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9c887b8cc5e5046268e137ecf9d0e4cb61f8b6b52d0e7342322f4491395c1f115ade823b6da5140088e82d206123d2bbbaea5ac74628e1f54913dbf571faf9189cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f25619e2827a9612e157d511d8c025658c4ba1a2c7b07b10c6fa570904baa4a2cfeeffc315ccbb0a80075c013ebd6cfdddf2d207ffd1f4283efe5094cef0f12f9ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18c1d5934e5ba6cd02d85592ce8e31e7098acee1741b33df072286e571724bb5fb25571fd8ca657882c9dcd7c0eef29ff8bfc522b6751a02b211a5c379620bb99aae4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d824db41a19170d5ab532bb1f79b3ab8568ad703b3cb9ed23ddbba12ed03c4bc20ec35e26829d1d3994028aa43b51e978340be911903ba64c429f18e5c47206c19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118f8927454a5293ac9fa74425f2c243c5610f834bea34d38b5bb5243d3cffb941fbfeb9ab4fe4f56c44e83e1cbd5c970120e2bd21a5be34d698cbd3ad0a46f48f974;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h168998bd65522f1959c3f6d6c07cd143cefdf1fcf1271e48772c8910ad51fd10b92602eb940ecbac949c005eaec3839801e1b8eecead613c8deb75a838dcb02604202;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa3115b3f51ea9c9c1a28be02737a1f2be7d5a49c41868d4df9b259a7b1c8cbb8435103ecbf92c2545495fc235bef1f1eab33b64047dd8097d6ef08b151fd4f96dd6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cb5f0bf2ab9c2aea98c3f0362e3f0880d25c666b81c8949e186d5de0d13cf566da70dfc70c7c3810e470194bac55cbf0fb307d9fd9f1a2ef5d2abb421d891c90c7ae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha1c61553b24d1f052706a34a69358aa773eb91a13feb68c6069c51b0f44e1a092d39456b94f03aeb8526a659b1b5b0281e484354141a41dabf37f80b3d0d5e2916d1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f0f44f239f28f19f2ad2ea8530b8478cbf8851a84c354ac1e4b2cc66342f09c631bef825d6b1015ec10ebe91d5d57f43a51ae88c3d57101a4a50398322f00ba9cfd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfab409234034905ff6151944488a06fccecb429aa0d41753407dff45dd17b46d815f7c2480bdb380076668a1d8101470f64a8bb10341641712beb0b15f7c312f01a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a8bec610d303620755501ea40c44cba95fc5eec9c74c1ae2fc63b87d7ace435e9cd172b8418242e6a7cc7b78a87021b80eec9e109ebf6d42704a21d35108cb90ac81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb92c2f083fb1dc31f7a7db22f41a3d4a176fb23106a5d49f8244be674417b989001615083b11cac9a4c6eb87b59c7e0810fd6035dbceccdeda93579482895753463e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f4ceb1cb96e1de9ad6c901c2a11f973a2593ad00eabfea00525c3766d816de0f88b00a659f0e300678b18ed9cf2fcf19a114888be8b49c070a51064c2911f5318c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6a6da2ddbff991d84dba43d10ee7ab4589a335f75c630b59ed3d3e38d8bb0139ce4680684dc08dd735625f6b23db365ec6109ea1f6d6571ad8174d3667bdae319c4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h147492f9eb9da657f1212819788b0ce8c660496e404ff488cd99fe9c40ef7643f9dda0f231c439f45ef66847874bcad01b0b1ff2b599d54db73082776f48a2a0e6ea1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b52572a478a86f02867272a31b109a5ca0a79d8fe50262c14caf20d8eb9c0458f3dcaa9f13e8d8ce9b390bd302338f2d16522dd6faf5acec72482c8f4f3d36872ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb09244cfd353d99920daa10dc6cbc9b8694189ac856a7a1e2ee55977766975111d2493a4fea758222d81abdd88b03ce6dbe105ce0a654275574bc72d5096dd756680;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118982daabb003145d8b81efa31b8fab59270b54907e6fc11a8ce2052be65d7999ef57329ef63b46409ce9cb150baff66ca54e9766c75a761f8eb5685ff756c71df93;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c46997a2182ff774a2646ce33a70c19196725b356ba632238c126d46df9d933e2688dbe6d5cd4002f0da17b2ed42339982f4cb155382227c9e04ee7822d031b74af;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4b9029405767e51446b7b989b91586d8a4f3774282288c762adc81c2a13494644f366146a2bb0e12e6f61f645b45e555a21501003ff4f60e12d56ddab6fdee06916a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h178ac7bee479cb444ad676dc4ac372348eef367a9b840cf45babcde30d95488bbd26e6391cab668696e2bf4c60af8e5b49344a13ec81821f06b0f7aada398262c9616;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8725d57133fa9a4441173aabee68e35e2aa4353a9ea8586d38db7b7c8f8cfc1047aae299b12fb35189023b6d4f137d491cece37197f52a737d54d21d69047b44219c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10bfee84a857b7cefcc27b40647501756dc83b0eb4c0ecd4fbd27cefd7b8bc8916bab68e632585fdab2f26061a15b92b8ba93b1bddd2ed588ab5579fd8efe36121e03;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1faa784496ec8940fdc78bd24dcf80ef8c1e9651cfa3d9ceb65021c5e3e4c9c4a6356369561299e47af43b9f65b5b40aaf3f7e80ff3c20d047f82344a30e7db90df56;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h158878085e78a1d72117913e3aecf91c3c2c6d97a3061032a87aa2fcb86c129d41fb2ce4bdf7ee6a5e304944856dc06e4c88e5a8025a1743391806b685b8eb93beb26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c5b07dd021bc5cabe8abae5638d3ca79070882eda5b50998efb1f7a3431430dcda88783c3327781c11223c2407308609ea82329da5a52d52d75c851f4f3161be723;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h996ad04f9262e930b108e994457a4e56c6dddc745d5138f1088eeb6dd5ec9d8e7cd4c8b7e5f4cda7f65caadc68df63c91285d7473542e20661f9c00b4f78ad9e4142;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66ea2fd1a7e152f1db46ea50a830b2bb4c292c9af64db4dd787053025f37d1f32ac47738a04c4cee18a2cc995a28e04044bbb8597d625b112b788616e021abf4f6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb6aeb4a3c11f37ebdbccd84fee3952f494af0ea4c70647ad9aea9c99b6552729666dd4a2ebe5881a84179b97e6f7bc15c918f9e25d6d61e5877782d04965fa1cf848;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h898680a030eb1e17ce86e957118cac398b02acef5bab5a07b5144e077704012fe78589273fedda73aa3293228ea8f01287f62551635c1c437c7450e04a7302d4213;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h146325ce0e632b12e8dac3de1dc69fe8cd0c8c72997f337d23f25ec017c50515b1ca2c923147a41a337cdff34b385281acece11996d2357b9a3b153383d45d2817327;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h29ddba707db73fdbe7336a38ff68ff29ebd7ff6289bdeeb15887a86912646493bdbcebe895c0b280b52fab0a695e2b1706444263f1cf18ab330ad04aa9b59242eb5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f43f36be286a4662d937479a93646884de541191d714b9d7f6bb83363abd62b55f9a7882ef1a966431f9af911c0959e9d518f1bb6ebc03e10f4066049a2a804d6ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h128fa2bbf43d4fa6cdae915460021b81b73419f570f1fd5405fffe9aa43df8cc703783c06eb071da20e70e023f0a3f5ee54214720ed8347e24968bfe3e7e29f23bf9d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf99be9928b3feba6215516e0040a60abcdb8c6cc5b3c88c08d7a24a569fce7c6328e693eeb74ab8b50f130bf2d319b61868f19f518ee8a87ff209af7851026399342;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fe4a347c4ef36748d6251e38000eff21c066b3dd28ff948e414b64a28806df138954d428baf4cddce29ea5e725007c5bc327917791a46f91d0ccbdfe418c6797592;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc98e61d29e2eed231f657b8b2640ceb7d496450eb36c4a8cec5e5fed1787218a9daa9079138efe312cea73f178cb473b0d2ccd5869fe61651ce1164538dc30965e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ebd901928d51c9e1a5a31fd45d0d035841941c1489e5bea46ae7aa68ed2307b0cf0d16091e2e68b5ae1f9a39e3c5f3e93c823ba174d26664b5008928e608ba42e3b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4ff37d08045ebff75123282e22a888879db233bcf18e60add76aeb2da27915204187cf20451ecd784ea442035aa91a3abe19b5343f90e3a1295c591a26e8b959c4c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc4f95fb8dbb0e3c630a4ba158cd7704f84860989c99d265e9df35c06e25de9253de26005ddf882d0b622dc5fccca1e1865a7e50289930bc6c39ea45f31cd0c10d1b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c6a0dd4f3224910600bf825c4f2310affaea72f8d41502da9a84c65f44c908a885eb1f74ba3f849892cc6597755a13931f6a9f31d3ac254e83c60842162cc15c69b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heba2f2b2ea30b25f29f9a5bfe7e95718835c9ac5320891774e0ea503ef79ac37de532db56acbd4d9bc0ba9399ebf2512e342cdbcf22e258c8af6511978eabd703b1e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h537a9ed3f3200b2a97aa0faa7db8fe1d3e34ce4bc3d101ffa7c1096808dd545f8c51203a8d8fc2eb28d2a1a337143e6c9266fd2754bd5e23f56f142c4da2610dec81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbaf54c51b13f7302c490da4ba14de50d142ff285fed616a86b863ef237a2dc5dea19c55cede268f6e39269e3f66234269c91f98c73e2583fb9b9931e34e052074641;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2879e5fbe7c365f290aaefc7ad2d0e0396fe353a443e640ad2f0a1fee15b45c035aa8ca3ae8cc9a27e1a43d070e4e0502ae799f23d1bd33936b85f555568d3d56b81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5fe9f10de59225fb6fe0734891302825add3d5eae5dd991185c359c691bf9ad272b06c7ac21533f78ecc19324884fe85813dd7b25f59672f00754924733b55238993;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71375991c76856a6658ad7554114d9f07f7af15980c9f461c44e31c832b5eee46e90608affb32c2624d8538157ae9ce89540e547ec48cf8a0f177e28162802584118;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f35565e51cb138eef87ccc8fcd988582386a979b2fa4eb65afc83b5efe688742ea5a454bba5c2198186aefe40bd28055926cdb9336f32f3369a2a156b392e67707de;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff6ce1532cd88dc35b2aa5314567667ecd86671b74ef6fc884ed4fc0033cd46248d030748a663b08c6933d3353a0385f0f4df32a03fe66f18e8a9e17031faead5a31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1175899ff04dc10b2ec6fda7814bddb631dfc1ef52f0007e091feac3d17a9063fe4dc6834f8f15e7b40836dff3534703dd7d80aeb8fe1dc03ee1aa39b1646102b7b69;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d59512adebc7d8c324ff797ce0179f8e7254aaacc9b151537c0cb0417c9d7f8fa68755bad5701ab1e1c4d9e3ce63f1f091bb61bc5aee7de7eddca3c0f862a547c1c6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b947fff09ec494f8f60f15a91aaa177bf12b47c8bd8acb5100a988c5a84e35318def6bdfbfd3411057f8ab09b66390d85fe7410e23c319c64ca148c7f19d0e57099;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d5858d1f04a9ba6d58f638b3921a83dbd55c35d7e8588871f833f3b8e9bfcb8faaca68828650e0873ffa3b2f5f0ededfb54c43f22362977a4ce271a488035c8c2b21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h75de69354ee3b47f761874bbe80a1006448ff53d8f5d3b41ce89c959da2a7cd85eb29f619bb8f057f84edf436175317ac5aaeba813e81adde24d063911df547259e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h400b09c2dd5072f16e5617a695ae7c0b2e55a368dc45e72881f50b70d600a844f4bf1f3d164e6456035002a03ce6c3d54a3f0242194ad548206a9308610938691d87;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc17cfc2baea82527b16d837c2e441bcd1b59e7d3d9ecdf6924e362bfb618d81320e24e3b428008fd6a68882abdd8e03e05f5a742c4886767717b8aade277b5cc9313;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3fd021292802270a7d2584222c1a2e9905b03e071f15872bcb5bd0a253b8892e6390a6bd26e0d0debef1be29b1fca6f5e66d53a996bf859d00acb41e7f2d211f56e8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f01bdba1a40d5360b5ad5fceecbf4a0c5c9a32d265ceda470b86d8c177cc75910749f6854940afc6c2cb83e20487acbc3d8af318399ed179c0ad1fd2d32a3b6aeb4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9da3f5f3ce48f3ba96c3066ec26c3c03322d358958a26fef060c412a771ba453fb2a034d8dbfff45a08bb953853569e39c0e8eed4cf28bcf945b9851f2d305dd787;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha108c8667ec4ac848e512263944158e03a61886db9809843a3ae752516b44fcd5aeb508640461f5b96f976333adb2d6fedfed1e1676a3f1e77eae6e1feed0e3139d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16291e30d137baa2915afbf9a8087d4ae164481784beeb68a2d9bc22ebba2fcc84b3d379232aa5e39ff78da83a8e710b905000ffb60c3aee5f1773073900f0962049d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c88eb203853a789ecc1eb9767692ad3042866e9979f461e4b47b7d03afddc8ddf30d2b2171262e3cd3302bd36fc4009ce422fd48bc11ff1e64d045197bab07f8366;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129e42b51004de540f79b2b0c0df63033fea7759e3334b51bcb7895474ff6dd545ed8fe1b7fd7a0e97ff8f343d40f3a54543525665d57d738ed91eb68c5c9354b5672;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h673fe19a5cd599b55d2015cb6333517ffcb7b87a74c48eae1baa0982710b40ab145167dde4af7c984baaa745eef7b76a9e018055bc038067276d9cae748f08c7c9c2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4c1e8f8d475bbd43dde57f257f6d04e6bb5a15471639b02c9e4485f82d1a77583b704e6f68c6ada2d4fb7e783fa913126b5ee70caf80e5eb174d750f15e2c2a70f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d4310511e3c6733cfedd97297f01381273ddb9dd7c50052115281f729512138ca591f2ad8a5cac21ca51af1d1004803a572e644b167b3fed0be9a2e9cd3cdc0960e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h469fe669a096e342bbeb38b31f5115844f66d0ba2c1155751308371dc7064ac92c3c286fa013abf1f2d9b32079e88c7e9b2e1c84da53ebc2a96e06499bc38d0f6e80;
        #1
        $finish();
    end
endmodule
