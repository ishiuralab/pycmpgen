module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [20:0] src22;
    reg [19:0] src23;
    reg [18:0] src24;
    reg [17:0] src25;
    reg [16:0] src26;
    reg [15:0] src27;
    reg [14:0] src28;
    reg [13:0] src29;
    reg [12:0] src30;
    reg [11:0] src31;
    reg [10:0] src32;
    reg [9:0] src33;
    reg [8:0] src34;
    reg [7:0] src35;
    reg [6:0] src36;
    reg [5:0] src37;
    reg [4:0] src38;
    reg [3:0] src39;
    reg [2:0] src40;
    reg [1:0] src41;
    reg [0:0] src42;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [43:0] srcsum;
    wire [43:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3])<<39) + ((src40[0] + src40[1] + src40[2])<<40) + ((src41[0] + src41[1])<<41) + ((src42[0])<<42);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f78fe0efd272a2ead68707624c0d5f401d12bb1d756d5ea6f0a4b6e3e92fab7e3efe6de47aba43441d3b3842425282f8b479d7c7e0696d600f225f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha46b748df8d6abec1f8cbb55cbebddded058702d37f5499accf026f400bb00238b9ccedc7d2ed30b4f9eda54c69400183a743ea31afc651c5922f775e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e34315d93197af37a49439fbf716a65aba62adb09d1227ead159aa9534e71fe8a1ea421b88d8b24b659a75459415ed7956f0b2f094aaf2e46dc50dc1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habc605c42d05d939393296214e14fe6e52e59096844cb7a47fc1b669ffb2971c1e44b7ebb2b113193a07f8fb559bcf91f9b94f8e7517ad8f3341a6965;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47da1b5a165d8b9108c89e717c0e690a8fee356e53b58b5db353c8519d00cdfe435f87c9f917127b1af354ae58ed09354fc06a7f31684eee3cd257b24;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb14330f069a7a865ec6efbc8fac1678363fa7d45091aa29d68ecda8b0d0331f10a78e2a67f4e2a2f296701c395f9972ee964f1bfe48cab1e9efb4a70;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1aeed8ddd08fcb6dabb471df96518dc82b1e99fda4be8b9a58e86486813187159d943844d8039d02ae64b0a7ccabfda9137d50813a17b76c0f186e57b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ff695a85b6b1b37d50de1e97ca7350513ef78c41a549617a56b20496acd61d9769c0a604ccca214aba8ba101d812eb7fca31544725ec25fc2d7791f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b2d1445409910f66c3d3a5348b6bf0dd6c96b951432f426d47a8031229ee4607b1baac4f7bf50efd4b217360371386f019a39d177da6b893753d7252;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a3dc6e68bb7c3aac35c86fd7d2df8032a69ada199101da57f7a8ae33ef638c8eafb474556e3f61bd0af60a3a4b8d0f84185954d2a2b1abb01ee99748;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbc08d4b7d1437cca2b0cefdc1aaaddb23fdb62d5a4cd69b89c5e1b2faa707081b480f61f7e619e14b3ac80ff48c77173edc3db11c662281a476cbe18;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h677bab747cc64e83ffb6e9ef7050e4b986ebd06e1fe2210fb75693723f11490a7907c02a16ab5a91aebce7ff1a4c4b57bfbd67821e79dd6970499f100;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf2213ae95681b356c0eefcdfe1ec20b70118e721c84d200db239337b998c522e71f4163a31b4adcc9cbacc3a547b485b8319dcbd0b28343dc38eb587;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c9db631ce94b2aa7e78f2835241c85f59fe1394da3b1507c0ed610e80f16bf3211aed7cd7b759a0e0afd698a1494494bbfa9a4cce591dc051eef2503;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39fa4824272879c202c5c9971ee367230ef85011fedbaf5555a5f35f91d8471955bc5d834f5815b062e617e5c48c99d9b8d42923cd3075c979b9d0964;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e1274c8f4fa76f32f9d41becc6987228bd06eb4e8ed90f260774ed371e716d6ec707a0491bf5fc4323edd2611a378004ea04bac8655ae05742ae939c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hccd49ca4d68117113fd4f4fe7a292fdf9c65bf998c07dd4be70f5349e8a8fd53d9683fddc046e3bbb13319034efc10202bdc112554531d592cb04b7d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce584d42d5c348741837a469015e7a68b6d6170b9fdc975193483ea4d08ae1bbe6c19c13f5773ddf85017d9ce881c1050093a4f124ec55a4c11e8b667;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6390a236fe992bd112159a4fa31b96645af560508362bf6a0ce38649738069aa3eed08a23791cc4310c4612a800f1932682aed386110788a6967dfe5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6c6efb816de6cdd992082b7ddf383317ace58729399d486f27c4abeb574f29df2041bc105727734c060face938e723b1f24c9a9239c8aac9848d9c4d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8ef26e3c1a142b6eb42610cd3b4299b41606544143c71f8a300d051f94aebde53b759f4cf03a1bc55eb3158af3afa0dfa1ddc0c95d5efe1239d9ab43;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53f906852e7fca271ddd1db2e8603cbfa7c35a91aea27258df6543db7eec2e92546691d879fd08b3e2016e831d8ea8e101e3debb060aba9b93bac9751;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha535601ecbd4e3b9b52029038ddff5c434f7d0629d63b1aa3675fbc06e938a92bc94d57fdc85b868748a3712492c57f6e409c88544c02da52abfb9a65;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f11604edffd99cea81e13d24db39294c1bf69a7dc4ec06df1b52784f1e12b5a37ff838674447206f2ccd2ce9049d5e0eaa25c78779894a4c2f81bc9a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2381ed8438aaac52875feb4c637d409b92aaabd1e17094897fc1a3926860b24b9337fc23781ec780bfc03b37f29a1978ef7f0bb8e8707851cd9801305;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9241135ab6f024f0a1b8f17a6f9f3cd6aacd4491ce2ed6ec355e68d3ce820dd12be18cc158583328b14e4d4076f171951b2d04f5cd4a9630194c3f987;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6d6650c1ac9af8a3faf6c6140eeda77056511b9330486ad4a806ff967633ed82c7cac4e0b0385f8f3a12af126d0f120b4517ef976c6658ce943f210e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a088fcf88b863bb528fc2ac3f3e0ca8b4480250e1732fe7b2e140afcf6ca810d29e25267e8e118670e21eda923f8a180b2502da2cec95e7d448cbdd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h519c1c72559c69c31bfffd041c97efdac427a92f69d21d107677d6cddd0c702bb74b6ef7c5fc5cdaaa3d9d10876de2e2ed37f89f57bdc73d63ba10885;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heed8cc6198243613d5fdd84769af335b3c1c629fe5c1492332f32c58876d59b71c1655517338e51a40450e5ae905b79b7dfc39cb088b3b24f2c412dd8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9ee3ba8053291c43b2555ce60266644bd7aedf2119d833497d728846efbc8f336dc3e68768d29b6756183bb8323fe3b06a1780fccf03af059f39e3c6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67c0f59e558467dac7aa4f7e3471a871e719fcb9f1fb13c1d7dc5596e91707d498f09d3709947b804179ee40101b63001e3dc791482f539823b38668a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf19b755f5dc1d93adefcd29fec65c27082ff89241676096ee9b0a1ce5a2782b93d3e7f37c7493405616bbfc2f34f62a6bb055c26eccd1e4f6b3181c8c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60afcdc7dead924da11b3169ddb6b634a18e417b661511161868f1f779e7ec3c84889867b4c10bd9b19eb6d20c982f25f971e4b246133fa5a149f365;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d608d4339cba204232f940eb7df6c4f4da40965763cac634e842924847298c1d0aa2fff9c675ca37edc72de903c98f47e10d6836e104dee2daad738a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb513ae88ec870b8c6d898cd6af10317e79d54685dac30ce5a88c8cd247cdbecf2dc715ac15ce99b104032858e1d6a39a6d386a7d90f19f0277096f831;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3dd7cd1081fd5ec2134983e64fb7a294ff34f3018cf72cdd60eb905e36dbba8e4c6a7e5e6ed38c5c3764fff82bb51ac96723987ead458c1c99156c997;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52020627ebf39e90afa5ba5cad329bb864259ed8cc7931d7b82cb509e82f5eb99178848e5bef82327eacd2840903471dcfc3e51ac2d719a1d484270a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdd3c6067dd408b23917bfbfa35958043872479924d604129322e45ad9814b411c920f5c7f41302edc4dec8e36c2c00b75ac32e34e02d3dfc633fa710;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa7ac8c0e8bedceaadcabfad7651ee67ed795eb40bacc03d857319651fd7dc152d486d897cd416fd0580663b0b6dcce196d6bfb23b56a3b7d1e771872;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30a3fda934cc04b494c307e4aa396da393541818ac67e702e904830abd29969b15281a763013a310c7e7af67b1af2f15066cc7cc52f0efdb2683fac57;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d27379a6bbd1cc0df068db20383cce4acb34e45888108d2cb654f0b780478a92d9a50d25106674f072fd9be5831eb1a8d8a1f33c29acae4bf8342019;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5bac935de634c952711be9794ea20148c38738ea09765f5548e9d8b435613e18c14f0c5fdbee5aa0a7921f927a2011626e1d850d05dc3a169a7a9772;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5be61966ec630caa7aa769de343179248355479ef47d12d4400c51eb5ff116f528597aa556f5b2deae390039dd6ef0e8e3b576165e1ae133fd855242;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h839f16e27011dd16fbc92aedefabec5af1e08b3858ed8c68c77d9e900eb4c0bc0ff7ec1c12e0ab64a38331b8315c64d95294e239bb9cbd9054defb43b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfcf5049a6b15351d204517d116adcedcb11dfc083e4fba5c06879952a41d4463a4a956e12cfd7ac9a4e721c6b54060284b91177c50d8f80352e2c1405;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha57fd26279ca3893a5b6ae899e983755f28c38b6dfad2d4904197b3c7eff34c513fa5027f8ec4acf7688475096b097f5fd9d0d40dee1e110d3cce731;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29e064cc11db45f6bac01965a434599ea5b03b3664ef315fb27ee5472015662808d753e1906a69584b27a6a43892c94f5d52500a0372c824be54f385d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ddaf826e0a156c16476ca6382e6b1454196a0a85cdb4f3c39c5a05bba9532c6087b809d8ba1f19e5228cdac7e5d2d3579e994436a842c0d1ad46102e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbfbc0e141ce1ee0cee552922bdab09d277574b3bd00d0ec391d142367922b0086354fafac57775b5e1108b2196e89d9679f01a52af0518dbd31a856a7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1833eb002ef361ae90a4b2fc12ec34d28a5d57822e104696b4a68b88d81e4eebc7f7fbcb8861ee6b6e8c2cccdf7cb452e1a05caed248fbbb1f4665008;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h957e5fb624ad6cbc6daa469c0b80130fa7f02eac05c2d02ff95864fe3b6692a54658e04a7b2487183faf3bf5802c0091df79aff039de84f140959b986;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38aa13b0c0fc7d17b1c04b90b057aee04912aa677b2a4f51c149d89857836b0c5da301ca1e1d782d29f77dd41fb7bb674148e0b59339cf9a8815c35e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4fdafb34e242f6588f4bd9ef45996cbb9fc964041b4be9c7e8dde030192cec89149e1c7816f4b9b6ce6dc52c464116b607c3ada784f05f1c54163bb5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1498caaacaefcdd66cc2e199d6d18c31b41df4826a314cf8fedffe4c2f2ec811f9aaa5943da162a4406ea27f85f7f40c9469b8a0fb1ae6a00ebe85bd4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d37246b86e554be4d22780f50c90f804ba7d6f3c4a711da18192bde8bba40e15f4e6d33bca9780643dabf5bc3367f355668a7dd51fbcac5db24c5cd9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c78d71dcfdc60f3dfeba6cc9bb49344d1b3f5f230b7793e4a1c0a3f3160b6c17ebb73796c44d9cdb2b3789e97e7b4aa6ec761aea372260e092b189d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e206c83a6445e2ba81bbdc1fec23456c53f3fa8fc0b0551db57815279639548113a11ca964ed4cc58d4e96f1762a782829d6607d804dcef32f82765e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc104b354d45081ce516b09b670cc5284c8ff9416104098939910de8d25f9d32d3ce52b8046536290d285ae7d02b2e0ab178748c42c17d1e920c8bda00;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5379a5d425f154b601a7899ed064ae325471060f5ffb299475e11d1de6e159cb261066ae108b1921505d47c9146fdc7f760291ba8e2867795f07d53ee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h811ae21a0e795c21b1cdacea08e92110e5dd51a5610de6c7a0faecc87b07daabe2d3fd3f14e8c452775b560156d82caed836a5e2818c6aec05990a33d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e233a7aa68c80c0337e54e178b1704970f19b738311a142bba7b15742ff91fb75593ca905a9c6ea00bb88a1003be9ec99784463ae278eecfa3779404;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcd44771995ae22238d0b79dcbf9efb4ada2a8cb706a3790f23dcc5b30b799f2702f5933de1af52b29ba42614c4cf943170d5ee2ee52cc07f2d12477b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba1b5d89fb8fd95cc62514a951d3dd048d19480ac52e007a123c3c95a92d8d095ff34f791fafbcf3e1170a816ec1b1e9fa585ef051b089e7e02dde826;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e14ba867fc4cdc55249b4961cac8d38fde0d7503dc03095caf9de91bed94941a82984e3f2dedf9e2018aec7e12c684747e10d30ed21c105c17a9223;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2900d9105429b2b9fe813d745976f22e83e8bf0215c9ff4deb719bfe86788f46fa323a0bbabe26600441b0a0e021597e60f79f634fc636829bdbb8ed5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h412b234f2ebeda276374ee847aafaa4399aebe7b7ae4304c506175f4160fae476fd0123d3c1583d0fd3d3cd9d598fc9faba9c18a9e28b64aaff6a6685;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b5f9564d1d39a1508d916de52ab42b523bd6aca3606966a745b20727a4f5af6b77249973d07966280de8ec07a7d82c5c5924f268b07084f2c92e470b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7fd221c4dad6685b9654114feac944967611efcf60199645f2527e17974560bb631cd868d95f3e8cd250c6777f688ff563cc279c463e305e787748da5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24a3bf1261f2c0d1f64bd99422b2598e9213ae8a3af3ad6549e07ffbb39e16001294e5e320c6c2ea21c59483dd30d9b9bac847109388153b2054430a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d37d8b51ec65e15be3034d19d9aa21b85781caed3b66d52aa0ff4521ec635a0d96a85b6053891e54e1cf63fe0caa9b896d363af194b361e55015766d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f2472fe5bbc9a477daf6033bc749373d45121b1504eefb9a6649732e6f186b4bdea2149e89d46de681af6b77c6650fe923f7fb6c8ff2ffb25742ebfe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34a54ce36c13394da463fe41bca8d0f1785a324792073283f86799d714cf993dd0a44f6ca938ac7018bf846b6caea3c60dbcc239e9bac08f53f59a5d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6be7661d0e270f87ad8d0daae341fd0aa1f6760d261abb7506566fdec6323f45b6584892c50dbb4b3cdec7872a5b12df647277b8b948ff63b56bd2d9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h829810f9b2a0476defa6ce0c71bcfde089cf568f06533de93b009c296e664f533db7a16b16db2df652adddcc1ac5651855981525235efb58c0b3f8833;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h353dc32a60ce71c30f74ced07379630ce51a5bb0e8c3feddded8727bb2ff831328aacd08eda87def4413b68af22fb8d9186a4ccde339ed1bb7987dd03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bf089b3efb5148cd51cf675598bb8098565656541244e50bb669824a13fba1cfa427d9039aa9d46ce3b1d2e4004a305bf5e61a0e3d84d4944bc2477a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0c7dc6e9aa2e92f07dc73e84a5047441622afe7c8f7aa2493f6386bd6dfb5154cb28b9517489bd7743223ef7f37685beed2a5f3fb0b65f5d910a7ef6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he144cba62685eb187741e73e1b1848307f5762f33c020507235428c7755f2bbc48460b5b5aff4b6219ea8b41c396a5e633b8a6e52974af37e75970d88;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec111b30cfa53d6ea8d0b993b29f43c7e0113bd10ea52af0997f82ec0fdff6c764a29c3ca25ece8972abf2c91662861a01280337c12006b1bdc543bb6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h724b4e810dc6a3cce806c90e63573f7ba8ffa24890ed42febdb29d3515aaeaf9743e460236c481c91a1ca430f677fb4d0909195e857ea68dc98930398;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fb7978cedaa3417326c36ef595d5cef8ad19d544c67d02dd2c65ebfc55d2939c5c66687926821bedffd3b1ca80645c172e845889e640358333c09e2c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h488f5fde2b234e696326d7e70c8f8ba2f36c9a7e05505f21362fdd0917e56d28d33a629e4071f33d5a28354245a0d15366af54109fe702bd3f0f6c46a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf67dc1a3e904a6dce6240a558892679b63b15769a7b56017d523b79659770570ada019e1e91ce1cf222367774dfd01fafb1b218c49bac049350916ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79c7f3bf276980131c14bd0d5919212876023530bb73c3f167fa4ee96af8dcda9a6b2e958dccfe1fb04e2a40c10b4f72e6780aa76db8dd2d43ec6af47;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5682f6a39b8a490fef00773ea1eaf9231ae904e627466a51802e38521671ae97265ffce811c9e4e37366b4806a155ad92f29ed9379290bfa14ffdf31a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90d7aa0bb8f4f4fbfc64859e3a65fe7fef300d95037378b3276ff2afa05e0193de1c03f0f8d4610b695e7b71618163aa8a224a49852e2790200f52eba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3e64a0de06df02d04925e898a64cbe417f91ebe7777dfce74043a58d725c994694ff8bd245c81b2a011c0cb342d7eabe06f94a4088342e5cdeaf676b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f9380b6ddccb1af8721e96660ebe73b5bdd0775024abcaa733f985199a1fda48a3783ce1fdec857eac764c6e016a47ad62dc9efaf9964a7b109b7e67;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee475b1280723d616c13eb12d4d9ce442726cf5e8ff0ffa7656d6d19881bece201df0f93a26733a7c0724b9c5c1901592dcb943ce1085a8d3c348e4d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61b8d67e02d9663e1456ea03dd40216e84ba1e5ea56e8636c7e8f4cc9e8801a1c30040038f0117e3f229c67d072bba51af7c48339776bc9b6d95a7f3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfed6ade178e1ea3b878c156de95c018c188878da3d83e5283017b516733495524867801b96f51897a616ceb76b1c5c6de0629f1f5692223155649c186;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcaa392d2a626d78b5848d1765cee550758657b72f4ea41b6f5832093fe3981d16c7c16894e50ba069e607f39b024d9e3b5c3f5a288f9f474614045ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h493b43c581b0f2a84fbd0b33d7fed276a82e1316840856bcefdc45ad08fa19bee2b78de6cfa9f9bddb497af8f0ec381208e1da0e125b0e5dccbbee431;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2bd0e289cf4be00faefe8be3c30b144b5f0aa65392db9ca01fb47e8fa3297b797ca816e227d0c3017d44e3770e1d461b559fbe7b1fedf2744b5aeec1b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99efaad5b8670a29d73e4b88480fa5df8d891ddbb7f122b3a07af8add109051fc88b51378a76aeb267fff5b74bc8ef6c9fb8e2550e5c2d18bd0855fb3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40f71e1a2f5f7d7b640ab34dd4613c4117e0d0aec9dba30b8f9bfc8aadba6f50f7ba93c464720a422a73f5189b3b528d7478b946cd63a3a1411a2ca61;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ffeec6851a075369091df4f4b5d14a1c8d39691cedcf6eaa80b128abbd44e9974910819934b0c6356fccc659001f86f038895318bea0b52c701ffb29;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a1045e422895675bb8b8249de088a3b891d9501890ef1921c7679328337a314cade9bf40e0039858e4067582edc0a7931cb8283842dac837673fd17f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28d6b209f2863d544c446d2d10c2a3ba3d626a04480708963b93693925add38b707654aeb79203e1f3b73c53c323d717eae8e5187224483a7c45454d9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa49b1673cb2b9eefde3a8a37811f569d4bfd7f1665048cb28cece5f380733a91965987e0059ccf4ab590d23e1178b7a2b9f321473a42df3403236ed9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a0bb7758bf1de7f956ef128b2d26c742f512d9a3b65d122457cc08115bc31a3352c683cffe4e07c778f1d5b6d326d1af4fbfa24e51c38e72662fe485;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72c3b7b9491395e75c2ccedf2c19c5a2d9f3249d5d30c5b7549590a6d064c0d0722f1189222a2abbb433df1c28b17d7c84321f28cbfec9383695781c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5214e80a65b3934bdaf6742d50d91bc82c31340aecd35cb090365f49d54f32383ab03d24a2f81cc92069b670e99a063a1f8adaa8c18d62e1b1e1ba85c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd843f225516161ce7523c240033c8b4aa20ce86e67f91e3088121154d520d9580899bae1d1d624f4a98bbb769bfd79d168f1c6e79d749a36ed0dd3aba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97d3188109a41d2b3161d6aafb205c695ab35b8ece94017225dd0bb2f63e74528e27be1708bf71349109180022bbf603555d7f52462cfd66fa665096;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41360f9aa27d88e860bfda1a27adf05e196ce773ec79d96161ab77e882fdd66d2f5ea414f51402242535ec192ec46ccd7d781acf217f6d5edb9be3113;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9add5b16289b911c3e531e2288ee490049452095152b80e0bcdff35a8aac89590e6e26e5e9cf2cb192c3541ab4a662885019044be70630f06db9d587;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8c88b8750d05dd75e403d936fdc597788a18c2aa11f7e8f9a206a11c6bb82c9fc58c3549e431c73d09f1ed4f1fe36cb53e550af4de4f561e036b5092;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3858e3705c368d70a450bba49dd6752a62989e0c53421f76381b90abe92b21f46a5a0c002a2089508f00731777aa1b9ef7ea02ab99ee5410232550c4c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedba64779eb48eda07b35d5a59c775b200970086e34f0d0a41a4d6167762ce6106feb64dd784cad6b0484800429e4eada9e9a0b7e5e3d457fcafbd0c9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce47d638205cefa10d0d895a58101108e7544875a17630eb711248cedee17fd95d9302e69b2ad6e0ff76bb6af78ba45d308d22461e8dede80149058e2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha98baa856342195bac06bcf1e3cf457fa8b06dcc777c78f473d47ac15d1b6ced5a03b1e577e4d1c8566ef63bafeab7c5664c3a9446ad8ea64104bad8e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27bae43203db9746d939299dedd926f83c04760fbb24f9fbc2e1001dceb3891f1b5257296a546956f9549a0bf3cf649e0f098a3a4ea0a971ae4bc8fb5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ecc9ac6d330532dd431187cf493405d26ff09d7d5c6ce5dc5c8dadb35db5b79a79d138f3214e02b2b0992878efa0378fadd16b1f7d661e961b120d47;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79b768a9cc3ffdd7b47ac9889bd74c39e5d7726f3e29d7cb8335cedeb5da15581df41fa0eb7b0a4aa15a1ca8f410870e7282ad5826603f4d9d6ee88c2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf265a3e70532d8b0579e10cdbbc808f93b1b43a3c6a618d884212a1f09d8886b52c91b67c537b8d145282685091b0e466e9207870c4841a2d9515c9e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1963b8fdff04b9357d0291561d18c65f49c0138188a09231a04bd12089ee118f3112a65718c242bee2d2e27042e062b53814cd10602303d340e6ff781;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66bfaa8e37ef019a61f625562683850bf689ae7a13a96bb0dfca150e4ef063c38263aabfc5e08e929253c40188748be2a0d308a5f8cc4eb101f578353;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6f23b8591985fd8ccf491bcaeeec991ff79e0602b5a10097349df207352ca92ccdc7e78d872f78a62a820ad0c8efd31e74521f2f689d590a629f41d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b13fb25e0e28a8eda1df018474605e498bffb6a0811b2fbe9a5ca8601172226472590b036a662690846d3adba2cdf4a0f6ece4ee0015dfda4b31871a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bb622f5f4209dc0923b1da8a75487990c5db5a65b7dc8622262286bad28f268cd2504f5d73aaf1ab7046dfcce80c923ef89f2d52e91e599894195fd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had85f9002ef94748e3f36e06db8326afeee1b3c2258c00bdd1d45a6f06a96583e8ab3a170f263a265ef30aff9a16f8ae2dd0b3330f46952c89457d506;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5bdd69e7ffba9fddf3aacb95d4ebc5011ad7e7743ff12e26ffc1d87730dd87c81145475891dd8e0e124b4de95e1428f0a95f501f7785dfc18d688abd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7eb0f5206dcb5b0f09a7af724012db0ac7fb04602d52dac27a8b9dafecb60489f77f9a1700ced288e1e10433741abe5427ae433dac0b54333192eeba8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34524ca9b22c4a4852f393365b0a85f468c3524386a6c741800893e20dc76f81a6d9a35441462d6d8ad2327cf1c30dcca29bf90d00b115ba57684c283;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef20990ceca0669e1605e17801b9cd8eab8518f7cd4feb84ffd08a0e92d2b7062b0de4218f735b7e8d73cf69f25a4b71d535203d4c07ae863d3399704;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb027f9785125354aa84b7d5616e1bc95af8cb4c234a7deac28906d25ce4eecfe1b0b75c6157a5cc4fb0366535578667b3f4825489ac44a764957cee78;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfbe0a642b6aadcfbca69a4058da09e37e7d66ab4c3f96606367e151d94cbbfcb84cc9441adbbb0aa8d5dd3a4c4bf3fd25d05b4d23cf157b4a3a85932d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2153710b3b499c1dd538dfe904494e2fc30dac9cb5acc6684ee9ce445c155fd359f80d6712755e0d12c632c26c1d58ed2581c91ae702cc0cba03adb71;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c46f9807088204e0f7f008f03f4d86731159f5a9ffbcf320baf194ca95a92e6e00a7ba9fd2283308cba985ea9b553bce9d3790fa03a4c07e61ed7db6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4910874a49bc734b0311dc3bc882374dba3cb357bb694b2ddeca1e38b5a303d0b404c17533c2a5e2c085e1a00482ddabbb143541f71b3c87ae36b1602;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb024d913db42695c15ef3e4f9d1a948143c8f330e61288bd65381890c1bfddb999f2220b81cd79c3d5c8fbde6b7f33bbf2c991332938da5b3bbd0f45b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5816ca49f5b1ef323aa4cd37d155179109e8810669b2976f2750d2bae196c8c66080634a540841ee24f17bec5a4da4a852f863510a2965ac31fb978f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb46a55e81ff84dd845be626d0ffbf50677de9d63b1cec04e3db737426cb44822ef8d277dca8e0a91d65f696cb467fb5e2af85cda5675f7a3d4fb50768;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbba0249f789584b9247d5ff88e4284ff31500a1ffba808c10fa6b47d07a52cd80ecad63467c32fc1442ee926aff401aa836f7acafaa4840bd7bfd8a02;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d1b9607a90762be6593f65f88bb6f7fa83087d5964b58b6e79b64a173e39715c6d0b6b3d87d3ff6791a8a6247e1f8672daa7671ee00f03a38d80f7d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c128fee12038b0fa3615b32c8d1538628058810585a3ee9149b55074783c0bcaea9b3a4ea243e36d422ab2e90494f6f8e99bc85bba1fedae1b1ca7b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52ffa3492891de82029a0c681e698bb9ab19f3ab162092069189cca99c3b2d7f0c44402df6cc26283a43b7a60b4ea4586007bd88eb541e30fee0a3fe3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9771f48f4f98cd9e58677d2071f31179fea6ebea0f6f062f8233595b847cbf6f51a0a0f698c6883a3f59e34314e00056a15da68c7632e90c3a35ef74a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1503b1e047490df2f7e3f13a242901fb1be783ee187f2a0b5e2d123861b9338c22f7e15fe7234186f9597abc73e09d209f8d4170a5bf83b2e7b70e247;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h744e66bdcbffed9ea20d4568cc790ed73b7a934a4175fff875edb465e89123315d1568178812cc69e2721dbc2ea733a96e004b214ba282f1a61064958;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb2d122a712f05b8b3536066d48c4b84d99c321b96ec93636c4be365a3bc0eb6b4869af5d5a5d76410b0f54d9e289a16b292b7fc2c684f351b99bae4c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15d438db47ddff4bc188ef473e6f782f8b1c65f34fb202f2aac814eeb4684ae3c776ccc3da3a488c0d930d2738330f85aa3399dc27825150be6a904e0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd70882329cd14c812b1c0935f99578f6a7a23026a1c729abc3ac5d96be49b13422027b039e75162cff1867a1b0c0e1fa917d44867bbd5d33c64f4b8f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66ba46dbea77bc011ae9fb732a181f31b9d8a8cb838887eff883ff341a8a69722970dbe9b19262afbae8130c24f30471e4ed550cd8e25cdba368ac88d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb51612fdf9a4914a061541ba5f45f9e6ebbbcf85d003845cfc1c868eaece614eb2c1b0a54310b3ba50318952d8d9cc41c65b1ac1a47afe5d4c12470bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46ae724952b98a6feb6686abbff343e3656a227b21948e63eeb344d7f3deb49394ae51ecce07e0efb6ce6e51abd683e4bfe27291cabb3ccc1f962bd59;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86a1faa25dbd3096868722c76187d6cc049f80fde931185e9512d02b5de2f9cf29d306f30bc7e9edd2933287e2b87d54a34ebe875589a713db33849df;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83915898b809c53b557383a6a9e98b96780e797ecbfccd332b3dee598bde5787e1c599d7624119864f31cbd3e8d3bdbb6cda27093068ddef4c7161fd1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75622f775b66925fc96868c113df2d6616f248207865ac4cab4497478eadaa2f84bb831aa9e73d4e4a1ff64247e846b2c9709ee5928c89ea717285d99;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h767c5bf6a314501a75a39f752f9465722e8ffd47b23460e588ce2577a70e8d6c7fb378c32dc3ae8f9965b6c3c2a82398c91cead902559f9cc5e5f1419;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb46a07dd102f22460bd57e5f5e4ed6f98b955b559d1929cc708aac94b01ecc619815c012bf458d90a9b0f67b57faad0aeae64eee6df549ccade1342e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf9d25a81be64a3ec31b2856ba40893238406927946feb124553ee7baa60f1d3a60fbd1dae67a418634b19a2029962fe7df3193c86f5fe4734529a2b9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf57c2173d24df84781dc171aa46075aa4dbba96ceb92f7ddeec7ba20c3bb1741c0320543c9768c4576d334c6a682173cb16264642369b23dae6ec351;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0da60df8f956e76eb047421c30ac986c4481635c86a4c00d99346a1e94b6e52da510db7ae05a412b67b4dd5298fea399084cee62b35be1a7223df57b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7342b036e5eeb6a67e5da5d4bae7dc6a7c8200f71d1003431dddbc3fcaedffe27a9e0408b43e4ee6884b4c58a5079030baccd35b50318ec32ac47e85;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9936120a3ca8b1598a44226b8e9642ed6523cc671893b111743dff3ed48b94cbf85152cc4b39454883f7282cc21c6480db715216cea6334a41105fe62;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac3c82debb11dfc7bb84e04669307186ca9e05f6fceeb1ca938d56cbcc736c6034e0753645ce98b1a8ca36db63ff029512002c01e7b24f9078337bf32;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff8ab2ff996be649155d7e98e34d57a706949d3caf684181482bf57e3e794a15e0f0ab38a8f0bb166b4b06b7f7ad1020db994a7651d1fe5bab01cb1cc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39dafe055428a44110a6039e3827fa246a256dc9c17e2485f29192cc86c74646104e0f52a93f34d215a2a2ed477e7489a296d33ec7c9d6408692d638f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42bb16cdb1dab95298bcb274c8ecdbc6ed9587b445f9996e0990dfb63c38945cb4d4cf916dbc683864a2a4033ca4b0bf7b1d435b6ffed6a28dabdbb8a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28403bde0d9adf32c7d77da0f70c37ebf487059a564d99a8818424b9157fda3e02bdb6d119148693f0e10a567ce71e4eb08e16b4f7ec9ec47d49c17f6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7fbe347797ecc5b5b6e46af8d7cebb7f0cb47307da78839ee8096e437df1b38c675f3cee1b0e74ea35de53b37d50b4df9f3d02095204c5a48ef17be04;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8f783f41a71de42b2dd772c380e8fde663ce77cb28ea7f2d0a6e0bf6b598c34581c3fc0d50e5f1c2f829db380ea5d5d50e3ce23cfa06928557d9be83;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c817d0ffeaf465f494e51a91d83f046c56c7ee4a750b6e91bbcc9feb78e3a35173f72bc19cb0d41302b25a9d26472b3bdfb2f1ce5282aea3fbabf032;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbac23dcedbe913509a0bd44a04932102fa7941751776eebeb5e2d68eda1903f8aa91d3fcf172a37d251f019f59f16c823529e7d221eab9ba6bfc6febd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25880f498a6fc0e3826a617a46b976fbc933c4e57631242444947addb3e6e5d4d23ff822f0b3c2b1ae8dbb936373a68bb92a3b64d7afc0cccb55d2557;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb38fd044f37f90d6f157dd7a385c809440d4aecae77688ce2e4cd7534fb3d724e09bd06ec0bf60aa20110d8cde9f2e07e18151ef86d9f21fb1f017309;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b04a125b33c265df6e9de03977b348d17958c0ca74abee0390fbcec37758d0173f7ab771ac46d0c7d8cb7aa70a1ad780602c07a285962043f3d419f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27f34c02c22d691f8feaeebdf31d1f81ee3277d736a6051dcb50ef8abf8dca689a41df9d53450934c8dd6b371c3e59df6fd5443637f1a6a8ed65cedb3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9447130461dad068bd8718463bbd175c8991d3e7eb7b140d092611b60b75991be6de09450c6bf0b4feb7ea2cef8acb0d140d217a0842338e953161df;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99252b19da91a093ac2904ba8d99c328ec373b0186e82dba43697f8c839a4d3d0adcb4dd2c96d4345fb6d97325de5d61fafa21d915d298b02661eeeaf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f5da42e96b15b9f9b348e5e720a28dc8d66f6ce226e79a33c255234601ca51678900d2c6587f9a18a54afa7fdfad0b1357db751e935e1156f1e23527;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he438c80e78174c5e4be22d0ae12bc6ac7f2c7f0fdd5e9eb946bbbd1b7f7818c8dc181628594b92065502e6b828ecf001a9060fb17743f5c8ca1c02967;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63b45a02d8ca94e47fc4bee0278bb80c3db6e7b3ae8140fbd6375476298bf4d5a1e568c3c3d6301242509ad998f87eb8f732c83bc8ccd5249015ed9ad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49280d4f1cf807a8bae4c33de901c7938fcd992bf2a511dce818cf4fc84691a9c7e784f250d17c90ae95b8f16651c82cf854b1f87d5ff783f849515ab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf249cd9adbbe76d25fbed6b7a22603e9049943ece09f93debad3b0504a6e514b967919b921e524f2645d5503d1ba3ffa696c38c179344b3146a280cb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c82b17e000d0140b618dce4bd9e03e80dcf2818c51a770de277cddb3ec918cd6b1c0a9fe0e0fed7475deb3d24ec35d5283ba422162fd0885a8866abc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d4f088edebdfdc600062e1980d177b4de0ba2927ca0771798ba9ba632b35be0e28b9ab1e1425fa69876295936703d20c6bf58455ff94cfebe7c533f0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8dac6537c43a6bab275f888e45430961317a7e2d27144022999f064e7c88c98d1cfebb3caacff7c99d83167ffd2477b15ee66c5c12c9eec29e0df247e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9edf65bdae0ab2eef8bd8d14dbf69e0e6419a8f7d16c446e264d95bfc25845fd9f39d748183110ea54b98787bbd6b9719b699eddf0506ea94ad94147f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd85e60166dbace60a19d6f31ce7d1b2947f42047648fc3056b4f00537c38ed732caf314d22b62c69b7bbcf06828c025b0606856b5e4d2f01c530f1cdf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7028c4da8df48c74cbcfe7536d856bd2dacd0268d90eaf59cd4613099cd192996a26d8be88587d84096ebd65e4aa7bc41ee079d951a09ad784ebc582;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7dda51be1758c45f9330eeba757f6dd913d503fcd4136d250fbb5c470a1714d4805b02fae07345397078d2a75a85d91f2801d6182496f09f7ff7f12cf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he85e0ab5b93862355ed6185b1fef8848cd5c826ccc39e80d7fb4a207fe33204d7fbe4892833a610f1ea0a37746949df9f137ad0917203fe6ec18c6b6f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47e8186046a590d0ec3b74596068c47b76dbc571a256f0e4e6205b3ecd2ba35bc2d132039b95dafa3d76bdaa4e2c6995f08eef2b21e419f8d314cec90;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h883d715d88715178f3f5d2475c4fd4f5e84e1901c6e92748b054d025162245d2276c80d7063202b2f32b260b54329d172fc7fac9f46ff52ca34e43679;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a766d502616902dc348ad12c1d3a9bd5abd95092b2c8f61eaa9d8a8c85593da2a0a5bc341b249e56d925bd3361a5ac71f37b49ce246110ebcfe7a58d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2610a684989c29b64b9085d7451425e9593582fbf030e14f723fe66ed586ecbe6bfe6a7473a417fb2a4cbfd169bd5686d66b5c300d49df54b55c219fa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h905dd5ac57f28b66b64798a42690634a238d272bb0f05f2b437338e43c93f4b532d6ec3f713abc7ee69d4e57f077a9583dd59ac6d199a9ac1e48c2e64;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c100d9db59b37df4035ae46c640d6c0b11e66ae6ae6e54075974957ae2b0d339bb55b07d8d7f84f75bef3eea74c3792f123f0b07b11d95ff1d936a74;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7cd70af691568238841fb427e4c3e599d16f7d40e697eab8fd82b275925d428ff013bdc0808ba69ac00cb20bdddef63b0a19a30c647ce93986a8c549b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fd81320b1c858b54d96cd8d9e5882c87d9bfb3272d54c1a3dda906c59fb5d9b89fc3f9fe17e3a168171325a2d37c2fb62eb354158edd39b249e73fbf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb53de5ebf54829ed7fa50761120a75d189192b968f367fd7405d4d863ce2f4e274c47002e3e96ca863f8b25ec7108c485d11722414804f090038d6a34;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13b20f4789ba99153902d5f9dbf5e3dbf9379f4e3a04558430e103d1673919702a229258fd848b79f4288a5337498e7c6783791e1ed0dfc5b9f341aea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h544b73b82bf7633fadc787125d66f9ca572abc1a2dfa7f7a5da88fc9eff01bde9b54c9cf3f34b8edc33bc67a9f8d1e16c72973579992352e73bf19bb3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h452cd13906f973e5a2c4c18158ddef7d530517387b0e1ebae68c1d09f393e8717d64dcef4fc1b83bc1eda08bda5f544add9538488a435cb7b0d5e47b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32f813fb14eb035f67d441dab67a7f57d01708fc6c6e23a480d010797e031aae17065ee9ebbbcc5ea76b1352d1353cbcb3bb9b28e49f0e47580e5cef5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e7bdf256c7e6d6f3e8a70287260eb80b1a5329db50a8bd0937365433d7fdbe4f1cdfc3f91564f1d40fadd4eac4bc7efac02a4dbeb1c6877414255c1c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcf9ee20820f330b028c966ceb45bf582a5178f9429af3a20eaaa5674e79ce210b5a4215b3835a29eaa9f2bd30942a72b95eb84d7870d4dc21c5deb22;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46bdeed32b3b9d27d3ded1a3e0aebb624b6aa9f5d6da3485e598ed2f4a89b3e169f1d254ec4a2956e9885cff99404cfda6d9caca4f5a13222213dd335;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2841e1ca387cb2612cb362eb8b48072de8d28347b680b54a75e42a0eaaae291f8574207e8f6259e29e56337b5cbdfa1d2ba4b1cdfdcae3241f341beb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8f3ecf951eec901f25caeb1dfd6df68de9a12e89231da675cdaefefd10c2377373d20e92af6fa1470cb39344d3c434c3d059730233fe33893d3efabd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37c8ae1c105b1840c9af8047f08ef4ad786bf171f60d9f272c2bd5fe53904b462252790ce28feba71d0fede9082a9a7fa0918b7d0a1e8431c3fd8a242;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h566c0ad3387b9e8398d49ec0900f7e020dd76c3333b563cf774ba30939080066c21c747624af187813ffbd02576e7a9119f8e03f8e788f2cf06ed2c03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had0307c0bb852879d34b6f7a7dd5861c8a734a151f02a147791d93c36cb8406ebdbd9f0a3e3549096596af092c6376696b53e3e2313747287355de770;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he30eda95234310ed622b3ce95735e0809465cef9cfa85edd818787799332f2f650ced35eae53c5a413dcbafd959563846f03d1c4a0dae59e35631d718;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e68bbc1cc43c5cf2d3c67544530af8c16e5db9e3faa02423590bbc1bddb79eae73eb2a642e27fd2905e15784bab2f5ea385090ec6255afca669d2097;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fc875bdc91a86ecfb34a3f9d38a71146f04d6d9ec5ba7496c6e015d5152f05ed4bdf95d0dcb8b4ebb833b26998eb2850ce636b8f6906e00efae715fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf92fec2800d9c47fe501f880bfed32ffb8e427b494763c2bde8d4857367f7b2a0e1e4b7bc6afc851a1480f45f2531a43a26e1706c8c33dfd4f293f975;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfaf6c68bc8c6dafd6d581b0c3dd6396734e9f7e42e412a2cef9ce4e09d12f430d0c91a26dc6b45f30db62b5d7458b71b161af4286a684b9c8b5b79fde;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea520650b1569e524075ffa2c033464974876eaa9e35d484384c9e4bc95a37ab49770bdb3222db48f18e46d96dd7525e00749ea0f9ccfadc420281fb0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54ff3d5651e2d854b355aab87849adee5d6cee0d55640834d53d486d69f6f2395036b9789e23635f95118a92720508bba55dac23c37e179525109b7ff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bce880cd496b9c735a44c47e812b39c1728a0aff9c7e12df6c9d38762272f00d97ac7db7fb56c1ec2a138acdbf450cba3c6ca812f14bad79038bfa58;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce247a9d0c20945817b9d2177510921f44f7ab6f631ef4961b9a8c99a77c5628f20e30132cae718c7469755d490c6abd38dae9409fef08901f27711b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had4112bf0281c4d00ae7cea8a3b1e8fedfe5b370b8a5d3cd01a90a9d82b492f2dca52f711715ab24a7fc711dc23eb3a8beea0bd57baf07c17da34b417;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he539695b0e5a2ecc38cfdd8eae54d98a637095d977f56117dd0ed3f2e6f12418e9d27775bae1a06b34d5ea196059c5c72f21e213f0fd5c81312e9ed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9c06354464c00800918e59e5d46ef0b6002f9ac08ff4b19a879273286b16c8b532fc10fdb109a5480cb03d0a7dd6f34fcb4376eb5f44a234d75b90c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0900e0d32c2f2186be5d978a743374cdd5cfcef2c8fbe1d6e232d1e3bc0af5e874911892cc7c65519151135d3e452cc08065132222a64fcb7d64fd4b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c736879f8737ad24273d0e8cfb3cd6a81e26ca208baafcfb4c33f0c6ef84c0dd05e0ee5309b334ed95578e98e03d04501ad843633ffcf09ebe9402c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f58f0c2690846f06fd33ea96f45d48cda6167798cb3dc1c8bdb5d16c102fd1cdd33e2455fba6ee214c97f804ba381fa3dd2587047679e4b60f1f01b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f0acd386dd9b79e5f4136ec0a6804b8e87e1720ccd9e0d6d6138a7c62ab45840171cc61a097d59fda68115ad8364eb09db26646947dec22c8b70b7da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d84bdfd1e0d66f1903d764ba3ecfaa921f96468d41ca70f2fec02510be68bb567e5366b6a9593fe36775f34efb43fdc1a66dc94ca0e46f4abea1e1a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf40a633ef280907b4cb79fc5d0c96c1addb120d115afe881f677698a3f2795792f3b52d7263653a55b75837bad4de93d1dfac5de0d8918440bff66db8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd55112522fdbaa4566af897289974816f2f086bfb578cf7ea13f851b38ddb0e670782b711e31d430036528c69384c9bc9ad0315d1669209cd697be0e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a4d2f7506fe2e9dca65d1b5f008951f53b7ac2673e2e485a69a85ecc82cf4d09e3c96342e46d639cf3a2f0a79f00968ce7bcc2181dddfb70a85443ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h359b2a40da7f054284d367e084b3d7c1e35ac6570ccad2f25419f6d07ba285ab0c5f4af60ac25b39923837b1447e45992d20fc4beb531e9de131ee1a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb08ef94b0757cf178800579040a86f535d48a98b79b81ffb66bb912a52fb6e0c18bf196c444bd7ed13cdc1c38cfc5bcc3e937327545b32b94741331ee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h197dd358143e0b7c78b681cbdd110083777e8d1a59b5bd9e4c4d22dd8bf63240acc1e3cd5fa267ffe5731546d5154aaf43bee1bb647662c3450160986;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ce7c0348b0ee7426320e98f2cf58bfdf81b6211963341236301edcd7157a0b2f3fd82dd9b21047eaf74a6ce6f0dc06f494599ae681764e244443bdb8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha45e83bef6605ac55059ea233659f4499cdee3e4913341eb74426b249f852066ffcc2eb2211517f1f333b3aad32e1476d3933fa34c90859ceb5a1d1f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ea9948181c11230f308b41d2df74710fe648ba9549a21b81aa032284a0ac2266deb657e8ef2d3549567deaae52ca80b950418ebbeb9f2a800660231e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb31413f61684088a2ea0f8a052ffbf855dc22b3a80ae291ed56d2f912566617bdb6c8a8ae84c4587adc8f5f0e16a3af7caad6b98ce9d7a77c4728f13f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h430c2f07a757ba77c24f3553639f7b6c2cca9d7608ab7b261026d4f0746bfe67a8822c3f56cd15d4b2dd96f5e3aa1b4f1eb6c38568ad1491ff516f40;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bf84e306cab273b9fdcb5769bf533c585559d33838cc18dd7a219bf4190c99a9ab3f23380d5faf2185d14fbef90da3734771730a5a4debf0b48d609c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8cda675a43f56558ba23410aae529d64b272887983bfd7698f0972fd2db1124e1e80d34866d465405163a4fef98a0e5bb111d16293081fe880384d3a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0ed377461e004a40ba0283d1abfbbd4256fa5f37912fdd4d9a7a8319d88c3652bbbc5b8cbbfd3e8d78c15f693232186cd9b786697fa3ab37eecd1b51;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h625f8f74c49d225b0a7963fa4c8c38d88745a2436282ba3e64e0c5f69d547b29ff50bcb72bdf8979d09acf3d60188724ee7033aada05979cdf6d260d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h130947cc4ea032c60b8444609c880e7fd2b87158f99171001e8d2a96dc4732d9216847da38b61787209e43db0610b649d35a2b96844843d206a8eca74;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1574130dd88e1d99329af63ca296b2be3d405d8e93553dcf5f315599be67e62a21eb635237e54f4e60b8d6aaa976661bd211382dba09a97b6c4b249ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ff4e4c321a4a5149da0cd083fa0a30f33ffe754eb1003d1b975f5e981bbec7b37a896b2b33394081735ac631d3041b596010d6b2d7b516fae82108aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8af045c7385f0879057706775f706efae1304b376a8b55fe198353ddde2a256df706e1015ade62db9d5162d81f3f060bd169d186d5a31b88cb704dca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4bc003acc7298c0325385d2cad63086eb8e44064d57c39b8d1129b53146fad5a2057e405e3d3feeea7c53354478d48c477740aaa8260c4b6bc1da7e0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5cf03b5258d0dcdebfb427009db5810b63a53b4358ae72f6e01b0005e3c04be41a41746838b4466c4b5b58b614729c0a1d556ea792d4d434bb7648e7a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b1a2dd599f6fabd14b58506138e2a553e913298793b24f3fac8a21d87c6d26d052af9201aebce5cdd9d2d7e9f37d75888b0feca5be474ea6b269a168;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12bbe95c079a11f5f5a58de77285ee513f670b800a658647df483549830d7305d75aca68b2fd7f3c217e484671334e4e92c63de8bb1314e031f528abe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92cdf9d2ca024248ab0d798354041c23bf18f0014f1a223fd859a1a81f9703a21d71215485a45ccb635f082e88d1b4603263157c8fa5feee870f3ed1d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d2fbb096773f7b8123e506663b28dcb718bd420e8d8e28f4956ea6aa3d506e418adc29185c460c8f04031838c060136ee4ccc441c0345f8489bb64b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80cd7658f2f1fd66fad46f248d2d907ddaf89360e3376f6bab0577640e4505c6f256f97f0c87fb3681ed88ff310b1fb85c79191a633aacc1934678fb7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5eaee3c4467412a990d4149594e8ebba77d1c1e298d736cac45b32c65adeed28dbd26b46df18253f7e4dd3fc314f0c6a16c5e50deb9d0923562375143;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha16ed64943d0aa3c6bd558bc8a236b60d4626b7b44796447d3b438a0ba506f494c341e855e7d11dc4b01f93657ce67ab782d086a99ebbdd9672ca7023;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d7dd2e47246440512c838479cd378ae8dd9e706fc6118837ac5ca3e59437fe930a96e3c8e5cae8b203a147ba8528924ce863b544c80608eed70d3012;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd502fe92d976193bcb1befaefc3f1333cccfe79dece6af273dc0c5b0c7d12fd4e4e8ee6b3d84d6806171b1a8774fc21598a0463d79c216b289bec7c1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b9965c69f947081ef7a70dd040d2fe685e28ac25b2043f3a9c47681abedc3e1b14e1e7293446d26b399c0db5a779d01697d66db72177f3f0d13114db;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee7900a8ae9d055b476bd900a43ae382255f23ef0c8656592b46cd64499bd11a902f6656a397e975c05b90f50074563ef7ccb62f931d08a2705695775;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9802c083ab2d75ab21bf235c4882f9429f4eecbee2ab187e3b964657d03adcde8536642b47c7eb1265c000a239f247c6ff68b709cfea5cae31197cd3f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5da820a0a147371fa2a455ee9d9c6c8e21e73ae2b8a38ce695da0aa30f472f597023e45f3f489d7e4db41efc874792a8fbdf368de814886e73bd82618;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc24db7638ac99acb1ab5133c4fb0c2122dd866849c0e18e183f7908037dbedfd1cd3d19e3fc57e3e4c7fdcc4e755380769f726f20426367654afd263e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb52cb27b05b5490d814b8368f2877becaec5bd96d41decb8c6cdbb52439ca8cfc62bb07aeed5f7482b1fe86dbd5121671d54ce244f9039580577cf096;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e8828383841cd31fcdc1b996989956ef94f6b35fb598e1e58cdd79826092d886bc08245ad328032aede3a0141ae60cf40b30d2c0ca7b825c99506eb6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2b7caa977866b048e89bb680518acf33566977483c5015ec8f774aa5ae2734bded82be539f839737890f5d4ae20f29c26076d585797a20e5728f1021;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6501f4b22b16f9348e573042de6acc6866a4f94f0ddfd3022a897246535a4aaa70429ab8fc1f4adf0fd1aefc357b7c3cd35f79717c9e6abd31bfcb76;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99acfeaad14029d22129e11436bb2b657a4517559733a876d68fda2a88f645a84ffc25ee79266b7f2652102911b5bbfcf93e1afccb5969233a340f74d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had56bf80be384cb1c4405353f35f2b118225fa8725c6114b2247315e360a0bed3120ad26428fae64f4444cdc51041248152d5f3bc6a28e82aba5e8cd3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6116e421ece89fabd5fa8ba7f527ae8ff9a8ee9f63cb425141b8a615d7ea413cf4f09603e374c7cd279944902e1b265eb04124d5867ca3dcc94d65e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9535e7fa75c67980f61c25f23e80eaa3df567500ffbdca0c8a3b9c6aeecdd213f2b94e23c9c211dbe4b149007ae08b51072081eca427dceb8024b936;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c27f6d5f6dddc1330f15a7a720811790519f3a9cc2de53755b7b8025a0dbf2456902f2a495c26fb43562a4655ce401402a1cb79e459fe40c3ae3c44f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3355f8f5b7e0b698487ee50c416abfc239a63e0809c35229db79e7042340d385412c670409b6b54165055a57aab25c1075eb7a7a800cb5e788601f959;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f3d084247deba3752d69b82b8fda27aa9a94ece552cd080aaff2a1f3a035528147d5512769d5de3208b5ac1ce6511ea3d2bb82162f5d6f330dc0294b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h422430bf31f8df743bebac93d57a29f8aa1d810a889e24f84db002073bb1f6b6b7505abf819b06a89798c895b023a6a424b40edf051fe5868d4199e1d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4aeddd346a486ac3b0b6d63afdc6603e8fa8d20649996d9d9d7cb3a28c769c0f20c71969e259297db84c451861c06e1864b62901751920e5807cbd518;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70ef04cdeb34354e6c6ff03f737738ce7ce4cfaf23afb3469e2302ff0bdb79acd392d01b265ff9d0c4833111765851881a73243185577236590b9d251;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4edff869204d4c961e4a25787b410b9814bb2c9831a7ae94f0ddf2d55be8b12fafeebc8e6cbaf3465ee92d935b283f073e0fcd5f34f8cfddb7528a62;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4193a332ef14edae93bea57736ac1f353da56ef238c58c4cde97eca583b0691b3bbc0db4bfc170da7f30418f6e630ffaeb53b0a0d8c113b020f67ef32;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8a3e22756015a7bd312fad46b2eeb2cbde86106d75c3948fe44540221fe013dde0ec4d6032d8a7a89f63687ee4468e8060a9711308dfec1063b52202;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba534bf9d1b6e0b351c8deb570ba30f406776acc1c4011cc65ee36bc51c1e48ac3382331cda10575a696ae352fb5a587564dad3334fe23b9c58907749;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a79ea082180085abc88f0e4a2cadaf6b87d5d20173afd7281b1d69bce96ae2a664c6e2d17d4d4c8e8bf2f0189e7ef0d728d0080f8d00815de8d882f0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68e5087be7048bbbd2220873c042e8a0522be56f3ff16b0877496f1913a3e78838f9872aa79feb70e2c3df3111689de2c25634c830de6dc064965e24a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he195c51d688dfbbb6f30549b3d8b49cf1f7ec73e4031d54f394c229def4cac4236108e14a792a8b6bdecbd6bcb56b9e677e289c835cde12fde0a340ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa35db8bdede71fcb4eaa09bc5cb54f7b3b2c35e2045585806826a1f9b537bbe9842834ffbf6a4683a62055ba602e8488fea5a5acc55c40cf342deeef;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcbecb4c9d7528f6e326cf58f593a16fd0d8aa7cabb6e0920b1c5c46789ac1796fee5ed4a80edd1314877748ff8299980181979a8820212c5c0b8acc8f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2dcb8a6d43677da9f8dabeea55d0dc396beb4059de12493306ed26d39e87b288fa1b47f30dfd02182cc3991a6f33d133692e1f9238f08a4e9e30231a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39e5b121ffadc582ea3b5550fbe8baf0a7e01de94db9648ec97cc921baddf112f517dd4c48472d837120c6b35d5d5527707b5eee2d456ca19a898cf82;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c3782198bb45fc27d22dad976623d1dfcd0a37f995c48f8682ed38526f369502eefa463528b6682582401ac30f1fe1550ae117ab4445826ef63c3520;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4de606c757b2b72102333dfd21b151a4ebebc951e2236bd5edd6241254c25b48a14304ad6999bbb5597fb7ddc5d1449d175527ecd9633406811b5b7ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7062c7176e96b94790c9f733b1af4eb8c68cee70103fbb258ef1f0fa62461b9bd397e9ae7382a5649cb7e228f7c7508a06ce5a62e72100a17559cf600;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64d4b460e3c2bad8ed2d59bf0a3db1562697d24466b81028b61ac2f7b8845256d8090da800e4d389c6d4892c40beacb2edc22719fcfe9dec2fd0ccfd4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haca4da614771dd1da494c20498f11f50cc2b4f041524c7bb753142eebc927708f8ff37bf278ca415507eacbe760f5b835c22e3b1a636475942667c724;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bf3c30b99ecbd012ea71afa17adcfa207a3e8337c1b97f38229d9a18fae2e61459a8328b3d11214059a2e1dfc3ee05ce9c62faafed03893f2b68a51a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd635d30d10d487ad3ff844669971bcebbc2ff082ef4becbf3a6e189bdb5f65d17dc3f1d88281ac20a4d00a9fb72479691e7a16957f2596829638725ca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12628681a3024f0c06c1520cc205b0e0efb27c23ec50f9543c592528cddbe0a4d6a2f025e6c46e04c7c87b3bfb72dc959c632e9123743dfa0eae6b391;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11d6d9448563681bf661611c79d11b95951e021cd64df20f7882c171e48b77723e6bb8d4f6df7c2888c2e657aa761ac61f17e6ba1b1a5bcb48ecc5849;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17d4ad0df2719410010945e0ec546f62607ab10e9de6882f3e470bf014cebbe4da61d6b3871116d9c7b7be06531ffb214dfcc15e9c0400d42dddb5f6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d896dda9d760db2005cb1fd98272aace71f81eabf22d3fb6a25deb373ad575978fb21daed0914c72e3f45489d274fb7647c785ea50b9c856e32bb958;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50a76e1a12541b6c159219c8402d4d856f7c9da78c23dea139879f0f4c6b2b81beea32a73c0250fe661aa6070466dc4f04c8c7723d7ea1b151d520bd0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5edee3471523f49237f34892faafc7b72dc37a35261760343de468eebb73602459c9986d2a6e46524f91b94c5dad1aecffaf819c8b307181be885052d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h175ebc55df000dac775ce8e62db7b634d09c09029f3c73a00497bbd05478f5da1d461c076ff1b51e7e4f3395b2884e52953fda5ccf6befbbdad421e3f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba1156b29b28c47fba6c3fb55e08855aad977aa9fe2dfbd5b00b7f805c0b7442ad4cc3de23d786d209733ef006b44a9709ed1dc775cb7725a816fb1e9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11265ec3d13e973548d4a133d36972a1ee7e53af18c99d6cf703fc72b63011b2fc61a3c7665100c94e6390ac97a5fb06009da2869e5220088483178fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0f2e1e04c91e873cd1ae2323dea2bec655e874f514c04a523de228afb152c79674a189bc9aafd2a6e118e8b1fa92d0d6254cca243567512cb6eef752;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe3d78f1844a91603cd2a8eaefc502176324f1b533d3e44d96f2971df617955d2e3e9c00a3dfeccded1157d9851f2723e7a23b6b71470fa5bd1387c04;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae8e902b9b5e2892b6587cf4561798f491bacd545cd42bb957838e89b44c1c8c9654c615c82f8cb3c7e61189b6d78436ba989f06136a17055605bb7e7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a378575a78c5c3a85ed443709dce2e227ac5c472ff3071f533ac1e2ba411cd8e3aeb5317e4f4c6145938c7d9a2125662ee8922aa87e720047c503770;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd054e9ff054dae5f9850d5f29b06c715fb205767f2cbdce004c05046224b1d14ff2f76ccb736a2111a3f743d9f216eab3d46e20d508cb07d248681106;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a7f34b1c7e1d0f2fe0386919f41199eb6841bffce1a53e25b3d50630596748a1bb8b1ead11568193d074606eef8656f335695cd1083997e3d80c4379;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16aade34a385b0732c1fc48189f6cc859f7ec4efd2e83002674d9ef5eea1b1d105add0b0afb4cc057bca33d70cf3bfdd230089345da9fd50e21ab7d89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ef651920a0ce0e055b41c9a128e56c13f8caf24c9e831849ae3cce8ce8b97e505af1bc1055f9593d20f52d1cc89d91b776f9688db9ec0132a80aac2c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9423eba03a7f536873431a16b353f1a7533fb1e2ee3a1f5e3c051c0e94d3fab3f8596975dc13116791508b8d148a82eb63f818e25bba2732b478ac0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b4d539330494a3ff6d4c9f0ecd09165fdeb6e7d0a95e2a280b550887528eb0b4dccbeba27e29231ce88fe10e20a13a7d6e1d9ba0ccac06253a359e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48e6f2cd3f6a54989aafd3ffcc1339295b2fa004bb3845918ddb0e5f66c6549b1c90fa9abfae7a802efcd7e5d9ccedd828fbf19769b5db98fc13a1f0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha35c6133890cac1fb2dddd8f542b1dc334ffc4aafb640f58566863c8f06bcc12ee2da15c295eee353d2a5db0a5b21d53bfa81e4c8208ad7aa9106461e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b5d0fce38fc7d446c042b3a6c95be4dd6e0629ac0abdd00a5f2813a83663cc3f6e943e9435b3da9204afb571ef6cf2f66d51ec99d8bbc7fcc0d9be93;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8265e122bdf9d22539f5d9bbfd8c398c57b4760e0b24f62d91e0b2514e4d96e90749177eca7b0de2bfbdc82946166c91e0326e69af0e37c3d9016cdf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30cf66b84b0dd5b8cc282bf66445c67f74a54f2616f024531d6e3ade220e3f4b9f4f621daad492708f052c3d4ac68b78473b7afe15c72db28ae3b2acd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18ca63492628634379e38469797be9171e7fac230788668e1ce1e6cec22f9ae30b38bde5bbee2fe75f6c3114e9bfb576a8e91ac52a6fefab1a809caee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h872f5f5a05330cebcf45f38b78e7c38a18c279c64a1535935532f9d1ebd2d5b7d5ecdd922b17538b2fffed03b89198c25f057ca8ab3da6a78efc50387;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa0029023a624f0572cc9e170dee5e1654f6d83c1410d5a1293adbf62054b383a58861af273f93b3eac566b17b03ea38a5d20fadba7365c962064d18;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a74776ae88a56ff5191cf547b3bd909af6c56da07f291068096b843778cd96eaf057895993f3b782b63784aa2d949e4762d6231357eb2a98e53783ca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h764160e24ef8259fddfb8dd7314d44e9f616cd2bfd38af65ddc22d0fd22ba2167d78cd0309406e7bad85f0f78a6630f671e2d1e19c60ad50547b73ab0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha91600a50e9d8c7b47f4657c7477df6846aec295246b570c979f5a4123f5fe2f23b77cba68905755d54ef43c66a7aef8a55504d95046d1a54ca95bea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2770609bc7a80bdcfc203ffa0a5c2702d5cc2bc953f12500d4e74073b494e8a4a18d3979b5e2a04da89870556d0ba8cdc1aeec60309882f04c0bc83b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdcd1512f9b62d5d845de440910854b5fc7585e8ffb5512c28553e1ffe4ae92b2a4a3c1ed8b83a920fded0a90d102fc65c46969d65a91480e2b1f6eb78;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5583e246d757dc58f1c83ba2d5bff8e23560405c2c5bb9f46b415a9dfd364be911e2a94474e0715e406f021425d82652aaecd80bce532ddd36895348;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd011665390b96cfa298e501462748472a10d5049e53c71ef339645964cd0435e45fbc98ae87a07d6f6b29f706bb34c3be8c58abe8b9396e44854e7b6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a23beb40e1a18f6356d175d847edae53c781dad00069e71d933168dddac1593a50609a0929daac4b0d82338dd719106272214411d7cdbb7407002b1f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f293632ab2a4924fdd8e2016c33ae7227794bacb9302f64e963dc4d25244c09be296af05dff92792f061ade11ec7d43c4229a53fc900e83a2576133c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7585520bfbf8490eaf0751ebd6f8d8da898a05a8c1d54cb9d509a7ba967fe2471704a9637d4c154dc66af85d3f5a1e9b44c81dde988e0ff17e609a90;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fb456b75d57578419d6a5540a28809e75ca72d6b5a8a17908bb4c70547d9f9b09f44e900542a5fc91da0160f6b57e10f514d84f21f2cf71b02f1d23b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fbaad0934d270c87dfde5150161e63a80c62148cdf196314b3fb2c9dd293e05f2dce7775dbf6aee8352a4c19a783a7fd7e8658aad0fbd91caccf0e72;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1fea1f06101953516a97bfbf769a8d3129f52cc81e9555608ae9e8ea9923533ed51c95a16147ce55f55bd77b8d7f9fa48620f2621892c7ae0708f30;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b59e37e7d8c570fe66c4e39f6cfe28c4d4219e5517176f60f496a2ed3a7993e546021db05852e3006bb9d790e3691933e6e905f9be26d3305bee2b8a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd287997975f8e0c678ec2b02cff7ff97c1c4e5805343556727bd319b4f2f1d3d5bb83ca3a0ee6d22b81a42398ae015bc61462799d6effeeb6bba3172b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9c360f9b64284884ca2f6a532e7ea1a0cd8d5348b8aa70c939451ab7390a2ea90ee44e1d87c592e0b073ebc2217c1867510d8230534a02ccc3e95c3b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92beff52de52cba6825ed737a58f59dc1c45f685199af3243e24448c41f7375e16e7a3beb0ab90e9c505979814038f71e39b8b3fcd140b8ff763949e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa4da211329517d6c68e5662ab156661767435dc0e6123df279f914d2dd480da8bfe6ba36314a8fac44a466c55af1be9602c02d37df62cd266237d2c7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb9f631900ad1bbd14c9a3eb6e31872a765c1b33fa143c35de1fd147bb35834407b973ed503b32efd15793c5ba60e8b4ea1110d1ce0a84df3a1ba6ab6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab56ae52f42bdbe86074017ae4852a2ea62783905e85c2d06145b9c643c81bf33afa8807fe8ab8c852e0a6cace4c340b1deb88df6048490b7792958a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h760aacbd6611a10964335fb2729d124baba43c362fcdc8b7a2bb8e2e91019b54f27075cc0c571988d2a21648342fff3e88bf725175093f13e06846aa4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf086af125a36f6555c982b459e99909373022e3ad5d6aea3857186defd6bc184438a190b0f2df9b6b15884bafa6b866f677a93de82abe047bb419e97a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ef0f3dfe8c53a9ef26a13e1cd995683e2f5213e7f16fcbd10c5597a4db2a102f3b73f9314daab3dff73401fee50a05859b98ff0962e49abf37432005;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b599afe8b4fcc1193434c0c40f187e04a70d21a9aa2b57240d3adf557e748a03626c13e1779e8d5eaff0c9155d303cfdee6f6a557618abc9518a0d21;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb18df8d7966af1b9e8b9d40a413a6cfa2ee9a9eebaaab0870dd4d176fffd29b42396f5df776d6bc777ed0e92f091fee5c69658bb837ab6f33e229a2a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a4d13e3a9adc84b9962d67f5f7109bb8e6b59451ef4b61805a03dbb6111e762dbcb78256c7392e6ae5fab987aa9ab388e61e382efd8ee80a290c0ed1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h233ee764eda6bf3ff451ce984fd6284ab0eac641f8f173cc298438736288fb8793222c25e22b63cac45348a172fea23e3bc07b2800abbbcbb72e33b4b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ae84b9454d2a808d4b1d6d54eed841104672b2ad4784530b0b9b516ccdbea477246a5a15ca50f3b9bdbf8c0eb665e518b57663ebcd54b0a5beeb8fc9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h389967b95935064b96e88cc8d7425735dfc19c41b97e819b4f75ebb4c5f52abbe67f28758125c4dfbb7c552f4ca31d80ea6c6429560a08fff86f154bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8485a7b602de1d1434d7441078cde2f8e600c407cd7d46c0392da8c6bd8ee4313614c07d00847222bb8e21bb7e4d12eab0d9eb03b8491639c93ed4ec9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heda592264ca765435f47b9a10870045c980a4d3bbae8954d9dd281a3b7df61a457e429f8fa594d70d930082a6d397ecddfd84cae009e56b419f64efa5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69f5803c3ea2dff094011a88c4df937e89ff0527865fd13a9dfd6bad656b775aee1a16568716c64f4df7ca82daf343d846d61a53e6a3f536d9b69ad6c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h829dbeaa1d62ad34002a87a06337d649649d5d27b8843f8ff17635d2d8323f01f23edde0bfb825ed8289f918501b69c4dd65b9f907c006a4bd737ed3a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0449682aa6bae3f40738b89f778629e75fac8d31b4fcb47843f08e23a6f49440228c0505038161b5580f69f7fef6c860ef3814bef60c4333ca7753ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30464d4823679acc10b65a547f0d2a2d6343cf4272095bfb7eb2d8df9841b52577c01ffd0ae58b6ee854ac768985131986741451964e7afd6d2f0091c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8299699d1296965f6a66c47d252ac2acfbe90474e073268f67603a0de8642a8b7b00def4feb8eb83738222d81d1731590939ea7c7400564b53429e6c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ed0582e7299cef6902b741e31ea385371d05a82aa07f6961f1e09173edde80dd4d50ab6aecfb7d85cc1a2bb85e75b0b1c0541f2f4906baec67c1c5a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98bf2253f4570125ad2cb2a29f1fdf5648b23ab032850e7f129985cb1f5953b7f1a7418ab6d63be1257d0be5c3a15ec3d6a9836307748c293dbe38158;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81f38633f391664572d5d7f7238da8fd52a842d2834bf304464d3b1373648f57e0320dd2190c4973d613e8da4434c18aed987c3ca3a1291d804302fcd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ac759ad78bfaa1c88ce188d1d0e0715b8bb3d83f3d13ec45f3b040795c3ef41789775c133f5ad122f81c2aad63329fff4c0cc3f355ae2d199c3f6d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2d29ef68200ddc521088ccc3c881d0c06f6cf3ad6ef82695b6c56bb8dd19b8b0e51d3e1b5e1556cf65f2cad92d5f30cfe27919f52accbe27a7c5de19;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a0d0f4b82676f86386dae4611209c3279a99e33f1564ab73335953f92118fa9863e9d214ba5e647bda24bd97feb02f4f60d72e0314d419e74bd9758f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88f55a12ca6ffc40902c7576968f5aa169336492fb8ed5b9a435da222e7581df270280ba67659f62aff32e5f896730172fd435dceed12e00c7aec94e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h391f268eab6dbda4dea599420854ac3a346fb0ea14a38520a715ac3f765c86300f5e56488930d887682bfbea0fe19d6ebbf604dbcdbe1fc53efb292f0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb08af814a9b5f356f45a4b666f048837a3998c4663c775b098dc61e942dd59aba2f44ea041d6eabb6476ae0c033b262101e0087336d0691e619113178;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69e89efd8d1b25674dbc93680143ac5c30079673c9c7b9775f3016d1a24aa1e17e688d9303c1ce93e598f4242b26280507c60d10ed8889cb2922408aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4ac089293df32ccbf64da45187708bfd0cbcc8272e7bebe956ad5a07e7d6bce54098c1f8a6168a61550615cf6ca807eb7ac6087853ce98ab61cb9d99;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f83a141e47ca2e8a5c1a6976b654a3a7f1d7e4233139ed80fdf19372fff13346410a5986198993687817871675c5d6a358adeb00747f67090ac6dcd0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a6c0ae6ca8971a403e2a9c38c238997fedbce7a8b082e78e3bcef1f9e531946bafac19c354b0d20be79619061be3f7af174f7a2083ee89a56f4e254;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h435991a07b63797a910645cbe803dd1eeb750963cea605eb1c038500718058402be6ac97b889c08049de0e405ee4aee373f5c4b3c8147fb7018efe6e5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hddab7376990e794bdd37d6c3527e966548a71f8e1a0a29a73d4ece1715915dc803ad4f9f967eb69b876aab9a5cec9da996982e363a83893fe4b23c045;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6feaa9b7e62bca3967e651f5dbfc26e681481d6c205c0abb6740542ca808294cfcafad38ec4ec030f76c0ae5416ac77093a0173b7f753f5e54e49db;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f9f740a9ef42d14f4d5dfec6b462292fe75b8fca6b449c0bc7a2c669408f1c84103a4e43d8c8297d73ce177b9fd74647d82d12409d759ebcb6bbc68a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc43dd3951fed66875ce391549fc7e7a9344815730bc84fb7d60e60ab7c981d77b3b265faa7092054ab8d5b8b974b1945e4c56f7bf0267a048c6e59652;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33124a57211396aeb4c08241a3074a361330008e44897f57466d2d99315a23016992137caf87a082987303ace20d86893506f5ee565679205fab5b9e5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73b2665377c17f9e93d30a136232a9b2315debeb9ec327c8bab3df759a68e59b8f88bad6d466b3e424fe1e7781ba665f8d012c514bd6398606c738353;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66b0edd37dded17b18405642b1d5383b2cbf325c5f58a0d4b011b7d66d5a0f6d485b8e902bd98bd1efd2d55fec26e2c00c811df63a0cd2d5b0adb3259;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8cb74fc82443f0b881d46dee7ee0fb3a7c018ec713be3a836c4fc634d7e839d864b853f7f73daaf6a6799ea58932789c96d2de9e373feaea686ac7553;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13e66a10bde41a9ca03637184745bf76ec4103b2dc91a16f43e66f177ab9567d88beecc6fe72a6cc560144e4dd57f681f208612f8c82f3ce539ddf568;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd54d3164405a63a34760d5451317e7f7635b86a6317a8331bd4b8ef832ea5e24df04cead16e92c4b93a569d7113722c670dff4049ae91ca086d13c09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d59455d042f766bc327c87bd1a1ee8354365b9b156fee906fce8ce41b49770541eddb60bb3ffc4fcde6c95e623d8e217a950b9abdea484781bde7994;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h948cf7fc02abf6d1aa3f679671133dbae8a79b5a3a0260aa32e79af527dadbc0f772f2251545bdad2500195a74b07139cd9c7383268fe7dac0a3cde13;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e31361d920e7bb823b1d075212fa06c48e8ca36d53f2c9c25bb21eed91ddc1844e9cbeed65a85fe546d7eb1a3ec222ac52d6d913546828ee279d8faf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d7064e4dda1f058838b7e7300a9e14954023ad8106f5febb2754a7df5e81e8c91063b7eaa0cf0373c5c0a99a062230c9d5f5aa719b2a8b34cf4c0225;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bfa5b494a77f7ec7d9c09d8db62183f66a3bdf5b651e9aed3fe11f391fb474b463e1d6b7577a4a445311ae9c8c34811bb1f7c8c738c800c8907d4b4d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4f11c00bfd63e4b23a9cc58f6fdd51b5fedd48ee351f85cf9867128371fe34bc4f0f52f48d128482a178193e914228eb6b9e735801f828574f691b72;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8938ec35d16f4cafaa59a367c157b6d67c94d782b5864402f1603716559b7823d4083705d973ce2df63c11bba817efb6077c4b5004e095b2c9e8dcdcc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6053a88c52a6d0d5ac7131597766fecbb01f5af1bb9f37029b80058c82003f3265be1458555676242825ac92c61e3ba5cd2aa80f3de0ca5820d095875;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he347972a61fc49424c04b40719eec9086590b2c6cc7ca142c8aba5a7f0f32335ca93eebc567b15ce53dc42ca69866dca3735336b5e8d3380a33a50ba0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5453622bdfae83b9ff00fc56cc6e2d5f285b611d80404e667bd7b9f452c0ab0ca924c19434c1f148bf98066ed76813bca78851fa400521814e35bed29;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h512b5a8245a522bf7998c5d07062f4d88e8f3646d5576dfff579773cff3aebb98fb0313648e54c6a5494c93915dda41edb47dcbd49ffbdc585a5fc9a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac0aae63d8865e0824434877eda638d27f965b65c47b449cf650a20a848e61a2a42b8c65c84b2abc3ad909629c1f4516abb9f6a44eb7b111755413b7a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3d564d002f00060574605963b06b3c75dd7812ff0e90c92f9abdb160bdd34cd7701ad144c49a79fde83ea8a9bf307f5c3bff8b59788951aed540f8ca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he17523ca38ef67458c607a6d8ee3517c8f977e8c4a0539b25ddb682f52bfebf5047b5a99c0f02244f84242657c192e1c51ccf700544f7e7db5acf5f8a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf57f94a7c806c476d324176099e14f14b2e49138447d07030724187476fd0273dad34b8ebc6692c94b28d10e5ffe769ae2750049493cea562e3bc9dfe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce0fa0e55b45225fcfb3cb2f2347be289011fb13149c524b3e1676d740800135e9b9d47b2fcfa03b3e4ba17f5fd1672f201125dd9f9360c4316d006cf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h298794ff2e7c47af3fac1eed8e5e2a5b3f46963dfa07c03ad3eb9abc8812a312979c5ffe711787bd3fea51ef90689c513e603527e918b2b1a25624ea8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2405f397086554fffb0f16fa1c58172e20701c9f93bee728dcef265eb67ef6da2fa90ad95dbb23c9fdf814a955af6beaa48a327f24e83cd93ce5dadcc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e1e2b244a92f25e88fd7221da7f1c40445d5013d3bdb8bffdc925f2c7c2d42b67c5cb693612aafa6790b0945f5575269ea8e6dae973ac368ff422367;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6cb84261d71e33107a682bcdba336b83b0cc8e8a5ae26621d449f5962f4afc8883fd82278a64cfeba80470b59d6faa14e1e1a1f957a4da9ebe1de4cdb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he23d865be0755b19c5d4e983185f3c4da0047ac58d276d7d34d8e321ed0880738e34095f588eb3c439232134fbe4e4fac4f721c7b0ed5f6109a10ca52;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha416c5a697cd0ed1b793a81105756c24f0a8ba91a19353335b21ddd1566a8c68a2418d7e3e739cfc3bcf7ed073dfd237df2d2ad0268165d54b8d2d16d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef3bb1e6375678a52e05453f3a98f9ac66904c3d6de4d72ab1a7e5a0d96e620a903a4bf2858b8aebca42604f6dbd2859343b492a245cdfd0205cebf28;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc506ddaf485fd6df1409ab821bf6ed61dfca6650d9c58c55f8c232ae773cb5c70ea35d245006bf26e75d73e736b6fa7d08c970ab41d8ea082f9177b50;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4522f751475ad270a1bbcdc3cc89399d17db90180067d2d7ba0d8d68feb05a62a3a13609f528641a2d41cb17122b868a7c45dbee9e1dd6c9685aac07d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f2a292b65758a547d75a1ea3433024a08eed29111660171a31fc6ff2ec62bb8be2c84b7c5f45ce933d87b78e241108b5d960bb20048fd47a14736f20;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5e13c2f40b907a7faff4ba135aafe2eedd9e751f171ea5d4a87d7b516efc0e4eb622622ca34237af9bf5b6f5bd54df6cfce265ac8b1f2cb80658e01d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf19e488ae90193dc09fe67a0f62c422c298344260f4585d4e96c7e04b5e67f52edb89212476a8bf4d1c62d9756bdabe71b6789a8f77428acd86edf84;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14588948b41b0cc14ffc0ca7456fd1f2bf25f2cf0bd44d37adf54f943635aa62fb3f258ab7e5f50e79bc95b53b8882fbefbb553a755407ed0ab3120ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65956e0de0e0bafa214ab2603957d3d312ae2ca6a65d3bf6f09ab33452770b270845e83a49eb07a54761780a6d3010e8d654b3e462063b6de0c0b41cf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ddbe3e3f844e7c3c5b68284d158b66e54dff030ebf42a353555e0c88443a348ee7d98555351dada20119d8fc368d0e97d59e7ed37395603b7271afa9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7c0789d9cfa27f49352536c7b4871424e2daf0ae024fbe47f6a4880e166c37bb4e7128b68aa003762a65c602714f83d618e87fce1bfab8c4c2962765;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h806163a9f850c88bec3b6b4be754e5798a201c7cf0f140f79be4010152c1bc8a2105050d2033454a576eebd0f88aed00312c80df3cf9dba392f085a0f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h736de43773c603eaeae8ef2c7ff6a148dc55e4f62ee723a9a8224e04dc20723d1a3aee03f80f208ca6107bd3e02dd0ab479f6128c3d886cf0a1e20b4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc087acadc7bc7479c2ca08390c80e72067d71fdf662075df89d0fca9bdee6dc7832504a504997920c306d3d9ddc962a5bb38bcb6212a55c77310e9f39;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h967b65160dde63bbd09e03dee56992e41ea94bde0b6eafa67f98ad212af982b6116db5993c5836fd6277a198f4ffe20668400b0d42673d5ba6a3694ab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf33dc4afd9e996b6d48258a6d2614e1d38c594556694092be5a4e8c285ccda5f02ea6244fbed53f240c8d63fd02d0cb28677fd21434b98efed96c9f01;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1bc6fd00208b9f20c423701ece37ebcbfaa5b0cbedddfc4019780278541d1c204843c30e67d0396253bf5893e1a59d2ac561da0af328c3ed734e993cc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb9596fb7e662c94c40f9a8502a72fba935a84815df1556cae2af55b95c7c5878df9857e9fe13d10b326729e64c606fc94abe36ac64ee16898293fffb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h609a9b9cfb2aed2c05fbf4a21f1aa33e14b0fdd5196edc72a2fde2c74ac93124d98dbdd70068485c982b3fa475a7f7d1383902aa000a9e021cc5a388e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f690bacc41fbb7be28fda3fc319e488565ac1605ddc7cf6c453ff76d88759e03487d92144aa1afef4643df6008478dfd2f75aff8a27ef9f28b6ed447;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19e3c6d3dd91fcf69ee10e86848988f3729f1133650bbd36f109ad6d801c8fe1764a5932f55e417038cbb4fd12dae9df35bbe2b13785c20950abbb806;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab30c622aab96577da41eea976ab487787a29c66517582675443c33d445038cafc29064fc0ff588f249385fbfd74aed3c93dd6a1fc0252d668f69458;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70a8539ecc99dc25add8c5dda1c5861617204d70600841c45ba062530e73e2468fc2aaf02aa1f271cd394fe686075bbb5f02d096c516a71d3f985fad5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2caba0b95f93f4b40eb128d1066b1717ea66cae19a991495311498dd871aa03aad23d212bc1ca1c43a16c1d04800f6cf848c5983e30e34eeb8fa50f4a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50e33658999dd7848e12a4e0222f574d4feb08e7541d2a8cf1988640c0c70d20315e51394c646811d805e1126b43451cddc7d145f25f774902d0870ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he300577db03f8c937cc67c6b7e5c72b87d1ef8728b5fe4a1d109537cf4438cab4330e94db273104cc19c5cb8b911d539b3956b9a3549e83f7dd0cc34f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10eb353328855ca9dbe9f76a355d0c28cfa67627144d447040ec3a80d698f9ebef09f43f1501031353d493776cfdcf5867fb94cf7fe1dc55f73f6e76f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h770c708bddae58dd8c20b175de902b23801f955073f45b47b0493bd216a1ea85a54ca17a9a9e2a2e65d1b5fc77d89c48adab5c1b57739146e59d5ebb2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb16fc5b7c3d00621b903267d4dc859e4fbf111d62df7cf5b44e81baa1d87b7d71a8d67a3b0162a20dc3df54411c9cf9c1823391f282373d6340274a7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3cbf9a54b31b9177c8623d3e63803352fb7f59362343634f4fa1a2306cd46c67f81467a58e1ec921d50778220d583b7c3e4eb787e7589de2121cc0b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h243fe714aa04cb235a78f1a35befe10d97e6c59ccdf1c378173037741187ddff0ed464442b5feaa5ddd8e2d9ffe119c15e9b87bc851c9fb366352ef8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d67334feeabd4bd545b3035507f6d2ec74c573a923b957e55a568fdfef417201d99a9c12e40edf9fab874083f7e5b3c3044f3d363e6e73a615eadb45;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66fff7f199f07fa816a234c06488dd1c2e09e68f19567835a630036441648bf5ad43dd6debab86fd5eef9ec5bc6b1337d48bd97bb39d7332607c551d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4f723a461d267efb7799f07574c1bfa473617ff9da4dd4468ecbc58482cf9f6d3ba1fcdd44ea3bdc1a05198d284036503b4fe4a1cdbec0a6229ba871;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc56104fa6697571ffdf050362a7a57bc887ddda961ad8c254e668d520c78c9165810ed632f8b321045c8016a0b85a652b4820b7de1e54bff3c1f83abb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3bd21dc1812b908c73960022e1de27be90e6cba5dfa1ee4fc26a67140a245028f7ba2f90ea9b3e0e1681db48dafc1670c5e7e7841161876c64085f42;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25eb23573c931c467c3d60fdbf497268545da385d6ed652fb49eddbf329106b804bbba73a1ed80d6512a3d283c47d4598e4ecc3ad9f1d4aaeec5506de;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda87f5803b3c0b86856727f249022c623f2bcbadd0d6c4fb5ce9b8384f72171e7d966275501f69962652098d57f45cd61cdd00a8ddab92e77aacc667;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47dc49d58119d09a3445ce654af5affc9009d85252066fed1b3a69b991582b9dbbb0f06f53f1b083be3007a4fa4f0cb10ae1a82264c4cc53f34850783;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6a53596ebc3178e390ffaf21105927bdbc31866224a2300e4e0e898efc32ca16111f9c5fe66b92632585d1c5989fe819044bb55072e6e189b205e7d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf25cdfb83062f4843ed946972bc1f1a322112fef6d53acd09fb54b56afc68adad5fa90eadd99393bdc9a6f20f347c127220f72e02c52b6cbebfebbb9c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90db47fafeb3cc47bc3d36b1a110ccf859d35c8bc1a9a0bb0746142ed13d7074e6f543ea2882d3ed857715420db3f8520f25b4f803b5ba9ec7342bda9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51f98bcdf7a63811287003cc84420135f5b889a8df0a9970ba71d5711568b2298ae4a5bd244f027c1f19c2841a063dea7f5e20e4bed664700e231f90f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce4eadb16d323241bcccbadc32762b51e002ab265e45b5876a1b8c37fec2766a4182157a6ab1b598ccd2c936ba7846dd66d31613f248c4bf2d9f852;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8eeedd592b92fb353ff8edbb561826d5b12e0cd352ad53a68dfeb65cfc5813b3731ef26bf61d794557e317d33ce4c0c1e6d068fc1929e302086eb115;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he24c312b4100a188a33c278dfad1bc3c1d7ee7614f041c3230d72f9539b7b010fe161b65c52d32ec37650fbff6e1bd8f56b9bd9dfc7c9a1e2c748070c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdbd6a24196c4198d5a4fd69db2786db54fe59639e30e54c69a7b16063d42aeb9f633072c7e9ad641d79fab2d9060733f96e10aa82240aba64545a815;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdfdfa0c1b25ec0cd412f2687ca6fe1e5103218e16953ce92aac0fbff6b8bfea5de2dbd1d7cdc39acd9148ad874402b3cb741ee6cf0e9de173e586feee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h717767303f4eebc2c31ab4376f8cf30f070dc26c5f5990b23656ee0e3a75521d62cf50d2a241fa747ed73c4025bb7af96c72eb5f382473fbd8efd59c2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2a85f875e1cc52e5c5adc867ec94c1589cea815b7acb75dc049a93cc2cad1c4c64d93d9d546b3c303f1da05d23012e0679d15a99a47183d963656565;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h277e136b3322f3dfb372b2afc7e7fffa7ee06a4bfc7717bfcc7cba1905a3ce9f9ff5f288e56279761a4fedf8f3b60f46055a909a732dd71767371bf53;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7e17ba29ee4bf74aa7717e2c770d124a92a542a8d0def277291881044eb755175c2bcc9c6536941f30f52e89e52d2c20dd7cabc98d3f2e52387cc828;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59455378ac1ad8f597e48d96bba85c6579bfe39b89a227ddb88ab14b66cdd7e95b7224443e76d4ba48c840bb11f4e25a7c6bcfd2214fd5d1406b991d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14be1abaa9841b36ab2fbfa82682f7ad010571b759c49af01b3c54d8916c546b27d9c710a0ebc3f9babc095586c97e262f4967328072d1163752e3fd0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd01b83b2c7f2f9608d59144287dd38abbb19bdec29378665d699a4adfdde88196df487b6a992eb54a32d2f9fe87c4d879bd6f6d5eff0b2fd063e64485;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1b91ffa72804644816915a96e7e0e3f9624c5e28194dc7f05958f3c179fd45b6dd24a3953cd42c2b3646d582cae7848ffefc38a701d8fb2a8a626d7b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7de3a29bc449f4d2ebb98edd66ffaee7f0b88e58a34898c2427e9dfa9f3b373496e7ded266a1ffba60ed4477bbfc4d01ba2bd670a3ee9f4cdc3555198;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64caa22fa86fcc5e5b0b35760efd8ceff81d8ab7559e9d63d14eaaf8736a3fe7b551bf74028542879dbc8e7ff1d4902a99b1a280840079ff4e8dfc6d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab7cb693d996aadbe2fe2ffee86764094c2602490b0ba786b6958b6724ca6ab9c04e23d574fd1054d5e3ac8b150026b08b59c0566bd3a1493dd7bc238;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7ac67b5da64778022eb6dd8efff0830cfcd4b906c884a966a63c8b5651951135fcfa252fb58b101165def81879d52925d0d9cd4d6493b5c49083a8b6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ce78da163f110fe31afd6b27db7afe3f0849874b9e883d991f0585ff13ef020f190f890a258116c230a849d1cb9f9605b2240383b49e0fd99f12f61f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef9a4f24c38ff6bcff295b68821ebdb55d0f123306cdd5861507671eda3d56bead31504536b47ccd2ce8c27b0a907a59397c4058ee830937b2692458;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fa3d84057f6176bf29c437c7f71f20395ef1d13051ed951ec6ebc10c14b0193dc40228a6e3c750ae55b56870a476b0cea20ee3b8cc3a0a68cd7c56c6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf252ebebd25e56b7cfa9fd47446808c6e88183cafc6eb3cc974df52dfb88cbaa6d2d071b7d9774a770c4a89684e3b1c210f24991764fa9c816b726717;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe355a273fd1bd2945a4e77243492570d2ea5b59e312d8dab6456d1ec310ffa2517a1a235441bc0c2d92063143e2d52d05ffff925ad6d8fc78b41ae46;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcc0cbdaad0b6a3774d4a49f9db49d4e015bd7e1b1c377b83cfa55570a1c6cd1e971c7f7472d3d63a18bcfbc345a746fc2730f56abcdd9ce8ff3bc163;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2f9707759bfe475dd532a3fd989b6998a635c980d1b20420cf915aa64cb8dc6448880ec547bfe9c54f9b5edf01f90ea517f1ffc10a9f340afdb93903;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4638b7b673c7057414e210699c51b3491f82cc01bce93593c91c43f8bedb73a810d2b66a74323c6cca23a564ae3b5f7864d90224c8a34e28cd21926f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b52cb72ab72c90b856cd615af3a047d26b5c0ee991255d5612395c78ecf0bb7b44225d84cd6a3f34a6be494fbecf2ec61eaad5ffb75024a0c6e5b072;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7051eed22cde3cdf8829e852462141eafa2670b9e16e4dbc7c4e7d3a969612816a5ed1fe30c4e4787791e372ca73a07bf772778b1bc400477572c8d3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebc1c2cb51a7de16e470ad672faf15c302802359d9c1a2bf130cc849eb85f104cb52baa40d2037b169a9606c693359813f7958d04972eea4c67bdc57f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h101088807a67b0596bad20871c5a225a635f43fdc6b4463a096d4f85424806917c13e0a66ae536f68d13803226fa46183a9b81acd6324ce0e56a3f09c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f00b37b3e7a52bae837d7b26fc728c223963ab3c3ddf3e9de6f21f7c332f817876c0b9f7ead8abe13c0c0572d624baf877ba7ba1aa7099096826a777;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95e7a6ada204c70da03dbcd0d8682130cac50ecca671d6c8236f2a56d925acec4c14cfb9131e9aa5a0d1a274d9643ea05609263a9c84357d353493992;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7fb36cd847e1b48f81bd4fd9985d92198b485806441e4e6e3e948d096ce77f4c56474a2ee6cc9a42781012ffeb1368dcf74436fbd12e9a172029ea024;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c8c628ce846a1bf5ea69f7f465f6afa806b48967244fbc040d24c409cf7a9180501efc38f4e10b7a536ae95b90ad8e4f6110afad9457e1a4ad3cea95;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c966150ebd87c36b270a3a68da42c4594f67a1e35798d9592292bd0b800bb11e38d495256ef07792b2715ffe37ad595dd976d1d9c639f07bd8086b51;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65c59102d1d22190726a06ef30ba24216f8d64c8b2cb4dab8111f05aee82b89bca4eb105252b901c1f71d960d03da834ccc80642b96d6152e8972dc78;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6156366df027c86a3218fb770a0919966e2931c3b3822790a74968350de6c4fe6a8b83bd983e96098af92391c6f70ce8afc3407b52c1380202a20abe7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc10d705a8cb776692f4f5adf773476bf24b3b223d4d99f602d410bfd3f8bf5651a9efd442858de37ebd7fabcd4951f53f9c43d5d8e8c00dc288d85820;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc7545a6f790396816621eea5f15f4449ae133c3046b12c20bc6dee5025eb21a5dc282e54d03d981fac38b4028799a32a0442bd0d3ec4864c5188ff93;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5d188e5e849b7350c3f4ffe6089aa3717f2585817ecf0d61729b8382ee622661579ce55a4ac0bfd921b46d1c9b786af8440ac11ab957cfe992adc11e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6c686756f93f4ca28259d5aa602bbd56d1012448217f6d14ee8243ef23d056ecbdb3c7ff18d1a95dbcabea528557407ff0de45e2fe10914acbe8d6b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3c233b295f696c22ffb41ab8ca2ac12a526189a178af244996d53cc7ee38ccb2d9e2d71e6c30eea4f5364f6935ff95181d75186e1c7813a1d9be8f81;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h232957e2659ce2b1da810fe0405cef931f4404e077b82459186a741fa1835ff8a2cca9d8de03594ea1f891a06152b30db4640bed0cfc730a26a7e8aa1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5996ac98b12645a8d2b9defb61d0a227d31e5b624c317f8b0540688b8aad51664d2984439c92ec2d16a4d23e46c2c1f129b8bf4a23778a29f04909137;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc084dee8d78c923e4b2c457cd3bc78da5acb4b843cd3a75b96d9295b8f0daa5ce52fab11027bd3a9b0de676fac17846f90149205868c68b1139ac95e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8d9b1b0d503f8c538a4aaadfccbb6e94bee9b331070ebf8a8a5173477fe6921f0d53fc0f84989fd42be987e0a09cf2224688a5e9868dd6c6e4b10f75;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0f4f2dac77957b612392a05a582c08baaf02206527bd5f2c501347b523eb9d1fda17ace678c866ff861ec95efe0cef8da1603b8156e03dada209e5d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86261949cc1c99bb5dc8bd4338d674e88e6d774bafe23b4e3d3b7638d48c84e3a022d9f4de921f41bb1cd17e160f4a951a4bf985d42653f0e8f82751;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h379a6e047ef34435cdd059628e36d5a33b4ed6aef7b16a8277241c0f892de4522797ade01746c7421155424f2c9507b295f89c4684482429bc776432e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf79d8fdf388ec42421945baedd694eae46c3e54507b8f7e013628e849b5d65ba0e85aa3ca0dd6b9dcc428843c134e45bf52c3a881744b8d37dce3d31;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6cd74cc761a29bd7e0f5d3b5264125d32a77560eb7fd0771a99ec3ce6ad262ff933e96bf9a05a4feb28189878dcf17dc9e2c374a38bdbdd39cec1b7ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33eadc9ee7fac545965fe6b9c914b8a5b59dbaa17ff4d12fb40f4d5e63276deb6aeecfb98b8fa89d3e2641eda80e18950def475214a30ecd0f0a5edf6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79f315af8e6083bcf03aab26e2b984dce8a8c8e34c0a1cf70e65307fcf32048a999425ceda2fe79fa7996736ff094518e618fe1a73879613c13784efa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3075973737bd68d7975b751bc169ddaf605b43e271e42354f12749cda7a51bce49ff79d7e027e908501d511682f27efe61e87fcc9ac61d81bf63dbcd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19e95a71ff5fec2bb86dfca08dbfc6864bed28501b6d074b23d60544dd616fae73babf52536a8a2fdd5ebb71e77bdf4893669c4a8887627838ae5fb21;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8db011aa25ea6c0a1216da8a77cca6835a87e060da4661498c076171ddf264e3b891c90acf5142fa5a52c6edd96fe02b33daaf342509c49137a53242c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5ee38e0d340626dffcdb7784cd85f4ca15da79ca740f632c839f47f4fdec9fc891f570b45ed2c99f68e6de86d414358e310b0d0c47ae2a9f693c8ba2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf88fff23e44e28e742d549db67258e94d9fe76da9efd063d3b2a0485eddbe730d25b859c4ed705594b66fc850e1a67b3c4c582784cc79b26954498231;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8b9f18a7278b285d86b0b482e0ab405e56f8c846feb2ff272760de3439d43cc5eef8ff4d33c5d6f3bda14344848167abbaa56030b096d2a869640643;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77af0a008709d176bedea40ca217e8d6e587f630cace7d4e34ab9fbd1f5c5ec9d1315ef1762c62ba54b7357debcdce30a6ad8efd0f4842a9f1576d149;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2f43758662c26e0101faec9a341ed45646f1bafe4135936d25940d62594ac8d9a0f22490b5a73273d3425347ce7b167d71181e41af593db246e3654c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc715ae4689e810101ed44633e4dce0ff9e5664fb4a088e07eefcb6b63a1bd3a6e25a761a04cad567fd2d93669024d02c4d93cadd51074313001d07cf2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd110e7579a5925a29a48bb2592f0616b4e9eedfba29c1248c763e15d04ae4b5a87002dc0163adc661051239d1fba83eac229c51a94263f481b14930b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heff2363ee9ded495de471343b9b0a5632db4eaee0925e56463b2e345a538223661668b396e2062a7f347d946800800e814864cca34375121e629a8d43;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1bda8fb9dc0c25449259e8edba55094b8ffc161e13c95979d7182979a17a13864d85f18d69792f8ab6850fe63d993dd8c4e967539daf5e11c1cdd6d12;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbeb11af4f9d4dd290799b810b679698ce610588fcac7f14cb1f9fd8848264c175be0864178fd4ecdfdca24b7899fad077f94b93e29b83dd980bc1dc65;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h256f38c3e793f322900edc475787321992c7acad1495bebd13eecbba90cd7b07ae0af294036a1cd727c7f6880725217c7a1e815d833d248540c882d5f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hafde2d46a292fb3f0bdb2ad5331b4109698d143fc354de14a91b3262c2a1ec6e04206c42f154ce4c9c7cb0309aafa3238ab0ca3909f6830d346392365;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a75cb57239f91c2b31d1cb1c239852e1d5c8c29ff2b60f331943ff2312da16daf823424f4da18179c8d71bc00ee62e0dfb781679c6ba776a5d3c5017;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ecacb17a68a4570698f2102e019443d132862f94dd03b33f7cab7753e363f1816527cf1e8eb6b9d0677bd2484bd27b319452ba3351a904f58c0426a5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51934c42a6f144b748643ec4210892ff8b3712c2bf8744eea15f2276dcc600d6a29ee6462849e2b848c7f5201062bcdb015da2754b163b95eec05421a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h149437fcf4122549268911d3f166fdde65b7c0e2a17ba11368ddf403211d27d60d6465b58c22205b74ef60a946b15273993f6ea70a588e2b2eea09ff3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41c2c2014dde800c8c94bb4a4fc710e84ecb528b16df503816dfa6a5a95a033f26c2add892922ef1e36d18ca55e78a64bf9e1d95792f29d02c908fd3c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7adb0e0e1d0eaacba997d8daf4ceb98b9af111bf4763745edd78065ee069d053d9f5144a00275cc6876de4ff114141d77d488f4d2826bc3ad0fd928d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5709ac8abbcccede737032577f2641d4d6c3df15e8a1e75efc479e5e4f30239871478931ed86d466b3a936c3ae5b83518d3a8fa2859198b11006012ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1806cefbc2e468b9a5f77131057a3c790121a1e26f8d1c0e3f0043528879d02384b31673e677b53c6bc11b71ff703979ca9e8857d5dbd4e0ee1b1ba0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bbd505bd3a7e8ab9f4d1b8a40967eeb1c468d69b22d400ab179cc1be34484ffbc939ca7d3f9611ab67d080a8b3f21e10e564193c8ade48688b598395;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0b86b2ab6519fa3d96dff32c6acda9ac2cb41897fcdbd04093dc9c4a390f520deca86b01a59fcd841c5e1cba574a6f3416c9a9fc125f5a95373e4891;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22c0a7ba2a06251c710da5202f7db6adb9dda9f67562ee3f6ec855e331ac9c16b0f8cc3bacc7c68adb5f2eb4d016f0a94127d29bf168b417071092b4e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb51f16736d75a00713e946553561d45f7b3a2365016917f2e27c43a43ed70ca9dd7cc15d50075b3c53b81066afa14948a7128a20af50e64bda3e3103;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee59a36f869201a04c6d759f7801b8a6ba9b8358779ff20f03b665ada7510e22af87137f4cfd30f0be27a958797b3a1659dc0368c03c95d9f4abcd252;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8be1f845e294f7c875f9eb886fb69276c19f6c256850689a25eb23e22780ce195614cd0c25bf71bb7b7204f50a38989e8007647406940af8e9ed62c6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33cda51ba7ab48347aff372e8dabc19c23f2ef833d001fc01d131a460fe846442105bf7a6bd2d66a92c3b893e70254106d20531c7e9aae9d5fbf3e5ad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hada847312dfd0357b2f2144af6ce63c97a77a257784129ddc23a75ca7045b343ddd90d7b731e1ae5f9050a31d89b3039e5e966a656ade0c7a957408a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d0e9eee8f2bada12789de4ed79f1c4cd01e2ff37fcde86796abf2792c8d6c7de91141f4b7b32edaad6b4a3460d1fe1990d7d07e726601e14d74476ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb7eddaec24149c3c287e37bfa2ec81fc3fd2d49734a5deabd8271a84975d22921304958f7b707f29555a2f15396a1e671d6f3acfa79f3429d85a529d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff5b5cb74256ede0b3eff9a8a50cd0e7f1270dae7570a782b9a4c03b96548130f28ee3347e902192824d7a420af839234cdc837abbf3ee8e135ff0539;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h565897acf501d95d6b6f18afbed23728c81a019bedfb86895bbafa52d71dcc0ff33c79b827bb88f9440becc3ebdddd78d0ec183d9f48b6907c452989e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ee122199fdee6a00bc59d08c9dadf73b5458ef46a12c9f24d1e8b2b74e95df48982509d003f02f42bbc4fb84dae2ef8058994ecca89d42e77bc25462;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha587a62f8da87595770d2bfee720fa1af9661d2be593288ab5750e0da92d644381d38a59dfb9b590e236a5e77b45a0f8bd431193adaeebfc1611901a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ff6a61091da71be67bd3ccbba4b86fe47e1c51c7c05b627cd411502b0c68456718700090a88ccf5ae1bc5370a66ee9434a91ac7b96dca6d1c5118806;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b1a5511a8d53760600eeddff945db639383acaca4f1072285825a67e70565ec50ac3c8952b272af655e3180b26094260a2dcea345416ca6ef5f6ca82;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha981c22eee1068a2997e3a23d2b366050a2bdf611694054ce0b6acd906de51003a4d7e2143b6f95e7e436d1498ac14d97277ec8a4292ef9818538f38a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc994dd9b5afee44a1aee1171b14aa482919a1ce124d028bb18178239418dc2dae32b0b908968a0a44362537ca16ac6b1cbf9537d1ef93f65d6a522ab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf18b99b4e6505d0ec29e201a6cfb3945fa0aa7cf103ddc6e42839425d16ce1b5c11e9a213e50acbc802c61f7904ea0e7acb0201c5b9af2f738bf74fb4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b7c4792a96e990f4ce4bbc1416728ccbf4c38e0ec810fa74aa58a3abf41a6744b779bd515e779c09a2aa100d8816da58e241dc07d627d9bd96bdf529;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3eba8fa89b197e4018757cb2e612965d81fb0a4241246159a64a33430092bfce7c82d8e95ff8a742fdd76c80586e485f371fe388d86b616a163b4f4ad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8941212948a9e90d990f003bb91e58892850b0fee9af2c562b7f2db9f7f16b81ef67f0e2376deff50b01145a50e02ee2603b1247a2b0ba6041c82645;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefd97819c2d6a013d88ca9211b8c72ce49a627872168a83db468b9fb5f711575f667f1b09905264ab9b4084607245918fd103dccd675cfc44f28519d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9ee4d2adf1d1e9622af949b59680136e4260d5cf383e92e61290a9e14952c3bd95d2b1b1904ec42e9761558171324acb2dc668bf60a2ac7cf1fa753a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea0e4fe5aad0b694fd2b896b6827d8a89795b272b9633056b77e4b11950dbba1cbd2700f5c56d10c1cb920c6dd24016b8718e9d7aad1f7ef329ca7bf7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc52f43960a3598099058b4d22d7e98f24eea4507dc9189e98b7b3ed5043a7f65c9268677e4b884a9edc471e0fb1b636f5822ef420cc96f4ff1b22655a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd777e4667a8cc9ca66f3072af65c06d47e5b79408cd0e2de7e936b908484db9efdb618bc4a9dba84e9189be4bbe6b7b0aefaf58028b454338bd85f833;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1cc3f0b57ec26b08f4075576b3e566c891cc905b7e537ecfb37f2b10f00147832d422bb3d30553e0295a6bd73d57bcee4fc02028bf50ea5363ce34d06;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2b178c0dac3a14a2589c478a4b5a078435c2d293422f729bd1055ce049a5e34bea6de2316370e270e3f307cd73cc11cd199f5e00bf4b035f66e58f11;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8957655c50ff2b2ef76baa091d4be68e144c5593ddd02b75e7fc00bd57bf2ed12a7107bb6ce2ff77b07b6dff4736d74b7e0e1fa49e250a0688619702f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdad926ffd6d1548b85ec1f5c994bc8c922764a828c43460194fd426d7ffc71ae76caf43f791c845ee2c503f946de59156c3080675272324b9b3ae2512;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7318376b94ae742c4aeb7ddbd45b30937600438184debb2f71eea3b3a73993be6b8872ac7cb2fc4269463397792b317713cf95452eb74f35825938613;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h637fc8ccbb2cdf97621c8ecfe2a8de6cb9d2f584c9f6ec0ba4e6dcfb8d8d6db928e8b50530ca8fa24224a6a962540d14cc3892f36c47bcd543c51287f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebe19c67e6984a295beb6e13f6422a2a14b4eb55815609d32c18dce2fa576e5a86f065252f61ac62479fb1f8d364f6ec75ef9f2e3a36daf453201b5c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb4605468a1e4edaef6041ea54ce23c7229161e207a7c04eafb2013e20cb40b393c70db1f57c9150c175ba9c5beda09751e11d2d7b56c097ea2e67f13;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9675b5fa5ff9975c03e67d8a884c4124ec5d93e6a3e2780316555614e9c71d5d61dcc0a8f4e91263fa152fc93bedc815097493b624a9833c7af1f0a77;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72b521ec40feb7e253e59de853761c579c5971ebca13af1bb424c1b9758248288763db6f482d6019c27718de5483fe35276d9cf4319afc679be177bd6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8de818904429800b629137974215cf6ef53c34f931b22107d6a8cd014079e601e9f76aa348e2e99dfebbeb63bece361b0035a2a33f46568c982e01906;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha89608f0dd8a6e9d8f285ff77997e63783c343b25f78bb250159cabd072d518957346ac05b11d6edf97c8e6e5d4d78de750b0420093e3612b7b678dd2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdfef3ae1a998699874fbad0d45b282fee0f650c68944f34f6c412841e2755853ac1f65290bec899916aad2ab6410721e549c90cd477982afb01762c69;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b29122a03b3c3fe4711a59a7df1e49cba671a5aca0c7258d5dc48b2855e466b1377c27b476743b07475aef1afd1be7d338c28b2f4489d3bd48d14472;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1a5e3f00d6a522159dbf18315ac200232efb4662856c4186a07124caf2d0a16b7c7f935ee7a151b97284f6ff154af682328ad6bc1ed13d217f414455;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5fd680725d89487dbe09149f41f18895b4c279e9f044a8a3d8c7c72881b49e5ea392e09dbe83b7b9800267f41b7b5e9f616c1e6279b974f9509c22d47;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd236e6e6567668444f9374ba0b460638c20da33349a6ad2d4060cb4b5f93c223d9a483b4b862514e30a0b0b4467ba83c95787915038d25eb54462281b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2b28d0e0a0a474a5b8ea5e745db4b7f68005642735273334042181b6dc8be790362310fcded158009f02a614a031cdeb54e1d175db942b85f7cba1d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9da5931ddb5974784eb0e61615b52e82797bf3c88ee5b0eaab6ce1191d4b61150ebdc82f761f816d5548abb9e4bbd1a512ee382744f3462bff68aeeb6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc76290b0b97fff0ae20f117cae3c9ca45ec5c5be45ae6e4b59b562e59f659bac6756d09bd36cdb9ec5fe4f2b7d73d4deb3d76f32022e55918a042ed8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f97803871d776cac69c20c7b2e0666c1d72623761b4cbda3df2aea93eea3b8af4ce050f96a61d11a8df598f74bb96ffac3c1c018a495b2d26a3abca3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf039a78d3da38a7543b4fb9b5dfd6553d9cfd9b60da5f9401c55f354eabd776ef7b8dda8fdb1de0e9cd935125dbbf52949f42d25c6c93320ec7c34b63;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21f5d85a577a2e99c52ed48c86c7d421c66038b2ca336baa18cb5441a3cde966ffc3a0e0383b029561cda51133c5eb5fdcd85a6d5b5dbd2f5265368bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7154d2acb7286c7b36e9262f2da6f9af5193d32c5a119e97b4c7fd20200ebf20171e32871013ce46eb528022f3ea34973c0bbdf8bb3d56e23edbd3a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h299e7f266eebc0854291e8daf19ab7d03511d85ad05bdaa21c3f7c768ad12223a20fe9fba867f18fb86b86a0a4a6243f8fd49562eea26b564e5160796;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcedb03508b673ac64d75577fbee7af875f22c909ab0cb649a52b18a7ec93db2613c64eebccdac1c3eddba535a2756da5649e553e1c599fea0734550a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a8dee038fcac60b560b720cc4ce21c10a22b0608c07922aa9fd24f4405a8d26f79efb9a93d83d3e5f036de63c887600e7f6e8ae63dd7f22146fd4b73;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd11fe2db86a41b62c03478e397672081d24f60936881182bea2a7d3cfc8780b5237c55b31202e0c18c86837c10c1aca69527316e0180c774b9a4679dd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae1af079dc3f560c52867e4de31a1ee83c09f604a4b38338ffecd0f297b25127061dd3ffbf194041215e1c89bf8bf81592b30d9064d968b8f418ead3e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82337bac1a7c77302a37b3684c0200749ab61567056ae1aa985be9a9f4e9c569cf35f8c6f1c3df18856e955f1a2822d894bf14316500094a50474cdb3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda9b02f38b1c9a24c616ee8a0c9acf15f3ee6909d66d565d08e084951722e280fa8962bdc9a01c5243183da2fe5210cf1a32132d3497d599762b4cee5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hddffdef5d9ee6bca2decef032e30efaed4234ce110cef52ba04fd71b68daa5736c78bf7f81d7e8e80a48668cc5b861af1bd4227ffd3291c82af2a7433;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he037011fcdac644d0692de57019b3ab97521d0fa1260d8ed1b59843d0009666accb3d9a48b9b56104fbb60e378f2c9bb5b628815240efb7bec0faa842;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d0b138003fad64416931b5de82d7df633836be0cb80a00cd07044ef7c8d0ea13422b9ab5f118cd458bf5647f5c321d3e3cd476530dfc1288d25f06c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc9153d56c0ff4df6892095e0cfe721f9c9230a023ff1623672c8fea0bd7d6214d05d2fdc4b157f440899c8bfcf44f232e582b05b062c28a01562602f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8b2795b677937669a5111b1e69826d4c7530f886a0beb4239b0a2be84c33f650305f7002ea39262de2151c973ebc34f93e897dfdfe800aa831301f60;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h556dc4554fc894a3fcb7dcb85706d2476c8322dddadb3e6d5bb5b239742d4d248bf7e327667e25b41137aec1278ffc01eb1d89257286bad74de38ea92;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b71ce87635116ed8cab39ed2a112e8c89dc9dbeceb084d692239519174eded101e6b084e5d0a01f5204d262689413a0788b88cbe5c004c6e2ba4d4d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6b2faa3f0966c21a5edb4db99cdfb4087e22bcd72a249192af251cf80ee5554f51c1df909e487591f07bd66355d4bfef6661e24685a3ce6a3a712504;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e6eac3d5791decb6a19da2b0a9574486583886f58dcc86d9987b807621c1ef0ede891caa44c38ba8e2055230b05bcfef18ff5c34bcac24ef61b9008c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb05cb56cb25ff9d1aed6ed1ce871d146586fa5385d5267499eb26a30e991a70bfa19acef24e093014c049f29879ffb70444d3e8d24205610e4e0805da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f849a74163adfd5c4ce3e3184ab7ecc93e84a4f6fd5eec5badc7e42910fc81abac56dcc57bd2a2e8372ef74bb10a631f36177049478e204bf03984b9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10140a6d2b3c2efd64f44e90640a548ca2276f1f01d1b541c7cb7088d885414fe1d57db9b07aa1e9bd1f2885f48e92bda6a4a00f3bf0f837a158f67b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2af47bd4300a181e7137bccb8884cf5bc06b6430538af9faac2b115517c04255b49314c36136fdcae0762cc7ad4621436b24bb6fcbe087a77be180a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha06caecb346e960f113c1009d9c396e782239d5ea530c16fd068524135b0b042bd5b7bad2343917be8a2fed010d3518c80706d4a7c9b120a2e6875e70;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a7aa1d8755d726242c32399af0b98b8c8eb21673b62247604228575386bc645909909645c3d941adedbca5b34ddb819bd93a172c8e679ac4088ebcc1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc1e686831a9a1ed2db5ab808719fd1155c2edcc71d112d2dfe394178f7cad52a388bcf6bd3dcf6c01355022a358eabb88dc317b3a9526627c11bc7d6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ad88d6d718db2655492a1684e948ccdd7aea9039127f2ad305bfd88a15ab090c7a8bf4dc79f9b159c7d0d2d08f7e81a2720e64fcecc1882845038b15;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he268f35006da91f6c85702906bc66595c29a8fea65cbbbd933129afb35537313efdccdd95a0c1da3f8986e52ffa2978186faa57da23cffe4ff7a8cb6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he47d160411696c6dc97913eb194896dc6353d74a6efa3ced93bde3d26b35f900e11665363d9a5b8ebfc0f05301e672c26567ad1f6ed79af630c44d6cb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa99fe7dd51936102b4516197824c140ef088b3044377bc8fc1a545c0d2cf9dd0cccb0b80d27b305b668769992c783571b94d651b9bfb5ca097d22858;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80484ed649bcd9608601f060cd548e73a26f0000efb35bdbc71337ec3a4ec3c8e9de071baadcfed1541c728607815f9bbb7012f14d61a24c7f3ca913c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d7de481d6512d5b8d31ecafd24e5da42fa7544e375aad89b796139212af6a87adc7503b6b5371fa6aec92853de7d29f8a79e0b275eab491d68c55143;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf3f6f9a6676403b3d4bf496ac92c9e8d045d4733cbafae9c2130aad6fcbfc5adc479dc4813e38ec6c582daff440938140d769dab43ca5e4fb4447302;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61f0bd8451b6bcaa04c26906d60d603a7f80332d1ca9b13a475678c36ef48f0fa6a061546aec5e1713ed58b06853c04aece1070a55f16b3d64c9369c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda1b2b83987cb6b7edb2196c397efec7c25f1376c726abced48054ea8cbd5ba5225b9fd7888a87adcf71d337edf9ffe4a42f96b54722f14a2f3f32ee6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74f900872c5abcf0728bfd67bb26ea6d388aad0ad220c9630b6b32a257bd7c455a8d38b8ae1a6aab998b77a55419c2f2c83b1bfe7b1d93e5dbd61b2fe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc660d671944bef3b56855bf65e354622110d054e1e003afb2f4cbf2c6dc391f3ccf160939618a01621a2be4517fddc4888294101c6effec791f88e8bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6850a5352fe09555cb8a988ff036ddd5f877df8832bebbca95ea36cb87e2f4c1aab98bdfe41501d88032982c1b273b11f4bd0446a8994d86ed9150fbd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4a718f7d1a6a21b0f407bff7ee1247fd4b73936673d444b1b33b99bd6694e8fb0803356b2f142eb228721dc6476cd3065b25c4a034ddb3c5795fca4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33dccfbd84bbf17239153fe8e6e6139126295d9165e5ea4db34687f4ce28f980349d1369485552f7fcfa742627c43712d6937975fa0dfda9ba140dda7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfbad325bf0b5cd54df23d45c0572eb2b3bee27693f52184a3b95d9e3c6280ed428b0b70a276af83901faa7552b3e71ebb5cd4ebc9a4f40c5bc57f8941;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ac28b670013f9ec9c666924d4acfa172e1aff6213911ac7283f1c090a8202e1fbc86ac7933c567015cbe05566078c2438939b343b52d96ba3c88e153;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92d356082d495cb3f361daf089f115873ffcfd303179af9710c3af8919a20ce5772133eb896e2c2f197eb1ae94de590fda66b9333655fd253fe80f63;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h966d4ddd062dedd3e12e13eb3fbd01a228aef0219ba94c99e683ff461b33d9d69f7597c4cce373238b6c6ccce8eea518557e2b7ad9e98060d7d2cccb6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8879fa11fa1a85fefecab8e8603485c231e0790c77eb767e972af34a8245a696051c85c9d654a7c22f2754e02109eaa51e517326609573874f6122bfd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b82c8d4144bab760640b6e3daf85fe111a21c9580c453317c9cf912d71dcef07adb7d0757045d4ae8e549de2de108985701d86c9b4e7ef30bd92c7fe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa55c9630ed2ba29a8a2eda143f76de488a87bf6646f764e4ca1a39629d1fe57709cfb9fcef91552e4f3b81c2425c7266d09e7766716b4fccdbe0aa94;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he36e2e19820eb20a3a5ac23acc60a37407b4ab50b0231c4556971f78ace65411b59f986d99c148bfe0a3dd2648bc6215be8660ba752131e70fa87a1fe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb7282276f031a720907b9520d0c35c31859623aec29c482075bdd720f1f517114d1cc75ae0e03997d18035adbc23bd2024995167db022c52d0d66c8f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a0fc798381fbb05a255155807bb34fecd1eada33700ac5b63d98471486dd55f5aa8b69c52ce2130e9e4dffe557cca9f0a6b165c6ddfe92399fd44fd5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9561410a08910a36fd04759e0cc73947d52971330a8601dac086294930726d3d2a2035b37e654919d9441d7ae0493f21b9fe8e29c1a3656afa6771956;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb68631fa50de23b9b2ca96feb1332b973466407c5e83de6e30850857285edb6f8de09a6bba71fe34c7289cce0c1ae39f90d4b31179f815fc9f638e54;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha43fbd370a96c70652a4959169ad9b39614b881980304f9ae510668022873efec2fb786dad21363905597d00dcdd3b89d748623535e50c3dfd8ec91cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa3cb981c995f3d7a532398ad7e1fad9aae87dc335830f55120cf7594e3bf188acc8ea24f01409c8af12fd6996f999340e813b0ae74ea5b0c0d33cef2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80be0660455576cd441df924d7807ccfcdbf7a191942cb677ab6dfb75d3ca84486fb5a45197eefed0aaf5300670675f73c35a0d4f597d66e67a0b959b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h916ef1b8accd4761944b8bd62d6485452e119370694b6690af045b8e351792ae4e7d1f537f376ca1953340cbe1686317f470aa1beaa5fb36eef77df8b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71e2fb3f9ce10408a4af7fd72265a4d026e26adf8c09fe0252e84a70b2110ea5e3a00ffa656f605f41bbdb1cd96d7a780d8e856a481614f98f1d63b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7accc6c487736f692f8db53110add6e060a4d948799ef2a609233d7c6f142d1fb639e4f63a2aa683479e9823050147d28c27cdbc4ac06f15e24b727ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b07800d6c1bb07f7db820e1900375be18e15fe22232fea601619fcf2da9f24ecab040ec684fd5569a4979ada1a99f6783988f23c58ed222ec8c54094;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3615328d5308386318ac705bcf4231d94d226b9181c5a9ce96a9416967f7e8ea4a0c03a2b64339b846eab0c99c33f79760c07f00e4d2e6ae15d17c29f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ac8c162e93e67528f61e5f6bb259b22ca57f83d6e2ff588b4aeb8e55b8bf752928f96ae721d25f499ab724a6351a2e40fe37ac59954656725ce37c75;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ada87332c8b424d469696d5898a237695cdf728c285a5b3bfdc1856d939597f6c0294984280cc48b693d5adcfc5bcac12525da3ffc012b2bdd98b4d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1da2c4d575d062f0a03e9449e92296eb1cf3c1830d860070efa19745ec0d8254c9aad83f7c7dc4244bdbf594df4b463fd913a75f51d906eb00c3d88d1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2dc78f7c78d19aceee3f19d1196d925656d250de19188ae3fafd11cc8e54a2c8df6c90bc549fe6afc369b86142ecba0ef67c5f4bbea917c3a4d91f616;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc57183962b864f8b12f43f41a5bdb8c413b8ce91841577d0d11aad16427a65db5b5e2ccc7ba1f4caf2b493231236b4da09d23a3c0d5e0f188dfbf1d41;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22d15fa545c94756729b595ca27bf543330486d8285b685974693246aeb26a0dd7e20a35a1874ecd1e16bd739e4d7cef5dd01e6a65f0bac540303b97d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd75e96d0d00f512d10e4b0caa26c7717a5f33c14e289254c615d9625a55fc9efc92fb67eab585d8a9fac7a51828bc6470de061b35cba74c096b1cad7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f481203c08dcc260c05301ff85a4fdd0a3cb32fdb2d25dc8f670826b3f02d92cfee3d008340b04d1b8c8c14fc90a08a9813999562e15a7640cf4a0e5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7a6d487f1a5c0f88615058d896e7d079491de929f6c0272f5e27589dc138c6b9255790dbb4d3abb601355aa0373474530ebe09ce324b05349a0688c9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc94eaa5114fe9a6ccf42459745c768b39fcb06998a873fd7b740ad8bb28dd74bed563dca6992fad3f38d43e9dd736232b10e415f15f66c9cf9d99472c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95143c1e2e6d562c80128def78b555b3d8c536e2d700f2a6adbfe4954f0644cc1a6d33f811c183be0d33b4f0c352b763c25f67a549a2e496b658ff660;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30dc538aa2ee4e5d14705d7f9c74d4ba82e71b08f288deb908090e4fcfb6c1b63a8beab42ad5fa2466a2f23e7356e1cd5125dee06e8623ee955686559;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha81dab8a771e08b666cb944efeec98984d9431b71526ad06963038e19f3749e7e93b747849fc19b9b89f52da9ee805ffe7a1e70daf56021188f8b0ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf49b040b52d5b5f5c103954183ca108e72ab3b9f9b7263f163378d22cb9975073d85dac04ce8cf37d9c1570442c938ec8c582c9e6bac719a472b2333b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7627ad4862fffd2f91e5f975f388a26b38a0289c2ac0f66d8235448487fee7052e3f052b176dab56f4054e36e2f5875ddd450ea9ae63742b4eb150f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9061a32327a4b7f95a01a8d26c83c3a957dc13b39ef2b6d9fedf74893bef8fdadb32ffd81aff95de108e363981a55f01abdd818c2d0637a05b11fe92;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h359ebbba250d9c93555fce41ccaf87c9a58eac3410298e66467fcf9fdfa3bb580302bfbf2dd03f0b3783e97ee86eaac98d8c74e9e8186e2f98b5f9a96;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae48342a19623d6e009e1f4c1391ef91d71e502fcf2b723fa3084a110dde9a01d7273821f80f77fbbb5be95538021520e7091a6a4aeafa7684e849281;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc67c1088d5524d19ce25570c785a9388d1881150c75834909e922db0a4199febde7751119ad82b0945f0e55ece6743d1239b5e1bd6d52a74541be1a43;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h880970e38b59156e1b2ac441c05ed7816f8ccf1987e96ad0e42ec07bbf03300e9cdd7a80b9e529b102374c4c77624275e9cfc6bbb07cc0d58cb3bc833;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h750c2d44fa5422a66030478e78a5d8a6f37e4293acf0132154f14f97c6836483c683327006789091846df4c5c15c52be78b6ce3c692add872c6c96b8b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdee3a05cf8dd3bf8e3982c903f9f28d2482437070542bb63a7593612396199249c9412231f6892fe4a6287a3d249feb5ee4729043a5d9ea80c8fa28d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he33c74a293569a8ed84bf3af4fe406ea282d8b13de74d158e9c35b1f905909b765b04093bf588a5a450ec9333763a87ca6e4d17914ed3fba06f8ca87c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8819be38fc5132ffb8882fa0d67cc1a13aca573c9cdc767dade1007bc77171c80ae3810805dda036342eb47a816af5c1fdbd2081f4bce14d375216dd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc23d1553592e6f55cd9352de29ec7e67217aab747bbfaec2ba3e2bc1ebe8b40a4dfe0b0e4054301e6bdf5f14192778b2ff4574abe92e31b6690ea6e3c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5db7f0424f7ac59c74b7187ef7745430b9654e18f31cbedd8f2630b728641105b9bf7e8a41fd05ddcfbd7cb1d906f31ed03a901bdd3dfd81a4a588f6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h505ea309eb940b14e173d40f830e69e92d7afb4d489c6f7fad021d953835b990fbee10cba569c24ae9ddb8f15caab5665517fce76c38406192408325b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87fcf61f283888ed5b830585472174ede83b286904ed63f4e2a86622c401626abb9adc411a8b73b703f42450c57aa3f9c05f187375b24123af6357d79;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94ef879542b069e2025f6c21a5043a160a1ac5a11476cc8fc47d678d566717ca08b1e00e1a848e98072e963311162caabfb9a6d3510ef800e126bfd2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7c402761d82ee0b2b2d98a31cf87f8f1d80e907115790aaa728978d9702538ab4c81fd35e18e3766fcaedb2ec08de7aee897cfe6aeb1ba0708f74efb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bb2d76bdb8c5a2c57e2f7dbb1dfa8495f94093cd615830069a891e091a714b57ec6582a9c417cba6a30d36199897bed6964abed6161c85bd551ba869;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38a2a1b4d8cdee3bb058deed0a8c4717c57f4a1a85ca52620abdc609d72dfb4cabb495aaa468492680ae5d63543d787196fbf7118731a79fec71a785;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee14b91ac2e913c695f9a0423f46e1bc14c0cdc9e660f1babde114a97865cadc3922c675c1382b59df42bf6eab0b44a6f5776529c41b08b77f7cc38c8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1022cfe15f8598c000ee654b3a26dc485b910e5f5c2f3dc6f9ba2b7998d534dd8a2e8d94c346950a072a36e192f3cce9b32bfecc855a8939f232e274c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb70928904e8267b69722adf5b913edeca3aeca17c6b05dd8f6fbd54c267960f3e22abe028abaceaf6aca21e7877e0a242e9316503f10b75acb1dec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd15576d4c3e0328e1d6807325655d7efccc1028504f5cb524d86fa4e4217dee763fcdc17a6d727c93fbe86c6abdc3c249dc07522f9a3a1095d181f7a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8130eab8360b54c91f0428b8f8c473f8a1121a6a86471f011fb5d6174cc71ef73ff398fcee183708ff152ab461583a0d1e30603ce31b5d9b1b6c11cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17abd7a796210b992949b3fcd32c88336fa1d3e0f5355aac9bd834bf098784d61e1d663c5ae4e8cee3f7d39b6ab77e31e6183846a5044b59b6577d79d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ab4242f270e92f25082190356d3c8911775a053acd0986f5f41d66d5f769bfdbc850c0a292d29c6e2af7c8c264e549482e14cd6dc73489867cc29e24;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25f1469e2a8735398d38a8d1a6001760bd52063bc939fc2599bbf28565dd7199b2d70f1f1b52984453d6727cb55c1887be6489c2d7e34503aa68fe6f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27e3e265a1d159609bcafdb31d233517b11a36aa2e26f766016a7f93cea20336462fc2c0857d826ea825725930fb3d0312345d6b74416cb1497620b68;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77669cd86cb45efac3ba1e89ebeea1a27a57edd5c5b54b7195d4ffd26b77091d006b5e08f3923cf3d15cd1f4ede3370290b0dedd328d386f03c985858;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8820f2f0e0f19574f216db43140ceb912bfe7848d12242cfff33f4391353240cea23836cc639125e7f7f66fa4cac488cccf5a4d8bd483dd62bf0c9807;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ff72a268c939d65ffe68ea1c6b178f2aec68a61c689cb026eaec4cbe390f5ee6747c702c43ebe52b28c5d15c505e01e4dfbbd9d7b80aa748f47f737c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba3c9207ada5957ec3b9abaf5bbc75073be54d0369263073e62e24089e5038d448c5c62787c24874b2d85076640f7e74532672601d4b2efc5bf6284a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1740ad0e87ea04d4d43b2df803d117bba2831c0a98c249f81345fbf700c9021142288bf4d9b2bdcd6456d81b7075345e71f08525ee135af7e12e6bb16;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7444c705d27b83fbfe504300902b65adebd9e32ae91b9e0f3bef8535fef52c339cc0f981ea103d82b11775ecb1c09c254f3fef0ffc5403eff53d73e56;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a78d9cd8ed7c3d5ac08b179982fef39f33b44525ae7f619d4bea6ebec2f87aba4b186a95c0117620af8138271aed80bdb1108b2ea8b0cebd20f6faf7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e641b746fcafa0c7feea12282066c87c082f43df4a916e5ad7936be7d42bff59aaad9baffc67d23492e6074e244d4907c3835dab2daeddccc22b6cb3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3aac98d814558773d5072ed105b1c19a159503597e1ddf36c1501c4983045e35109ba7aa8fabf86dfb47d58627647fe2a731b75482b16fa271ab7af0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f4ff3e429701b94ce9b12840f6d4435fdb9573cd2d99e89b61b9141bc9c23793e45d539d5345be2e77446be8ebe2058ca6f2e9c2a43c135cb8625831;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76f0045e0485e01188f5429a398820c507cc76bbc9f2a888306470dc7e831e848f5f650ebfd8b5e4ece942c723e8db6918edcae623923cbe6e95c940;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3283a32bea268b8f094f290762b6306f394d9f489a581625e298c12d69c97567827c60ecd7e394f69b1f0ac5b610312f7b69048d6d1e82048ea8005e0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf86e85bd711d9145ebdf4fa8e65cacdbd6990890bea1ef94e31f295224b79ca75d7fb17bb438b2af190e087b6c27c0c92447c29eb4425dc40dba331d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b257131bfb29ce2e8987b928d55870ad6c0cc57c3546d98a998ad80ad9334d68d4d8703570d65583ff2e65f66cf8042f38825a2db9dce33493a96d15;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72fbf027b79f4e3d7cf62e2a94fb47d6499d12eb8bf0e30a8e3634d2a42efc8c1ef7cb0ad2cb763ad91c9519cbe08243ca342db9451e41d79a78464a5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h274419699779d19360d9f41203ce27339a46acd15df3d0b28661a6e5b4c833121b8dbb5768b7fa890107165d569f34b0d2f8e86f1dc810221cb90d3c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c42e4d983657ece2e3805e6cacf434833a136700e65bdf8a4e9dd95250a52250c6d2e4c5dd0146027ea83d9d42d74536035ce6639d08216bba787db7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88f5435e1f2077cdbab6ba05e2e7ef9f2bcbe10776efe80d0c39b22965f0fe696f74eb3cd528e2c7d0179c9651b76c95ccd67bd5455d793b56dc158e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h750d916ca560a08d04e5e2c0f0f2d64420c927063fd154558664fdd6d2c453c1cdfed2aa5b53cb3f8454b0cc612635100f6a36e2324a2b7f3ba2ef3aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f49e4d05e68e28b02b528de718f4c324705f1864254b9faf9406c2b71e7449100fd0b4b0780b9409fa4b9781092972e407921c1f7c4307a1977b8917;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f353e296ca45280ab6e0bbc531460d4662d99ee0ce77b131ba7a9e2e2b0eb0d9b8f09dcbd8a5de60004aa761e19894501268a0e4d474c2d90f62fd7d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcbc0700cfb6f31d9f8b5d93339af97d469409c1c19c779779b31a34fe150ea020a603c95b38e23256e8acf6f928ba52e228fe1ac481373c533f9a855d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21dd384b214707fbc1c07e9635f59159965011f6d0421f87eb09288b024683f785d0f772af8b9002a8fedbfa82d215c9376d050fec9054715e91c825;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc196338c46d9371a5809cbd40b8b262b8f8ba4ffdc8d320e4524992c4745d08e6733dea51e2a163fecb3ecbbc63d8ef6aac1d7fa0002eeccce70b6ba4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f1c9c46ef1712b52c1144b5bfb059f305b4d87d9fadbe9c496e1bab7b53c573ed445a32e4822c6eee5e75e6240b9208e62836287690878b9fcf27818;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h941de9d4b5916633b11acabe2b9a8625c23e20cfd68a89a7fdfc345a8722b6088f50996eeadfd6ff3f2acadf281ea2b70c14752a1bcc349c94e56aeba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ad05ddcb8c621c45799e7a07ceadecb4596ae4b4dbe835ee5c1a00c07ae4a012a0489c55620a6763c2f5064a90a2b59abad64e83d9000771444a1568;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4dff7f5918393436212070c55f6d2686709bb7c56502215ad5643a1e0c04824206a2c8a859d802c6ab82c898ada1884fbc52484f11a4df6bb4c602bd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1129ef5165456e8674a52b00fcf51079390fb7e839ad80513a5f12b5d5ff8a529429a1daef2f7bfa389b85732c1e8f555418fdd770cb3d65b50097891;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89e8ee261a76bdfc13330efd7d516aa4e78c6c0eb5ac95f07bd98480c82ef5436beaa6797c7e3c802acfb1b070948e0dc2cdaa0bede6aca2dc14b3739;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c39395e3d6e1f6d959bb10fcdb0689f94e94efb4312eec339fcd986214af46389f41aef550899d5bae387d0f6d9308adc73c07f9d3a9c1af0de76d46;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0423a72656a7d5fdc62d76e44f54bb2e5fbb65a1e191475a2255bbf0e8692b8803b5f8b669a986dbbcb123f7a9683a0f7a1f198aff89fb60b96f2d36;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4f9a4f12ada829a450f93ae0023b5a84750dd9f537a95673d2ef6f5d1bde69997531b630baed5cbe22228b35420671fbfeb3172904d072b0246808d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a6db0090aafeb2b5bab7e34be9c21b8210734993620f7e842c2fb10e7ed2ad2750a8b960075e821993cd7fe545761b8d941be9f06ac2f9b51b31a062;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3fd52bdbf8d4bed8a40005213e1dbd24674b33e52dc3908fa538961a4f6a43df463c937330762907a7b76efd5ed638674003a16fdc521f91c479cd6b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3d3b03facdcdaefc1b5ff49220237c6267f3bf78b717005cadae949d2f772a75b9b14c0cb3da3d03a759057576f1f74328ffc6171d30fc11a7ea1486;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf51866156a6ccfc7f9a965f5fcd373d71ef6d88f5938a48e5004534c89238eebed2d0a02f3c50cfe4dd159298cba572d781e6b1a43432b3c841df1d42;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65ead36bb62ce8a757b5e651851bdc4069415157416a603e9710b2ba4f3195d4f2bfffd127f8ab0e6294bc958bb1a79f206dcbbd5a78ca0c354a11ac8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedd82688221ba32371c6b12b355a1376814f948b1a5f25285063383279bcb5cc93c131eaf49984039754f10cf86ea41e79449c477ff46d1792dc12da5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had3af755c36b2a17ea053904d199e4bb272faff5b695ef2fe4990664398beab41a0f0f2afbfac7df59e47b1ebd66b28e129408566615f0d6646f0efd9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d5cc2d655962dfdbbef3724cc79bb963b4810fc22710078d1b0faa5ee88f15625b64ffd725bbcec0efa8edd5f69b00a3296653d109f024b968edd144;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6734d6c8c920f2fbf27dd7916497c9ef96b81d53e79bd44fe1197f9fe33696f1e901822047f0aaf6371f4472086241e38d093662642e841ecf45c71ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h662b374a59dbab7ed757ba99d498f82fb6ae8ab1ffc2298799189ec8209f5d12c2d7a5d034044d83a36fd026506d332ed700018f304571ad26cc52169;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e189b68e7e31906e57b686b1513fcbe6eeb2b7cb1ce7a8ac3b526c14c53d516f2ef7b9a18aa869010b5cadaf10d466e9bbd09b39c898065eae2181cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89201081702a651dad2f728bd64137ff2a32db5420d9b9839242fb1475afb9a715ccfccca91158ec8a4f9d7d5a005ffb31eea69434425ac324e5d9cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h428f19057bdc1aacdb4ecfcd01f30055097299642e1eab347e7a0f8a8a190a36d008f1686d7472d17b924dceddfe1df55ebd60418dbea899573501596;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fbd554aab3081e784f38ea6353c557103c995bb6f452b7b69afd1f413100b8fa7d6da1c77a50337f0230492cce6d658c00661320b82e071565f40603;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b5362a64b599d2347332271eb71fa0f94edc13a478d1f577516a1fba408d00d25aee01433ef12bd1eed617711e3f91e18d8d89d1f060c98a5a93eeaf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9e266024b2fa7e84f198c8b0b07b4e81f54b0133c2a4cb41620e51a8b714f80e88e99e7b6afd930c82c324a0f597ad6f879a09180f87f407dc1d56e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e587256feae28530de40868a20e27a0604d373d366f8e8cdc4ed261f8c42a116d15e3135fca5a6365e4e1bfd0e314b37311730561f509c50e6722c09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haee1e2d7dc2e0488380f0035c36b63f765a28fd0f9042d5d77c1e924ab80cbfcdffd8ea77381c486e79b988c9662050ab3a7af9c2198daba71237085e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5f25f6242723cd0ed8b66be9ecdb617ade5e4b10cbfcd67a7c045bab266442d04ad8c572403bd1a11c4873f9dda568870f76a77d59c3eafcb0faa785;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h912d61c203e42a2ca21d0cb7d72394a7715e5ef56c0f962a407b7172c036aac7f951da1b1653567559e260f4c6956f3a0588066bd06634e5ee0447498;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc17c04308c76efcdcd8e327f6a0b6defc156a6bf3ae788ba5812ed8f98061084a404be9bbe92a6eec90c4b0b4e901a7efe56e0ba69d54a39a0f9740e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5fdfa635fd37fcf628212c692898c9b9fadb0e98306a720bb758d5cc7813faa5bb7a4d1ecbacea32f81772191b06be4346d4f965e3e6e8c2fcb24619;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87f22f64b931831525c2d6cf6dfe729d85e9dc4403169ee24196363fa805432f7cc080beb920c8b26b5bd29b5d14ff8fed4e882e16f89d3dff0e6f857;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha569e5ed7cb9f05a8895f0e9fffd9f50ebb680c7f78efee98bf70bd4fca052b9cd0cc06f0b33af870de7a3b11ccfd0cae45f2d3916f0533e94457b24b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5d76f1cd5804be0e774281b6f0501499ae0d65f7f95998a386e0f3376ca358f94f11bcae968ff6fcb33a1389fd30c0bb39a3b7b07f124c8f8b938306;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9850e1f53cdf11568bd62d7b7797099dfd540e3182a8c322c3879178a8add757b9a5946704fc33d891f4c0fe5b0a904f980c6fdd75973ad38c34d656e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef06de503f41fc05f52f417f38a2b224298e4ddc002669a74a1a581789ec5901b4cde85238c4677f023f115504391c70bf0c583441d5e4b47f9ee203b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17d88a74c8e5c571fa70e2c6177520dcf68687622f08788c1e038557c15fd317bbbb73255aad01762bd75f2fac4def33dd2c6cd6ed904500bee1f03f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ea88a37843348d7b26282efbfd0678eed2cb04e2f3fd011279f89b53c1988f9607b3a34561aa160ae393e3b15591bca63a944b74425138db4771050c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f297d8147f4d36c9c56f9195a041f68bb8414c1bd0400c379ef2b055b2e7f784ce87c7ef6022485a22ac33e78d156009676b035b161b854906c6c75a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce04f50fe53224ccab0f1403d6d8c2b4170d10ace7b19f1ae2f34c93da45e96eb3121003df7d267fa31d0777fd612fed0cf2ba0b24e5ee06a8e5e6994;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc43845b203fe19b4ddbecae07000c4a25843107e07f71bf5c1a51427351206ce60f5f0c00040c71befb297aa71ef0b2b3d754619067275881af17528;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bc81fbaa46ceaf49ab2985a87506ddff0a391e00a46ef3456682076f8f1729078d8d3730a85949b4716da8431633f2ef8f683308ba8139e28281072e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea456b37a157286b254ebcd218b61db93e2984393f8a605ce4caf85cac9da0e76cdeab83d0bf8f01f4231e5dd657700307edb5c765d19112479f7ae96;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he23b97ea2182311c1d5e4a45b473aa234906ffa81894c96e261ccedd98311e22017d17f493b6b99f73a2d0deee338059f3ffd23ae7bc1511c489a7990;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43850c15103a9aeb9f4d3319b7eb29fbc5f22842c84281bfec20373b1d3f2aed703df56f02b7bc7a1d238d40415b714cbf9de0c76df4d8f155510eb08;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56a79ac0c8c7f06ffeaaff47b1754e1f8c72bbf0635b737d97fa4a30441bd52e924418f82e5ac07ee29f401c5a6249ea2ecebe9acfd17224539278bdb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h982b47ae765bded212eb82152e7d367fdafe999ab8db1ced237b5ab89a46c65f68cd2044e7a48722334cf30f3e4c3b1a0513b157aff948f9f8993c025;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefe990e181164e135604551b835dd516a3dba8571f06f9e6d9a737186a8b729910f92168b3edbbc2b6ddd5eb8f72f9a4c96cd6b7c75c7eb00d0e068fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50c1d9e50a255ab97afd0e05348ac2710b3d250ed80bcb7e1d88b5a28de4e4b48b28091ec3d15ed0b0ca97f9771b2804804611a5ae8576c287eae2947;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8c7ccacd187648e9c8ceb18607e5fcced6b5341556b55d0782d1bf6855c8e6d1dc72ebc931dd75cc594830da7d4130b43287bf467dafb43e959d0125;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6761077c2ea077191192b97fe99c7da23e65a45fd28350fdb5210a77d7dea5cb5cadba26345302665d9983b7db35737b1ca0a33429c1b9a530cd71f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ccd02b1ba8ec74bde39bb1a8111dc84ac9e78632200673041c9c7e6cf1fc2ba473ae1d438fac754ab13fbb3376bd97c1bae1c6d830597439a7fb8e4b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h110202cbb76f3856d8edff66aba3cad77f99e9f76e9c4e310828215b9349b1951c194b882f88e95b1fdfac0f71f385afaf4f7774998551e9caea0fb2d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h472e10d995bf9100e16579800decc5385ea58ba3befb9211e877a545139901284d61a878709271d2f94f3ba6efcf8caf4a01f6a258aa1a11d12fb7e53;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8c506fc1421741d5c64311fd2700326eac1ae05f75e0e3709b8b81956fb75f5636d271241f67092d480252f086188cad8422e3c26950a8b0f5bb1484;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39c82726a17623ed3dfdeba43e96300e91ec5940e6e547da9acc89d26d1df23e62f3f2f46091f85a6aab53493ca4dcf4c7f4b2226feee8020b99a6718;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf66ed07dc28479e3a60a7cda9f06fb4a961fa0ffa361d751f6896bda01ecb335f541b42eeb9da201e813d360f8ae9fb1cb737804cc91dfb880a20c7bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h159cf073e25f86b17c6730a0a6adfd62006fb44bb5f8584373d2d87248a045536cef9d4efa3f56bb57d12bb96f4a719af0a18e21b8f8dfef1cf8ab348;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5cfc15748c97a0d5e133068f6d4dd456e7468afa0275875d1fe5e347d12a4e5164a8065d23d7962b3b7a5fab1e72942d1ce305f073d29e3939e694633;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1673813850fce73ca740e5ce1dd8e6ee8f9160bdd307da467cc02c4271b2c8c3236b6abb57c97191ad4c5e05210dbb5b9ed4e8afe121e0dbd82eb272;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf43be8bd9716a47c2b37e0984c4d044beeb8669efb77cde87c63266543cee03417a83a344689de3be8a3579a54de8e36029b7a5b2900ac0082bfc5f90;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fa3a6815691e616e8d782e11436f418559655edc0ff3b0527bfff839c5dc207b8560b896dfcf309c007b175c4fcb9388c399031436855ff240e0a0d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac09b1500f32052d61bdb4c40f2b0998d6e0209573c2cbaebfa04318e02c820965c9b15286f3fd80a8277d4d935af804d807a18eb647d55375f985d02;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb43ae5696d269d5ea747f5c437f8c218beccc49f37280dac23b6517eccb5aba55a028a4610b1dd1b9b88acd962cfc1ca3d8d010a1ce6fadcf362f394a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87b617802e781f234f62601fdd82cab59421b55816c6bb02c7e18c32d92559bf6e44ddbeb01dab326e955669d2407a0c87d147f5cc926231a689e3190;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2abe962b3f57be79f96bef872ee4182ac5c87c71397c1e3b40bf7aea9dd30725c54321a22c870054f88b8f6c2b373ba9fecdddb57cd650f4efdfd19bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ab6f522d9f671a4c385344dd485f222ca7a693a0aaf508d29ea7e0daf6defd3a362e34221269eb50ffcd02910f5fe2692a864ed3b9cd3550c0c301df;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h584e914c2833c999eb0c9db7ca645ee92116f09975cfc49bfba364e4b9ca7993aa0e46eb6c1566e4b8f1270a038c5272e512c6eb3b27fb183b420df12;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h702788d5b949c83989467ff984ce363b57f6cfcae93628969ee1d126a07359c3fb16a3da0d08d44f1cdfe84927f1a07d835d57949a5891ee9a0652cc9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7724a2f144008315bd283317a1a42267a66b7132cd072341323620fb52339d53e1bf13b2a32f137153b421149d8d408149c5ffff82db05935db470f4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h307b73933a7256f1485558d66f83e83c17eb2ab3eae6a948a755bd4f2021dad63ed1c5766c08daebcdc7b07d2f497c0ef4a9e6ed2a39df28f3cfacf13;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82d7baf7ff10e5f26a73456046683a887f8a4a05ebd63efff6bd4de963a7b753adfb19de32310d3d7e9ba07d5bc41acf161d5f0d72904f6e960161c44;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd06411af3f19f02c9208dd1cf5dce5b13e2a05a6d81c297a002eefc95ed8505cd70695ba1e7591f751cb123cbdb1de4884613f90c39f4016edb2e6ea1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9add8b47a16332c6bc35947a7dfcccecac469755d9be064d0c056980c11b6fb99c56341cedaa637bb57845d351b9cde61d640b8f97589276b832b29dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf540b4467f7334985d7f8c862d7e204cc125d100b4fa1c10cdbccbb93166091445fed8d1878ab2c38e94cf21168e91710b9af840d2f3187e9a17cdd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e5c2cc1f685f05a358fb451c6780436a2113e250564cd90be1cb118e649dc8ba4b2ddbd35d3e22a47c88a6def1f136159f5c113c50035bb538759bda;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c9ea7ec2c6a9aef8a89921c720606bd198afc7bbcc2bbc70c3d0c3eae7af865f0ca5cce429f4e25956af4bf6d5defffc4cc5912a088c5e096c568040;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed5cb55d0f3d07f5bf9091559eaf6d0ccd36617df53daee9dfe61b9706c28db9fe520aeed69ded9edbeb01062120186cffb75af6f42e91430477369f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc18697696fab887a05c30070556f9a49b0cd1e4c938417b3e12eacdf2358f38e5dca037202301d4ddcf04596d7c678478348da2b7e92849ebf7a252e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b065626f9e65bbf191ee1564ddf04463a735d7b9eacf417211c2b26ac25213159cd2442b09e528126113a8d4ec291a56585d8c41cdd42e5aec5dea3b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9067c482fb4b5d9f13bc6514b87541f04a7e27344ecb28e9ce4fa014907e1c7b4e9a71f0ed2ea5a3d85051af37a498a9748928bb4451a91528defa887;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hceec058570bc09c133318e2ffbeaa3e2cb2b4a6b8d080b77edb712afe12088f5b288f8559b2f45dffb5e7dbf3ecb3bbde85da09e8e5e060e23582b79f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hffc1db1d3a4b9de74fd9f2f2371f160909e331b4b8245677446f9c310f63ba1e423ba5e454fa4de768bd34c324999cee334eceff2e29c4a71bd134c21;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h398b4c369c61956c8353a837b1cc893fd80b7d27f50e5bb4caaa8570dae8d277257b2a6f44d3c390d39ab4b00746f31aebdfc62e19f6f80c64a884009;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb57498021596a3cfdb9bcd8e46be5c90021f465b46fe3dd554ec48024839d4a29b3b1a2e6d4abc9c47177f448a0097ac4e071ad63ba3613e532a5650b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc54071fd85a3ee9ff77f5d468863597f3c744062e975f821c3896036f3b9c45e29448df4363338ae391cec40a06c4349006d3fd7c47ac3f47275972f6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46d22ab524ac7903b8d336ecc2fdc6166c1a15b543767bc4928907e906d9ca53fc5d8e314155738fec78463b4c50aec22a840d91f7db5d7bf54ee3a91;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcde932d11c0738b4233bb951087d5d6cf9e7e3c144b019b0f2561d83881619700dd03639bd61da123e702a65b2bfee73b4897827f0a3bcc04c91b00c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38ac1152789e95be3f208d7a992c944dbfab5d24c35817875403fa27fe2d23bf82fee589f7c774837c102f58ef94aa4539de83818591b62bf4114b142;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b16a06150d068fefba7f23d4b173bddaf604c74c3b447b244c3f9f4bd5e71142125d21f69c77fedbaadccaed8dfb0889127a59a5d696feb125d97b7c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30dbeaaa9b96f44c39dc65311fe98dc8cc756fd04a368fe43775d6fc298ca3f5dde7c2c66eae9c8cf16033467e875833d058c6ddfb94c522b89e06638;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85de71a7e3e8b480b83455d18e07a27e2658ff1fde4a091fabe893b920a1ce54baf43cc0686cdee057cd9a2254a7016c61988029f24af3e0ad66b332e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f572a365e1665d5cbf7612caad33966d251a49472a41ffb793ae8ab91cad200eaf2b322c056322f192bf52292f0aaf1e01d9fb41b207bc9c8b0a5f6d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18231fd71b2a5461fc7dd3fce8e3c54f9582a7d6c066aaaccf5fb23e5c02d852c93093b219c03e6567133c64c85fb621fc6f22b487082ac4d309acb64;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc795270fcbcb48997fe887c8d26d4a0e40c216b1eb2ab83a3094ea53c9cdc29999cdc6cc5138f54c6b837e280c44bd4c1e7075eb36dc8aa42db5b726;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72d16f0d5f0b02a9d8618c928ce083b1f83fd47a95dcb36ed8a804950ff80a0dfa143b3cafe43d435bdfd52cff7b01bbfecfc4e640aac118619fbeb74;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37da4cd6902ec5a40c3aa1b644ba7d51c38edc7ae80546fdb63ecbbc39deee44f4885dbb0dfc1e40e1636d2ac227eba0220f66dd5774138d1abc2aa89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14206c31cac48c2872e9a67d63fb882721aea4576416ea2201dee4c939848d2eaaa525d28f42be1e9ff4dfc6b1d2256be75242f54c3b0cdf9ab7333ec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3566380ba0cc2efade57beec94b1a09a2cb2305dbc69328c0ea82c75fa5b19c58eb36b2aee5f4e665ba480600f7e5050b79223907e35fd742ec5dfa4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h562d6cc00ae27d83ef6642b91e529d69c4f6f3acdbde4b5d00d93528e4113313037f22b97846b397cb4a9980addb99e4bb8660f8d6f9c2187876ae61a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha63e140eaee45cfa77a8c64c95eb297a2dff2faa774c474919b6aeffeb72df1c66154a5cfab50f06e229ba013f552d66ba2eee33f110abf4ba63b7e53;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d65bcd0044f7314d7950632cb41a4a66f5385f8a10bf421bfce93bb5c45f6422cfb98abb6fa3fcc71d40a811721ce4f3ee4b7f3b71dcd23666e5d1cc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8140cef085290614443242366356ee09219d3037f277f7c027b4f2c3bf0f797a31f3fa1afe4fc63bdabef15f5d2ab007a011873ad199840d50b4fb6f3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hccc185802b723088dccb39bc63d24db3947886ae88586031d21369268bf577808ed026441be8cc5035857181d7a97679786fd0cd99d3add8ec67a0ff1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6e30767950ad4f690ea7d3a16ef0c113f8c6cbcb466b45140d64fa5667b63ea470b27df0c4314bc9fd110168feb207520f991c7b725a000d60be0d7d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1daf288c82b755d10b23cfb79cd1dfe294c5990800c834a1f3a4c25452b6d077d52308b9dd9bab782536b62f10e4b37a0cfa3ab6ecb68ea955135dd0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8dea79074ef672d1b348a120f5093d1ab2392c240df9e3a0443427c3f01bc82ec2e5a91a8055f34ecd8647a9d35cfef421815dc39e2664b81e2829c23;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbef6a45a11d11ca76c3ce4bed78a706707e1a8451b1ca3e8488d18611f1c3314fa812a4eb1ef3f83e07e0a0e0fc02dd0350672342abe0cd7180b42d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h434f17c723a45de29d53971ba67810fb811ccfb46c58a41c00ef8a439943e11c3bd774c7bfe37ff0e8b7c298c4e333e696345bfec7e239da5a2c2bd84;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13b6ef34e44557c669eda4bee4076e07d8464c6d208a2b735d39b7aec3fb739a1f67cd0780bf3bf49256306a60d2988f6d5a13ab4b757df985733b48e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1baf68fab998bbe6a201ae9897e6067c36024a6500f89f37d0c0c99d7a28ce5effa598f4c8193554d178a88f09fe3ae61570f53b4c02aa9da57734e0d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95536fd94ad2adfeff62f278123351909ca9f307addb92861f4fcd54ebdcc1216e08cb22e79268752d7ff3b6664c21cf43d18b402813f4fcd6794cc56;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hceffc35878cc2f3a93de51ff2fc803156a18a363e898f31973c0ecf83c9ba9008369b95668d816d41470bc9239b5ef2b62fd6df73c1f140262e9b0cdf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce5833247011fff6c2741f864785d1eb73ad37a8966ee85efe94b825f36f44948581017de6f737ba28e4f0531d8f5512bf4a2a5239d97cbd93f55926;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe03928d751c33bead7d7984947ff09dea8b5768df7a1cf64d42f13a60d060db752a40098714f8e04a7d70767c26c2153e5011240fb8f9a28c336a474;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86fd12cefd4e9acb318322612a062cf066737970b6321ada72ba1625ac24355783895e3350b618d332cc7b91dac34e91480e5ca36f38bb3fe3fc3306a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e5f182e90c7a7aca19e4d832f6203f5839baed25f7447d813f5fab9b3f97a33060e2b9a44302ea9cf56b8c9689cf8503ecd3eff26fe124f9aacbc16;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2af0922b3b23ee806a01aad32bcbe9f547147a26f1e5f496e552df45f71c6ad94cc8d1f270c002be012edb70adf3b62558afb4e7e2acce5c800532d83;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d5f6487d6f9d01fcb9dec142462b05a37b1896b3bd9b88aebb7710ee120b788c8770ebf7450879dfde3f4733e4675f4cba950f8def4ee6adde40ae76;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4648f2c168b8ea97260d250864f463206d1cdffa6fb6101c45187858d83dd2e8b6ddf553fe0815250064f4377bcc3c1ed10102934341de719b914e38;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf3d23282c8604544558f372ae7208d0f85f43da19ef21ef64e57de9a724e0ca70c8b2e90d7159482955cc1722abfdb4fdfe9f13e148e6372a2878818;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69469cce9e042e9efc103182cc73a3e3ca4e3989b6b7c44a4b86a5ac551e5ea85e1d8ce2ed7d41ef001c66d366697e36051fc41b6a68aaf0b0072b87;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7422bf94d56bf91cce98be2f3cd674c41c7894715ca89e86c7e9be781c785b49ba355dbe95c97eaad926a4d0e689b6d7af28b202eb7631894a5f8d08;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62a223c3f6f9e4d0c75c58a2e6428f2d7b7ac68891b4f53f3cb94afb58724e2c6b33a7dbeebd2e760389bf82f0fe894f3451c82e23f22a65593cfe458;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa0da0edd00f52f7dda0dcaafd6ba1a56363eb073d3d8bb12e4d289fe4f775b7178b3a737a67628e86aeb77ca4aac4c94512f56ccfb27e58652dea38d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde49f8c366ecdb36f930018bab4cef69c0cbd43b6b1bc3834947f98f3f328851e9b6df3fb835d3c24a6f9965e017541bbd3ea04ce77db55b098b23d8c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h219574c1c19ff06b2b0cc4aa200ce092352edc1c9822a0af37adcbd9005ab7ad5b6e7ce8f6f98e78171708a4ccc475dd9abb35c99312b14346b0c93d3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92e2d70bdb1d2d24814620c3d320b357c0ef4ff816899fe37cb9af59a7f0966f11d09f783cf333bc5096096827a2a6c0427870718219e595c81b06c0c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde1844a1d790b8500af450bbb750fc4f988ececb8c5ff420c0c7c1f9334e45b031ff2a52c6d5b476feb48c937281c92d3fab085d9d1b030a1503aa48;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6760fd40f6e1c33d228c68f455f82cc7d53689aa79c6a115a9c067c6caf145a7adb1e6e270bb8148fb8ab047c056efeb5197a7bb8c54af53705df1754;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba6fce6c174faf91375e52e00ca6a05ef81206252d3a552daef17c34152e3775a1b74d7fb8b3552e21d3abdb31e84444c7fc5672b2e0766d89b763175;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he420d46e5a9bcbbd47196806bd72ae3bc928d243b3a14ba65cd070b6598b2005c5290d0ed35f5098f0178a81b7df70a97b03288f6e5af559144b86eb3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f02c9dcb1686c34179ef4dd5dcea1a242e7425732e2cf3c58e443b9e7b75eb975a5b1d351d9fb84445c763f599a05ca17b51b929e4421199eafc469e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1126d4bf81f9ca277d941895ecf24ecbfc79ab75449cdd8558dbe0282e13c62592ae967d0dd50b44aa401210f4693a09f4afdf7b32a0d9bdeff2a451f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf33588efd2f6c580d54a0a0f6263a7eda953f0c98d68ccdd2e6d57cd446d5890a64164f4c81db185d5b124faa343938965295c48ef57b001e1fecc223;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcec41bd272dcefef2e8dfa083ac209a50e76e70afb16bbb81ad08b5d46630606b29cce0ae5c8804edd223cb655d4ca7916ccbf4d0a7756860a2b2e9f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6298aef46c0027366a1d22a3c4afbae4cfdf8562adf8acc74aa3d004490b614edfa9c6a13bd91ef89a8992ac6a408022c99c7c474181d862c9e94de8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa73fde39ceedd813b6b3abcff73052bf36a4b2bf27835360ca0ddc502781dee76a1c88ced8c8cf20a4f1587cf251def0657ea10ae0fc9ae04124fab7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9befd71bff26465311c682998b85be847ae1d30514c29590b906d16691a85c687cade5631b9b2a229a6da419fbb9c9fd617b41117314f727fd4d5f0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h760b44ea4d2ec4aa38e8c3e8e85d8d6c182a071c52423b43be6374bd27c8ad1f792be5b8bcf770fbbb183a4dd1d9538ef762081812f00ed214287428f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb614b88f7efa3aa7b2887ec55ddb06686a438b6b8d40bc37ef5d5d582dac0ff37910a67792e9f68813fcc4a8689dba5bab1b02cd7fee9e675db06486a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d1c56dd8c9e725932c9421cd4f1611642c27de7b8ca0904248d6dce2efff00068ace74d10108d9b01eeb8655bd6742684a8647dee5cc29b3eb82fad1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43959aea8cd2e471126694e6e25040202611ece034b698cdb09cf797b0dbc5630105a08178ef30589d3bc5df89cf09cb8ee1056230688b77b2f65b9d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h772b47d2858813195e88b07a7626feabb49e929d4dfac6af6431fbe0f5e386d89fd7f40c65234f191a458b4ee433d27165a4a28e1e0d7d838884b549a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3f99d196dec308fc6bbbd12aa442d21e2a4967ca06982dde91732baea869bc95bd55cfc37394b8764b8af121a096e3f078dbb2d6c7e27e09401d7150;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbae1d263d087495950513513fe1a284a1ffdb2ded074cc8f026e0f1cc63928fec53c3fc2dfc6468b60dd33f33705937f78ce298215c3635a5e91cf5f6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd96ea3ed95c8f1e5af6d457c3b5437f24e3de09f287e3c5ab4d53f83f3ca3f0db8dae5b8b16fe3d7ed340b2b8bd5bab29d1c9ba329777c5cd836bf98;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h550506bc4296c7411fbfceffcf31adf7c3e738b1244c765c055f17dc93ae3687e4536204c8b323e32ead9b8b884cbb306b9cb1536930c5f4bf056fe35;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b53c2f4c71e6a69d465595f772e84cd6773a3536594f26767c687f3d21bc73a44b114551ff2cd750ddea4af116e205fe7012ccea50460ced8870cd10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haafdd409cfb35bdd4fc731d13ee42afda3d367d557c2291b015729a2bf5241b858bfc528fbcab9eaae1961a6d1673049861d77a60aa07499788c0a34c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1acb5e63cf99a6de47870a1775e9ea65c3875a685194ea5656ad1e2e8a43414ece507f7dac9354b9ab7db7d168860c5f699d1ff8c0c8ae141160ec51d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he096bd9a5a49809d5abf001f0ee28c03919f9124f811ce66a8c45c4456719d005469e09503359c761971644b66e7f9342a06a4d0f85be1ff6bb24688c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5f8fcf60f8efffe6ebdd3b1de22d802af832f341e72cf1e2ba86d97ef1059e0d29240427a2713e12efdd07ffb0174a437dbdbe7bbe067f9fecf96e5a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb364d014509140666ef99d96bc6cc478936ac1fe805e4266be13d776a7e0d06331ee3cdc91965b5dd68c3a56d7ed94c9dbbb3ebeffdb6a15d15a8b38f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0e8baf87e22913a87225159642ebd37fafb733ead2504439a1943f2f06958df83696b031ab3aa930814fa14fcfd7a8720e2dd0272a3c248de0f16656;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52e0a6af552e6c6ef75ab6fa8c48ea0a69a907e913e93c858c5ea29f9f326eb1d9a0d44e63872f42008ceca3815b574a41882678aa246b78dfbf685bc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3dc9b8f655a2050cb8cae6fd4a4bee4609700148d3c2fb82a40db2385f60007ab20945fb11820bfdedfa78dade5138a25dbe5ea1772530b781e7fb468;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25277c2efe8fc7440690a6b3d890b7555bf4c2c65d9f274cfe329b04103ae0330e101c3ad2194e63c9f0fb1d475fb9eb70412b19fe6f60ef576bf7fe5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8f51443bd534724ea1ffa6cfe373f1306dc799cb0b34d57827324f3b08d155a73541da87a3c3e1c886ac273b35d376d861a247cfc0a145b65f0618ed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f9c46a699369016b67de39303a5d9fb24fbfaf7c54040bd1689ad6d24b916b1a5a041a219db365f08e50e78826ee8b1e27ffad0ab92eb2dbb9442bfd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb384cb5713709f19402198b7447356e43821a73addc494fc662781dbc33833f3692a4c23060cb66322a727aa9e41f9cf7932fb5bd71498e2611cebe45;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd60d10d4119d53576f03877af01c170ecc6b35ea3f450043f92dd1510dc0eefb9829a1c42837650aa194cafe2122046b5a821142d0f6f6149188c6930;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf4adbe90122348e6798655940414f7bc4a014068fd467f6fc3c22cf2e67b182e098656ab5954efeb48d0753b4b15f67e876ed885473fb177a106be44;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58c3466ca7b67654b8130cfba294b23aeb22407eaf7ae8056df6f26f3b88443298bdd7becc5cf4e18490cd8e82baa6ffd764123311725ee80e85f2580;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbeee0142ab1c5aebaecff1379d8f33f2f56a11c2e6bf851f027aaf9234abaa6b0abd422db8a5297f099a3ddbe8512f8cc2c2f50ae9943ebba9e05d97;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1e41e77de4e9b5f1b782e37cb755523559c096c28bc001edcf9dd4bb440e96095c4cc97fad116b255a0d844f6f060127bc1a6557cc48171d5b7f976e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92489445d2c26293bc1e8010ff404f9b4e74f883900e4ef5e52f325517d9f62616b761a9b506b1d66a24087ff65d609171aa35589211803fb39923037;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bf3c32c0a9508c347bb1efe9011f13bd2a81cf6f24a5759f6e625374fea5417584267dde42d307604b6817a6b301c4c005e42e50ab8ebb2884def603;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95432669a98a883cd03d8ceb466d034ed09e7fab38287011c082068e8a97c3c9a74a94ace1d78376b67c9db10be856a7b81be0df5be11fdce1aa93787;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ae68098a0dd7e2db98c4f0973139c312e34739ad32326a418f75bb045f93c33bcfff79662881b76ce2f2ed7cba72b8a0fd686560bcac48c8e929eb6b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab80b6ed6be79beb59026b1ce5ab005f08a1e621831d51207b2ba20479597cda663edf6bc4ef1c04ca9412392c98e98fb552571a0536e9277d96b6755;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h863f22ec0533e6b2fad01000595d823652575ebbc8d4c50fc239facd9e48ff0caa77bc056dbc6476ad897fb1cd1e2e50e40943b09a440f1cf016e6772;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8051628e77ab17868938081be58ce6f6d80c0fa373fca555adb2dd9d6e7ba1c36a06570f0c14d43c77628c226561d021afacc13cbec81544d9918b926;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95ab68c680f05d4a2c59c53a59812cad64ab4e9239260d1a482c71059451649913b2565a5c1823687c6ff2d999eea4871f6159e4b13e3ee212e723b21;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49de5de3c099860cafddf6ddb55dbf7c828cf1de16e5c9d753faf1d10b49c75fadc48b7e110360490e29ce07d42245451509633604085284243d69b13;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6665af48e0527dba03b1207c4ce0a6a8196e30dfebb740b649659d8a16a29332da2da5311263177d2e99320a06d745e063cf0b8afc2abd6b77a892f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16f44714d6643e009dc645cfb32d3e38cc949e6a099e8b98678dae8fa81bd554d1d01544787876b1d2a05a366c94ce6512f82c34887b23eff90aa72df;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d731e0f6f89971f93d753274dfae87c886bdf145009acd78e4af41c662648b9d1036f03881fb13ad72bd4373596e9f3d4a5a076b6fe11d3f2a1bb6a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d8bf09a4afab82ce840077a8fefadad86b3703a21f2d32533982bb239580ef114dd2a724a2f318c05333699d025327282a7b6a919a76eeafb2d30b9a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97015a33d87f0158da670a6395c933995d4136243810696be16f37d29b689fec6d49aaeb9528d260255c86cf12bbcf52fa18aab3476569a412f622674;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacc464c543e64f5869e7634db8daeb4f714ae704de36f3efb86d7a506ec5293ea2d31c53260f156c74bfdf9d3e631cf2a1e0fa27b4a2e30aaa2db9a90;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd28c1f8854ea5577fa5b5e9e4a90b890088e5077ccccf28e5fc08c17c7eaf21ec47b54d4a63550addcbcedbca8ae700e66b299ba68acac5e5506324ef;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc673ff15144ccdd9eb18bb719af4e5cd28b8b1525893702cb8cb0f88bd4d3f9113eaf6139427bf3315637f4501e12775cb3eb5472d8ca05071fa19d0c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83e9bd0a6488ecf6f22924df78c0fd4eaa1155e4e0fd2ce474d173fb09a3e359db77e7826eb9545c6578d9e0ba9484105f155e82eae108cf338e9b840;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb62d61e6ba7636f8e424dc3eb28d3db68e8a2ad2cbf8865695d1d49351d21cf96681a6267c1b0f85ac97899f25ce817a0a9e4b0488d4b3cd08f42b90b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c83e7d1c6501ac67df45a8a69bfce09f3666c2805e80d129385162c981491352c42538006c4e1fe7c2d2487a2922a28e3023791e516f6bb9ddebca2c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1156a4d62ab4f42c3c15a37de515a6e4bba9373f8a5206726b42a29fe643915b49d622932a12e40c5ff9a0f958af4a983a990c74936f9a194395065e5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5f967b39158cc17adc921c9de000aaf5f99b5d31417ac5b8c8fb587a23a185e382ee85b374ef70792b1b6f12290231c223cb9c23b7be019eb3f3bcf6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fa23face2f114c50037b40f488aaa57140f507f7c42ec6f22acad7b12e3c1b31580a3fc745c8e0170a585dff3277f3bd0dc339caaa62003bf7e98998;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h235a8f67b4e681575b8a95251fde7ea8bba6ca2502b12dec735cce0f611677a999b2830c4d908769be4d98a3bb7f3573db4c3415eb8f2b7df06333b7b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf94dda4353079a9c18a528d9f9c96f4fd323face64e9efc8b93785477bc268f00cf63a9048a522610dbe4206c4d5dcfafd8064b72bf8632708e20d3a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e273acaff458802bcace1e1bb468b639983b657bc3468148a85eefc0e95f8c5e64e615bd6615f2ae5f2288aaa06045537ef11e98b984c32411b55a2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3635b275fecd53ec2d65ab6e7986ca2b95119c423a2f1d9bf9f5834a9bca98ae4a1124f1d736f7806684fb33787501288bd5981baff7bc76605111092;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdaa492fe9313a7578c2baae1fed883027adcd98b043e88fb050faf091e1e7ce84091883400016e4c0acb902a49e8c427f434b0dec1c11bac0a77dedf6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h579b187581811b7d36e82cb3f73f5e263f48c88056b83369903e517fa81230f5ecef3115720eab093f6e40f7a659077e88dc699088970f138d402f212;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5e7509db25ddaa1e275bac6c52faba5e66041a47779c6507f24216306ab97987cecc402521942bc4a3ea316c7c68e715160ae2c2bda5a62ab5d51938;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h181d8afa6ceb63fd5a81d22b8e82d9ca8c547595ad49cad7f693e878a4465de9c8730252e88a09fac25e12d856270b5b5975f6730ec31c72da618cefe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9eec766c2bd88cc62bfbe8f1280f91c4434a07931d31ae231d0fabd0a629d12e2f76e3307d49935434738b514d2378e70e924273ecfdae1660c78b04;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3e46d0a84f7c930dfc16f8743698fe3bf5c6d6054194e31c95a1f3f2023529d736242127d8ce6e51481f7ac04a8b4ecd0a75a12de57fd6d9664848b6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had2493be65f75d9a7b74cf73ce092299f6d9fbd118a989ad688005fb5d414519a2aeea750e6a1588205c30dea8d8955d32043903c8197cfcae0535ccb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0aded091fd58ba19a29be136d71d323e9b4b92d499675a4a8e216bf6927867f081232c0547e561d8e94b61a0a07a5ac42ba763705e23ad81636bb409;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h357d50a301aed3d0505c9c48fe1a17c3e79d7558be66aab57b4bcc48554c0a420a2ea2883f35dcefe15cb03c2318fd77b3db29736caa4f019bf75e2ed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5cfc06e5b7264659650f78632a35081540a26c214fa9903bc93ab2d52eb517d3112b3b1aa4b9e5652b02d72196709907b2024add2cf7f7c1651fb5e9b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3abbdf20b90320bbb88b128dccf52d3a8eca2e06813fb765b2c7cbfff6a402b3d77d60f86fb6749cd72e36e8a755f1ccf0912a94014c3cc11f6a4964f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51f400a5e1bcb605d7a13d908b1d3cb608a1abb0b1a7af6550fd9eeb3ff4e9546debc71630308b95dee3cdd065d58c1a0607523b54a5d5c60c625d5f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0e7164cfd089a78e80f27a6f1ffaa21e4f0a4f89d837dccbf72e1e3cda6c8a09381b59d0fa9462dafe692acfc777a0197a42aeab5807094055d0f6a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8044ea034b45aea583c3b0b416940a2b2896fc01a1c6235d1bf28c94e4e65bd2ff71da8ca82b3ea5339f5fc75430f6a2773f4a44800b7662045fa36a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3882983f70403ff474c28848645b6a17b780cdd7e5fedbcb8ea6b9bfc1aba92acd79395116e73b45b0d0115612b5a85ed3f2eb7b3e17ce0701f072e8a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h426569251fe4e21252584c9cab7f8265808907b9145d22c7013361d3b7dd8fc9b59b36879680baf7fcb34d33fed352d3e99411cc4b4987da33e606f4c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff2cb4464932f92e9c583e420422ffb0c2ff8797a7180851dd1ef7a7c4995a6d4ad151f3d4e22d431e4e48ae65f699468e4cb62b60ff8b1d24b6d02c2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c508a1946cbfbf5ce6828725832917c9dc65708e4ae5b72a6d1fe4dfb30918a41d827bcd47c1b4136a4e2d9184f17a2562d9778d3c264e791e8d794e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35e89fc4d032d48fb68b49bfc25f0ff2fa470b84ceae73d6b86c1df84e461c89aca10b9c20d0087a864a3028eb853f6bc03830f56b1f885460963cc0d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h581867a0a212694255c50f1ae82e1664242865f28459c5ad2ae79e6336a3135bd3d17ffb41d56bd6c362d6abcaa1a3ac1523e410b0496d6e2d8a717a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc722fe7be3a0ab6083172f311d6a4f5cadbcd63090174d9a207270cd4cb49d45593570c3a0eb28346ed0e0166295c6b71159c1f2c40e50c72bf0d01c9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h560aac3d04bdffa8a6a3e0138e44e7dc14d5c24f46dd00921b22f96dcbdfeb8da95f577503b193889f9861a60447e3c63803234e07b2bb23a8c03d0c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53d283048f252d465e4c49fefc0e56ec8f0b9a8898bd960acfffce950c92c1cb1ad5d000a8efd968fa7340642f31b80f2c0e1b89cc80c24e6a67d3747;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc14a2e9445bf589e95590e7156ec85e92908e1c5f08453d88f7f405e5f9bf1576bb1c9e367a3ecba3cfdb5cb193221e6befe09ef9a0e0e43fef3113db;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15a79d1f5e56ce3bdc8d731190bf39c3c9fceda2874205290e6c1537e0c3ab7114376463d24eb3f8866376c22ccedd1449488fe9f8beacc153e00b3e2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9088dfd1940c491a34ce96ba5de78e47ad470697e8a9c01ae86025983290d315a321275618ad6bf9e520ee989adbef1c99d8131519ffd2de72daf6ac4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf86fc8811365b467c8c23df678234aa0e27c4bc6e7b325b3177fd0c66b10b9137dc2cd82cb7362c4e39f85f53b3eb952b21fd4be07ec747c0145d8d06;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc592e4d852d6cd6c8da2a1dab20eee31cca145f9246f71518975bb70fb32247fa137b8b8a97f881fe4fff6cc58fa8e44b06044208b6d4e8f1638447ff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae9e703587e8fe5f0004178c2daba7bcb7b93ee6992c4da8ae3b4cd54d3fd3f3e30e0b1019e34c56fae646c0eaf730e6447e6de38a4f2d1abb005a759;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h286ca98ee3008adff37f770221d11076f0796599f935392480cdaf296b3cd4d312441c7dbacd2692c40b89a47fbb5a04f1aec838ac50ecc31443219e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f631ab7fa2d6c9312f12c8f1895d0bc88dea9e9e2eba0ab26983af74706697557baa9a1de19d08fd2b23f4ad22aadc390de0add8b6332588ee948522;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbee3724941ac657078536bb16c8a560b9fbdb48da127333bf928c1da8c2edfc6631700edba382a70f195185bebcdca233e1bba14dbc9ecdddf82b3c37;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4aae7f1ead7ed626998b9846c4b62746e31fab765fb081c4a2fbf431f0d72c75c6a84bc921a36d0391b556b170be9a369a887bff5335e5190f833b69a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fb531bb0b7796214fe7601fded096613e7a64eeec838c1d922125ae4b151540c1dbdaba4f54684c970734902ee4c326b72d99e834fbf2c8d97a4d45b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2a31c0eac41319ad7b49de18bba7fd5f14b109447002a209093051a5b3193b196a737c3cb4bfc36b655bdc7af73ae17cbc41afadc7171c620ca9c5a7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a36cea1674ca75746deb09726247da09240386bcf42ebede121e8c407c89bd3af54a8f644b09bb75ca6298b02e7d2b44cf639a46834150f4aae0b008;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93d38a7184f36e0e92c88d8e717e3df5999c97c4c7281aa9defe582e9625d62a624cc9fbb3dcd0c599a162078cc23010f214373026be39283fff2b267;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68f43a0b1bdbedc3e898b8c9ec21613506869b0f19509c48848dc91e2dfd94d0aacddd2e1c7b9a39bda3236848cc541a1c8307604958ffacd2860d48;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c1bc330700dab3e8e0916ce163ca11b2fc38eca7201cf32b1994b03f0f69bc1e5b64c53d545d301bd54546c163218219eefdafb83bf321ef2bfd288c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbf531353cd40bb1ee8ade0c31699284f2e2d2870a1603d359ed60c4cbfe78c5ec17d8cb0aa905ca3478fcf0b3ef780c7e532e75cd96eee312d838bbb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcebd7446d7afb2ee4ff50f02bc4197b9d5f58c11143165d85c68e71115060b607ef17a5d7f6ac5e31a4c9a7159293ec3a4a2d5ff6266c25b239423f33;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h482562d9485e62fc3d9c7e5f98643b907030fde504e24be48a3efc48e6b6eafe6df7f47cdc47ef4d631a0080e5e82ee0b0da7340cc931c9bc7ca3d7ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf057513a4a5315c5a5915d51d066e46da65854157baf081fd6a3803a3a9041d77fb4a7a210ebd4278a418ab9c0f03211e6ea5d4b68b6dede4d5a3623e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h23a16ba7f8f76c2b076207c6d7023d17be70a8a1341ee8882d8af8e20c87d160eac6024f69dcd933c30085f2556105bbdab65136cf824c458eaa89f0d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1ecb90e6df8fb8b83af716de77e9aa1a75e11d2a90a36178261529715a84b53754c2a8c18594c51d66da5059884a10e993064685d7142a9c2e90ba74;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15ae4b32f8a618debc4e88830ef9c0b60008709856589a3bce52229719fe93e8209ba64e4baca725705fe4ac3bd8336f846baa4805b8aa54cb81cf46e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had42a4c8084c66a4342bb4677a9f3b382a6cacc6b9599669d7036ebccebf20a55fcf2b184ee7f7620ec467403c1c6b6e4fd49d9241cfe3d47168cf826;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95cbfa5f6b2be1e29f9bf3735e5b187c794249047f224063e446d5b76dc67011a391e56e62fc155b6bf24880de2475f4372f26fa68616dc6ec4e6ed2d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf37ee9b1461727cb093f903b5619c6423c2853a452828ae6f29721419d75c29bd8fcb2b9585255214c29fe8c1c612ea2888e324bfe41f755f957f878f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3afaa2db79d86ab3d8e6a92a2169429de1769e326334e184281a3f36ed4a22bd6b5d3d26684ca220b018ce272d72bf388e7c8940553c551c37536b6cf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1185ed484330df8b61a2dc44aef147520b362c597628c7bd548127da513050bf0be9272540dce7014cbb82396fd97feef65683bed496062d5707f8de8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h487771314f13f8c6727a0ae95b8c2f0eac6cb964cfa7ab02b1a9938cfc75daa88b239adaa3cd8de7aa51ea6796e5e0d17b1849d8a2dca9ce6331e5ccb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h588bbfb381dd1405ef1fd7c83f5546687e308056d64c102361a32b2c15eb70b531aebb598a5774d791d638228d3362f921c3bb47fa24f5beeadf5b880;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h637db212c6d26464e9998b4ae8ebfe170caad15897def101c4f288f1dffd8c87695ba200a11ba311716a69226353084185915e3c80bf6da87794da6ff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8854d4dbe8dfaf0cdf91706294fef9fcda706e41bdd390dee816a270693ffcdb763f1e1452e17442fa0e9e387fd43218287692373525c9a2f82854e17;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h203253298e2597b050af0338edc49b859b30df7715345411d875836456cd779cee44b2a5c7f1733e0b79924860eadf53dc3ef7cbac91fb9c140cc428a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72af2e8bbd206492cf8ae6dcff6476a92096ee87a3621f0e745244139006c89ebba28ab11b71e6434d9595a8725d986bf896d59151adde9c34a16b36d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he57d98901f4a8c85738145890b737c137faa8a20acc7be4eb79f83254c4026d2ea28bb5ea49dfcac1a11e29204839d2ba8771569605bea3869942494c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30b6f8128c087729c5c2e4593c39e8d3bc8d6a698251812bcaf7f97ae1a9145a9f31dcb3a05d9594bfd36b89ff12c8b747e642b546abc287a41697170;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heed4da61ce7f13d72b9723dd4a8b74ad5a5bfe38049b338b651c290cb6ac6ec6b000ee8b9f94637e3166b45ba2b55cd007af847cc498a00c3287bfc26;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc522bcfc13ce4f45e15f3d3a585a256b778e25ea9f6772959a56118255e2d1ddc9ed7cdf22f3d6311151f73419b2489961e4f4cb2c1795212e4526c6a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf174d2a51b53e39c59fca10bb375ae6f52f20bc24cc4500f5d6ce0fe8839ac97f61a574994b9436e40349f8653e4d05b1cf0f4338b41685d01f6eb6a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9dedd39a5e202f09ad17eea2f81f906f964999efbc1a962d4af5ec46c2f981372d7c8f5ea30fbff7978c829a61ab7bf111103b2e3a5a24733ba00075c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42d792b03c4e190537769fd69c465aefec1b996075df1256b443d29607989467267d5c403936c6d1fb1d1a316fac4b94e8a9fef8df40977f05a51ab93;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e11f2748d3d7c1fd6c93fc6e7661fec555695ee35c7a46f5f703bc8eed496e62a38ff7f18cbff09e6f36cebd2e27da5ff7ac6dfb005542ecac4ed6f3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f11a7624e6c2c06cbfd1c6bc83efdc4967e111a2609292d349c537f9f3e9e8a186212e2ea2308d57214a3afd3c4e907009d35a0516f27c6fe3a0b4b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf692a2ba535f7da3e0e42670882ce6d219de6d8a778a0c2803f1221da19be7f3be4b918988e9656579348e80752d4069efa80d8d4eb3eef897706a0f3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2136792410ef9a058ebc15f3af5619d2c7436478381e53a56a14a9880f6a44b6e42de7734cfc6c1b06c621eff8aa6de149d2822835b6d993b9823366b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42da68ac8e7ca9a5c1f4841daeb90588fc0f6634417dddccb143fff294e19072f109634a6e50222e087869a50ea8ef85654fecaf24e79c856a127a1bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb096553e963488e78a7067a22fb2b055dea77a8715c600c479cfed3b049e079f8ad9329ecba88c9c54d4aeaec7c8e8a12ee62357de0413fc75e548b07;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21dd8b32a1bfb43aa7ca06e67385d849a2adee70d7ce992468d75d18bd92c6e3fb4ea6ae2ac572551705cca40b62f20603b2fd95d4343f6ca5d3cc871;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0314e6ec28bde6dcc3f893b06e2ed9df8efbfc7fbe4dc7777c9728f99080fa151c8e21af89b2c71b5b1b4ab3bf174dc9f92465034e7e16b6142bf640;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haea9aadbf0de2bf933421dcfcabeae6d2b178efd6a5c5aaa3420185a411e8c15893044b0a58787b58900bfc7347e371af7bb96f052aa4221ea4ad607a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4789e4374b3ef71e4bc30e7d8986932a1b4f142d8223660cd32a7e8313f995149e1c76d59738119ed9c2a0d79375d5167d3581e04db660aa7eac6052;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14b864f112fe3946ae0a2d39457e58491d0ea02cc46d85490f64a5f040e271b2e620c085f7216cca82342e1f83ccba908165113026a2b3c4dddd233a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e0586b3bcb6fb8c19a96b733a05659b1c03a9715a020f707b4167c41a662651a35603673e4951099c861181bda07b5e6de4ff597b7a5aa96ce3cce8f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7de2a67d65cd01a2036d0f2b893e73c2b48086d9027cf9b5488b91f35b00d1f680fa3871ffc96d18683d7ebb2188a01a1fb8a05352626c5e8612ce598;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55cb561a3f0e29bd8858af9c67d3ca9c3be49938ba5468e841a31381dc444f724e317223d485f44337b66a4a25c72edaf25bbe9dd083af57b09afe37c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9be75b0da1752b20cba757f9e7f3aa9d7ee3828285acfc2bdb4e15d25b6604c0df5049f569211e29750aa31853eb8cd2e08f8c4fd63a24493f21aa47;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd198dcb6baa0d525370aaf969282b29873991c6bb3f87774d611f8dfa0a700fef72d2a292b2fceacf2f7cc508cf9e31478a79cf53e95d5725588c291a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb890b8e218ba1f81472c7266393c6303afe7c9ac714d0bffe0a3350e466927714cdc749b388b05fc9ef2c7701c2ae5249333191b8ae7203edba053d62;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30988e46022f89a260a87b6bd7f0bf8919db7db5bab7b0d7bb45664e581a7673978492b75274bddeebc6c9d3dca50da0c8819154f75645da58e7c3286;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9a8ec43d8cc16dd8cc51a1eea4c231c97ba34f0c0a054f2ec0934c760bc2f913e7b36064dba482b4e35449bfc228ec5190c82a1636921e6aad1b1318;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb08675f4826285a45a33e5cd2295e33790a3b0fc0035d666ec9557bd965a1b130ba234fa1b5af7a6e4a0e4f9ff1dfa29f2517fc5ace4ba5968b60c2c7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0f1a3c8a4a071e86097319255f6cf35776951d948f706d8c9e044cd7434570c868db981ff397a525fee78df1fc71c433755662c4b5267230aabf971f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h927088223f5c40d10a8f958eab279dae7aca40bb74d14ce7d71cd104657dec8ccc7b61237fc5497b13cef234b8232c785c99d1dff00492aad136a864f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f02852f669b0459e701267eeb24a71cd93a6107aed9f0de11a8bd28d918c71799c6ebe9a23a3beca09d39f07c09ec0eb9795fd2f665abd4d388162c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed0670cad8e51f0432ae6a9c1c79de2a8c7fb2e5736b553bd14fbe8ccbbc5b46e7e569654addef6990cfc7aea1fc330f112188a67ed10b467ab115029;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc586eab4abc1dafe0a19c15b99a4738a2d964cd8e4cf31dc264821629bfed7947922b4d3c094155be248bcf73baab6d00cfd7a53de00d222167487be9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41a2b15ec67e81fe05aa7a8903e638598ce402ac4715405a724aafbd7be0669d6a6b860e720f6ad52f4eacd2f8cee41987dd45a5214b50d16a64fae12;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9d2e50fbe72d1d28e064886e3d9cba2136e021466e1f4cf608bfb74d043501e608c748d209a7a2b7b0a0324bbac816fa120f764c06c34975912168e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89ce7d0eff1b4da74bc055c73df1e263d1b5d31f3f83f2ac891aa801dbdf774f1bcc755a6d909f3c04e4a174ce78e8aef74a40de74b97bc6a4aaa160f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fb999faafdf06db587c011a082da533e6a003f64805b84c48e3504171927a0ca91168fb0a4fabe88e61bf2e0d1acb54fa351c701c732c25641d4c119;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9207233c492e6c26fa8bddb0d2da5ed05cf8e67a54d7ac015b61cbec128f3b16b31eb75a1ae29ac1c6debffe0f1d7b5f52c76a1db2df0fe24bf647b0b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bab0c02464d7f353cd4735f0705b42f1133a5260b3123db739d61b3a3673909b869a41ef924c06dbeead9311ba55e9a6322b40cb7509a3e8bcf4746a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8c91c3d21d5f57702c547ef555b5bdcd67dd2c6781d386b0e66f3796e2550f0178c4676a782d2196b431d5747bc3d0a93c2f942554ce8e04e6ded80d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbfdd6e556676d5bad77693e256eb011c647260f9de605320ccefe0bc73ea7c5ee463e6e68048e4cf96cc5fdd783318dc4cc93cc44190e648b667589;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36d34daf50b8b0d0599f3c370beed2bcef547caf66f2fd09f648557a7a6dda862f1c9739da5e9ae4454aa722820b311491841a20fea8844c56fe1c23c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59d64ad077292fa716ac48acbf0f659d307aef101986936bc8439e426a48f84e6941feb5d706484c0f03bd29ad40525a436fad8c8e05d5496e5b58f93;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha29cd66a6d6ab97b52463b3fb8562d0eb48d6822f20ff9f00748d99920b32ea1947584e910cfb993b04bd57fe3b0297b2afcbb38bbd7446dcf93d66c8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b95c4bf7120d7181f5c1586f90a91054fbf78a754c8c5b6bf2f2dbe7bf00b5b8395d0ee381aaa9d56cb9b5d3d2f346dd25aac448a07c052ca136192d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd59b32da0dc01e7e536df391b4b9dff5350a8ed07e10b182ef9846c7ed2f538c226e02904020221a1ac6afc98166f070def34f4b683e190f67f0b9363;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50f6e90bb5a8901b548dc116e8ec546825fadad7d14d9ee5329fd133aa469ffb9f18f0e51cc8663b86c2ada4d71065b8a811bcd1fad9840c7a8979189;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4605a85db05520ba92104a7d3908f313e445576b1d1c14d11e7c798d8dd6dcfac2e012428572c89cf09fae574abdf8c7376cd2fd45f426a4a8aa360c5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67e76d7f3bd69694b53bbdf66af89fae197a3405c527f4b16ffae0fada8235fc1048c38d2765265c9b8418770d916522592f50feb3b3b91d50b0c33b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6f818cb1e855e6500271fa80029431edb7fd86351463680caf11acc23a92ce711e0144e8f4ff687f36b5cf7056287091e8d6fb5884e35ee68f182a6b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he437c00c30d8d7ea4999e144e8295090d3489ae762f6dd4079fbab52c35c88c422798955c62f216c6053eef6926db5c02c0c52c88be265e2373196a50;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5bc80c263e5358e77695d3031995d2d7d5b7fcca491c0cfdf1da43b709417d1855682f06582750998b5958da6c910e52eb07f14da2154081d652725b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8664e4d476d06c79a63a8dc8d34ac2169675cd0a1df7f5070b014540f7954f6891bf4123f20b6c798700236513dad14cd4ebba129948c5912f8a5563;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0e781153dfe804538a70fdb080a83543c647d6fbfd53b498d2333acbd80afaba82f5df723f877d2b028dfac66d55c6c62b5eabd806490d6be71e8a9f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h595b4280c545a5d8ea6c3bc78e4775aebd3be76b440fb48a8c08ef2bc64dcaae02329f646f9a7032fdd70065ac7dfa96e045d00be2652c84d2e365c32;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hddde65ab7ddcaa924ebec13b5f9781cabeb84674d0026d6d87d5efb59ed68e5f4779e5c9bf87c7f9573274f7f1fa0afbba5e32d00fbfdc80b8b019a38;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e63eab2715c1fd285e826ba91a9fa12fc378a0c391d4f1d2f11238584e48b70062bdfa4fa0702483af2f7ea7cff69891855b7d567fb9d3c00ee7f278;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6837c42119fb6be323bf1fc32f2467aa9036d30628c8c9a26e72c836754f640f7b28c140a58c5e26fd203e0c3ecba45e771ddf5f1ae603b3999acb04;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b60a1131cf410ed722f988071ed0ca664628612f9975ae7816541e1907d33f98ca5074b12d11b9ab25ccf86a80ff8d1bfd84ee918890fc1496d658b6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3748e8e96a87c4b44a3339f35fda7181b1d3e39c286f7262a5a2c1c91e66eff8c07d513fe1fab668ebafecbbfc936345feb4da15cb882d72248be0e9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d641249504cb7594448ab4879b6d6cac1a8f8a57ff52331fb613a6f93a44e2c833324eb148896d45bf92b617e8431d43584226ee45bbbe9e7afcfb46;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc81e149fbf1b20080ab69b7ab488370b5c6ac74f7b70a16c69b408a330c3e244fc2285fc4dd8ba1be09b799a22fbf68f3ece79ae9bc5a57dd09a3f6c1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91d9320da8874c588d7c43ce5151beacb21845213a9d9470bdd71a9656cf7bb7023387c57975904f1a0a8bcebcfbee0bdf547ecac62230494d940d402;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcd2777f7d3040eb322f4c83025163c2a16a0762f934600739e8e9632d6f08d9932cf11f022ccfca9ae119d7c179853010964561721114f8cc7863306;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h988d9367cb9009b08d18b84e498b66de64c852a7ed7db23dbdeda3c8d81cad2581c6c6ffeb8b4759cfd95ab3a5e75169db06c4141f4c4a9f32b80ea91;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0127712f0fe008390c60b062366bb0695b88f81e930e72c9e77b623aa6ec3f27174129e96d1406e44910a6c9f76ca3fa56a8b51ea16c0fac738f59f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac09a18593335d167b3f1f96bc1e8ccf4258c43d2ec3b0d931a2f24a93d0142c04978628ef7cd8003702b49e11cd99c0f9037abc097221b84a79d933c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h433af7c99b9c099211834bc09247059f61de6b4a495af29a826a10b52edf7c01c690426b70dfcdaacb30362dd90ff7a6bac6b85da49fa24254beb9be1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd12cbb98ba165282851824e347755d7cfefb15efc85d38c4ab1eeaea6beba7dfb5237f6625f9b9dd031bacd22c774c1dfe68f47d4403087d45fbc156;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2cdfde883129a517e755706b45a03f52b48c8709cfbcb4bf60f86392d00eb0ec41e26a982aea4315da3bdb59cba2a98e6146c3f1ab226d893d71e25a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3b9667b9a2229660ad0d8b3c7f8588e6832b3f520983615fce69a62fcad332af3d1b13fdfb45c4b8c6a52acd94e3e3ad3210e7f30d445c530369cf10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fb0998607fb97ca110c4fcadddef0f3616417bbcc9987b3b020fd0a299abbeba0d3e8a4a140a2a025c33ae509968b96379dde16615be5c0c452ecadc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h231da5d0bd05b1d78e72ba3080feef3ea9db4d4f9a9524257125460a31fa41b0f4fd7c1844cffeedd490c291be91585c3eabb956c1a7a4e59b25b41ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7739af62bc9ca7fc8f8dbb9879c7aecb61971c1cd4909c6d2bd448a6b99bfbc887957ff9736681a0563d7fa99748b255fdb01ffe568c5c08ff2a65d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h686e7d09844aed632aecd1e98bd50d88c6d5a00074c48ce9bb2dad562bb0ddb67926557478b8837e7853fd42ac7bb7b1978191b9b1f36ee3924e02c24;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd24b462f1b38ed1d4014fd1b29b854a67c4f0f83cd22b7fccb78cb319bcbed699972715962a9f2d7ef251e22cd854015c24451bf9b3b957c59b6128dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50da1da8cb5f6243c16c7985633088ef355f842277e188794a8e03f483100ac78d64fa45289773432df411b3ab5d3e79fbfefb0df26afa727b7e4fde6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90812164156b68a68ac1db1e5e641733b147d2070877ae794387eecccec5eba4c8a18b45ff63e76c2ce750271a02f97b7e936ff5422ac12e67f73fc55;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3227fbf00b3eb2d3f6c67b26c0faf7e21a7fb271ea1ef7e7d90638b44e5798b6367e54655c5a9f7c4ec5e269ead0a1ba0b13e4ab6566b9b1af18624ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31e4519040f709432111cdec9d8cbfd8164cdcc511eee75c4e3410175af852a4379f31660475e27f106b19ebc9fbe390815e74482104a48b1f76128c8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h905b2409726844ddae22b469313b47271f5079017bb4aba9177370a8d14254aa780140fe4b5436843c1dcaab1b7f80fb0f5d1b22efc02a419b19e3807;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h185fc6c3fed6d23d445b4c5856bf65641d56f1e6a0d2a3e3d23c8cd4e7b848483c817229b6cab7fa0d23d4f03cf8745c5b11cfd1bc43b3015fe571dd0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21867a8dd0a3821306c6318d3f1b592395a19f08ffc459fe5792c100fd16b9cd452e3373b8dc0a7a2e3f18d0181618a793854471dfcec8bf920e95398;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70e6b91684b6a67b3c60fb065ac69df1c32e86a69ac62ad5756e70a6f0f72f98ba26b40408f84f20533913541a5abbb74ef34c8845eb5bee81f81e963;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fc7543eb7fda0da96bd2153911b56432325ef7cd5cd3ce17c20011b2d574977a0da8ad1656bbeb90b1db782a6027ba8f1008ca222ed44c3286fe0325;
        #1
        $finish();
    end
endmodule
