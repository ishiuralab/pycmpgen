module testbench();
    reg [23:0] src0;
    reg [23:0] src1;
    reg [23:0] src2;
    reg [23:0] src3;
    reg [23:0] src4;
    reg [23:0] src5;
    reg [23:0] src6;
    reg [23:0] src7;
    reg [23:0] src8;
    reg [23:0] src9;
    reg [23:0] src10;
    reg [23:0] src11;
    reg [23:0] src12;
    reg [23:0] src13;
    reg [23:0] src14;
    reg [23:0] src15;
    reg [23:0] src16;
    reg [23:0] src17;
    reg [23:0] src18;
    reg [23:0] src19;
    reg [23:0] src20;
    reg [23:0] src21;
    reg [23:0] src22;
    reg [23:0] src23;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [28:0] srcsum;
    wire [28:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haeccc0639a1795fbf161a162c157d45c5bdd71b9959333dd280889c7c310e9dc18870794cd9ef4362143d5d207cb6701b9b5a6a264ff738c8906a22de6d39d189e9d838c3587d7ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf2ebf2beaa3f3fc0ffa3d62895cad3398ba3ffe2cd48c6a62459f2f7a54cf60dd77280a696b69175c0dfa497def7d68685f194a16b10b3c3a26238d566cbf4fce50ce319c14a09e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97a34bed9d00f270295ee081c6b519851ec2fd511183d6bea80f225955cadbaa06928593856fb57f33c10455bceb56077615466bd9091bca435e8531e0691c60d2af4facfedf16ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9491ea4c74a1a68f179e637924ae10b653cb00d84e3ec864811ceda20669a5e56241057926c4ab3cbd6e5fd32c789d5b08e70cc1797ad9d19fa3f6348219f2fec2de2404be19880;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9562edc8fd1799984719de48fc004d2bf47b49e16c2d3db7cdc93bb4b1be57caedb7529e8c7221f9c5e2c646901641bc7ea231453aeee3d46cee11209ac6a850ceeee638ae9f7ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h844819c02d939c0050d313577dcfa35b89e5b2c97a99b08a4405cc2d044cb226c0e407a8c00d90485b50ccd566bcbba69fd20f42e69d7198118986e8aacdf4a0303eb827283ea4cf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h348f276b2a74dd59e9381c2220e76416dbe9a5a740ba3850f2dcb4af4c16fc0a11b38dcb00076776d858cd660d4af33f6a48047cd46536f68381a974456a9508540b2bc9b3130712;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c6aa2fa51692d221b572fc85285959cfd997c4fcfe9d7ce54957b2815ee0fcd85ccb7d610b1975dc8e1f4ea39815eb74a1e1ab543f5f4ddc0877d2f03241a8df931e50b6258d99f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2c72f0531d989ac97aef9b84878faf0fb13698395e42c71407a0b4a372153f850e81b5dc388ce3f71c5829e31fe2a22a3dc5bd0aab9cd79140e7ed47764010514165f6bed2fd5a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4d1967400cc847e7e1f9343b29bec14c20ddb4c4bd938b8eb0c7e77d7471b05de4a0d21bc3f784885163cca6901b70ca12d3259bbbfa6ba094143d0147ee874ce93c34c3ef593ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3d0cd5f806fe89473e593dc19525cb88b400f2cca8a745dd2e3b78728e3d1064bcce8ffa6dcee4a062f7af96f3782e80b247cc3c756f379cb0626f8e8d8c08ef9b08ba9ee10b87a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75d5588d6ead0f6c3c32539b867f58a6d8f1f4a669f584308e4befbc61dd5d6b640bf4eb4b0d69b409a2fedf8fd6befcb00a460327070efca6eb5abda9ece08db2df12ea7219b72f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf34b54dfdef0f5daceeb16ac1242a2ad0cfc242dae72a37a3d0f399d2a16695e7896cb51f0e924a4cd64e954945e96ed30ad329138590b1f184ca9c1d6ee11235b2e8a0753fcbed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb4c6881b26cd1028437f0f675a51be08a5b7e8968b96af052f1ea4e7c97f492393e9af5709957984e4b38c1cd6bab5b0f396db375639075115c48acdaa4d81b55a9b3f1be108350;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0549acc4980153c8169e076df830e353a454f8851111af0140647cd2524cfa7bd525f83573fe88d7d7f4448c2fe6959ae3126a850500e5d81b89ec8e997c6c701fc08f0e7fed9cd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ae4eab13c479014551abc4e8bc6a8b7fbf7754bd8fb30ec387d4c95fe3f2b346f0edaad2ab6b414a2b8a2a9be92535677b1949a85994d21ad96cb3c7f0416aefbdbdb026056874c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb16b61b7a43f960aa39cf9f3df0adafbfdd39529b16844204e765e7b9eddf03cad2f3f5ec27f99a1cda19ba3de256a3e1d8b031ad8e927adc6ccc8802770668d16a7f0e8122e3b60;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4eb611044ba25f8a62cd0f65db04be806779a045b3b9e183ccbee1912616941f36c2a46e8f6d84e18ec9d99449f0e36eb17a0e8ed4522149a18fa3824da390e0705436ddb64b22d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb75a83c29b3142df98bceaeef9b4b3bc9d72277cd7293eec3f9e3dde9815a6d94117d56c36be1c2d4f9338c942909f168c8ac1a6a832d7e0ad8464de63c84b745c06980d7f851873;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6068d7196f3a53e58e30e2ee7ef0baf8290b554fa06145198b995af519f91e9ef0cf260e3a48b5ec8799c1a9008b0ffd0bf8d5617171558f84492f64e25de7cbd0fc0401ba2b5438;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h412b00d76b582f96533bd2885a3ee72f68acabe977e15981e833f628b8320227031b108dc023e76e1a02c8c397616e736a3b13320710be1fd4103d7a9d6fd447f27dcda77c33c956;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd648008c9a94904192395be0f01b6e40340b7ae4419fc963ce42ce33193092d2fdd9cf9564f6d30c8310eca21da3b9b5c95bc465eb58860c918cd02dee6f7fcf478df41edfd25bdf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd73f9ca9c3aad0e448003efd9194571ff26b982d4c7eee645fb058472a53a28b1490ebe3d6d0fbf10569f4cf0079d6a00d4a8f52072e9e024e7652ac6c843f39d9fa7d13468ecc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfe557b9292e0332c08f69577960e9993bd66c32583c86a076a9fe868572631b0c3cb6ad280545eca38e336983e92b3b3e635702d97fad6d1b12aa6294ea34c3bd05cc9cf39b6d6db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc0c3760c3369d9b235980e9cbd63cff9f77624eef10b7ffb7051f679664e34fb8faece3fe5d502899ffd72f76faf7081732231f18fd80a6ee501de2b0ab96ee2855dce7f02c78ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29819c8b27f3c46dfd055bf2bdcbbc924c23a717cb8f4d2b6d5b0041acf1afa45513d28b4887868c1ce9390eb60a657c0aea5e36720ec03a2a7ee962591f264d54399bbda5957c72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd6449fff25795beb8791f3ab9a896558f41aed188b61afd87a69f9085b0eac25099d96467e485e114349214809a69b66b3c19c68accdf882876af4d877eea63e82d5089c38c43f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha07ae4adf64ee490467ae7af722a6db60004be89b14753faa98630e078314ab42b4fdc8815d541c2f8b41738f055a6a2cccf0aaad839ff77c4c24b6e0bd204574b0c496222d71c97;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3563db7515d20cad90455bb2b4ff1dfe758c0059c05b18a81f1ade5a4c978f9b2ae18fa81b03ce60208a219371c718d3f8167e315b027ec8ba51871237143e1220318c1d793f346c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb87082a3fd9e4f4d083a9bc4ca4d9faa04ca6a7fc58027dee854a1ea4b56853df79125d256b9d1dc076bfe1674ba80b4568e9896d2f1675c9540c6ab5718b4e782ff58689afa4df6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h980be9d920cd5df055d46d99d19328f1311249e848cfa8cf7ac3964e75f9b4d7e9e10c5692e7d53dbd16fc3f27824393451bc660ece7bd26823fa31097d2735c9f2e31b20888a8d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h252e0e36295993395df1131123dc92736ed5d390f61d9bdf5f2e5082f3cdaf491929e01073b9d84525a22cd1a2290bfc3a9f2573c35225d4b0b32239723b6f298c75a72ea77ea97e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc81416dac5034bb8c3c8adee7fd93f5a8ab4138f8fd730b331d74768ac7b1dd88118530d25c97fe965724bee7c8dd1b5fa6ad92d959976e887518c159a17f00d16c30837686434e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e6f4a6df633c5c72c565e5a960770ed43d168dc20981dd66f5c9a170c366deca1c3e4c5ceb07a018dd0f6555e6114c0b77c434e4b82612dd42e08e132d99fa8d7db163db8b04ae3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ecacc956815f1a30b3b9d4879bb211a9e189af05b768b9f0e7e1da4f396c77afd1d5eaa6a9b912fd52cd405aaf743677f4f13947f8301ecef3a65da5a98617c28c5ad89d6328843;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he71ed87f26816e4901cb1550808a9b09834d235373b791324b7ac2c732dc7499ddc609301b2a1864168b12b74c6974f5f32f5fe5ad22bcd095e113f5f45f5e2de47cff67b15dec49;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c3d7194eda3c0129f1f1ce478faa865d917d2826eb6495018569e2a802bf052fa34b2ef809efe5ca79be44386bac0ad252e329f141d6c13561bd0fdded911d2a929f5fd1fd8fd1c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had3679f291d3cb443173328c12afc808182dacc78e6e0fbfdc679e223236bf4ab82bdc467af2b778cb5f94f6f93e9e27e3a9a52579d9d1478e6e2a6674947335520fa4c08ff6df3f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd361f2921171f3411927413e8601944d1d5f00903ec5ec304374438a2d8166800ebd938f1d88b60090a48332f29cfb1e382dcba6c338547823171431e2fe3e34ca01eb96026a8e5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83df517865340da3e1eb3c8ec66a6b753d2c8c40a03b7cc811f6eb7f7c4611f0a6bfb7ffc98d54c6630d272352e79225f19cf1af99c2a25553bcff16e6ba0785de3ce5c8d4d267a5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83c4ceea8272b7ed7595331db3900749973a67a06edbfd1476c88e74667191ded69f46cfcd6b778a9fcb519db69612ab9381fa05a7dcf6861968d4c763e3c01f521e4b3d76d410e4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb06aa88bed808759021e0ab8c8e9f7b4333022f86bb78373a7b985aca313ffa8724781f0115db65c372881d69720b80d302de0eed01aeecc828c2ec291c5ed1800c4f04b1c78017f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8a39799a229f8265589f61a2cc963f8ad3a7a70e4eb3abff0d8b0934f42fe94f0511f85a7ceef7ecf1743d5b3e6b667375b89391cfe798d6f290e0ccd2276030798d54a838c4dfe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e8e89450bd6720a0b13f0613ba8d6445b926f99670a4aeec7ef4b352e3a86fe57c3fa8a098b50b5f6202ae8a717dd0f95aa1144f92c9135bc5e355eaaf2b6e0d9c978526bf83dcb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb515b8a0bc89774222c8df755caa3809685a8a6cdf65a4a3027ff414dfedeb61f2381ec74573fb21afac7b2d795b81a7d98938a48c779d4bc18103f00fbdd2454ef50c8bfb60cebe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc30285efb5dc9e48d464f7b769533a149f4d752d22974b993e669b4f1b312223ac019284dfd1b05c44e784dcc4033046fc5190f177aa7ec77c36347728031a55b06d54f3fa658ffc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14039f3d3e41bcbbd013610b0393151846d08688f83aa45736a91deb3ce0c996e847187937010c1aa19f919c466c844e3f2efb71d68156d6b470b98282ed030b3d6c4a91c7575066;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c30243ad209a416a0d282368384106686560c31884a32b05c1dd81efc34c35dbedcdec72ff8d82dcf58639da4678001d7b0cbe26fbbf1802d72c3f0d56c3810eec5c1b7de003630;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb5510b814b609c3df70700b4a4b853919f0d2ece34a2a1e8276419d140fc4ec85402605cd9e6d71b0d0e40b9244455b68e750b0c08fd661df9e982620a0b44e9b93da692e419dc7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50b2f55ba94603498ce94a7a85249482bea8d67ad1fc94cf1d0718529f484e8730fc2233afeb0edcf737646620d6df6a76bf40dd482993b28190c4b876b54fe5c8086b6396d07745;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9854b7156e71c5fcd8ad91d4042a0d0b678e6d1bc0c1adeb58014ee2874a5ec1a2b071fce6b6b98d3f78f9b37529972372986d22c8a70e19be3653ef01821543caaa44e981e09c72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h861f30bbb529f7338fa787a16cd8adc7f71f43a1bfeda0d451c449b0773b219b6e8faa19042a109273e5396f5eb8a72c4f6ac493c6dc8899f8e150a61297812bffe545458670cc35;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8840a679c2828aa5c169de02ca5845f799a50d32022aa18274b20234e3571364d02b0e9605abfdcdec2e4bd05b1e4513921be33a463b9db5d69ad0f7e59faef9fa9cdb30624fa436;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21bc0f5ff9c8aa6a76f2219460164b9fa6978698dc24c48d1f0beac3fa758b8e2a57f23592fb93557c3eecbd3e437c85752055077bb2614028ff4878405b079f9f4854cd13ab1e28;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b28d170dbeea0dece778a3991c3db7a62b864f08ed831d2194eb1bbb7b007aa7dde97e28c774b77cdfa5a14e50a557ee23815f86dd960d39b669ce22842d1b2b3fb86a15592b680;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h802c72242f1560eb7eed393f4076a4d22b0a96d65c1c2d5c155078792343a98897c9a3bce60e8a5bc8360eaae3c346300981eccc1039d51d04d5aaab654e7c4b87b86f0cd4f47995;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a7fc6c5edfebd822b3c6489aed307a616641f5ca9ed6b79f90776f300fe6b1c5977e0ee337ff6bd1e7acb55694e32ace457f53a95179a9a59db4efd6227c0230dcf99905d65cb75;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h480ae3d5031cdf77f9f82ddbd54cb7dc497baeb2a1fac7d72a8e06992ca805879cb39760c19ee5cc3e70ed14e4ff1a6fdd3ec32000a94ad79de1569c81b6f42f63e34351ec00da17;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce6a66b951520b8d42f51235360d61ff395b66c4a0c4a6f96d9bd60c09f5e946c04e251f6b5cadf7d9fa02bb38a1e2ddcba972951b141f242592c4296917cad8f3b441c7f69c3a11;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h397112e1a313d301004cd09a19f711b3550bd6e4802609a7b38a3cff83b7067e690d2faf4ae8f678f066983b49d837cb168f972e24b183e0a8e649576f3d6e0524a2d59fcbfd5e13;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf10dcbc9c997170c3a36f11ba2856034cbebb2b3f29142157201fbe5805a3dbdf75e946534c09c9d556c770c1b61ec4fae8c10999cb5d98cc85287c1ac9b92d33d364ae530894e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1fb0a07f74e3c682a9ba7826c4266943d59fc4092c99f78d2fffacfedd972b37750ae82a5acaae059239e95015dc3248a5f6c8b3236def0f6cfb387fcad247ecc278355f44ccbe13;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24404f808c428b303229e6484303f9e2975e399c4e15a8a7c1dc6e4fa19a94cb9d35f741801ccd6ceb9cc21e3a24da99d2d047608ec9dcb241add3cf4a44ed50e8a0235f3746b85e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a39eecda039ac42d6cce90dfb07618b920ae9b1bc5a9e39939c7dd8b5c5083980ab5c23177fb31cd197a8ea139e3ffe4f9cbc6af4828d10a1f2b6c2dec058f2c4d29dcc0a716c77;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b9711051cc69fc1acf74a98fd3762c90cc057a1c9521f1579433a0595bb7af40d9171eb6162e77acfd5ed04c1074631ffff1d4217e2ca704fa7978e76797ce30882e4acd8a594f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17bcd560171a62ea59b43440ba54ee83f024a477c133f7eb7a1ca75d1bdcce66269239a22108e2ebd54d1ad4fe409fbc1f7378c597851beefd66c94f0c104e90655524a2c4aa226e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c839dc4f77b947e30f9aa7669e9ab777f922a686701845f8fc0c14020d7cd182087a227997be32700ae45be76eb79051ae68fbb3c6a2d0d70a92cebd87f291c0e419b473d4a1330;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc57bce550b26d17aa71afa3388c81df1b8e2851217d7946449a47c272e488dc69e39a3367b0be69ed4b1ba45115435847f24d74287783164f30139784f7d98a93d45c50d9ce8dab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9469397c31f0642c850e471b88a2fc98696154eed54d02e5006211cc453496ce8665581111b4e67e57640c7f96848a368f563cca223134c565ca8e1770b2312e5b64a2778e2401e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7c12fdac525bfba113d790f6c6fdb121c8d9df7d4b829613f297cc1db63fd96620e4e31d4b9323981a7e80aa9951d80e29a62ab40aa062222054ffaac69182c54dd6191d8d78fda;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef191d5e1e216e6415de2b6ff86e5884388bbe407e8ffa77c414613823c44419689ae8768f4952572094e61a8be3d66f8cfb83b594b564062c487b32e9b4166b9b8a56eb937f0002;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5e1b2c6203cea5c741246051231e0c3f88e09fc454d5a3b15df6dd4d410b7815e40e46d336a075c799e927bc207afae01fc61344bc3397b966741b63a0ec17810ef78eee8c99548;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48c1b109c7a7d66d6cbeab114f4138f641f0af764a328314679eb2ac43e1288c841a515e591ffba675c3a4acd1070074031f17963708b143af2e5fa9c856e84e840d44089fd26061;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb54c7fb46c1f79c1746c3f0de267cbbef6f1f6c5d5687c94878b5f518ce482790b5326940e32b90e393b55f21dab9b670049dce3297fa18788812c9a4c1caa654c68578eebaa48e0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha220c530c97fbf99d14a650fb144d3273111becf8e8e59632e63460b6da28ceb1d8d27d3277f9765663c6567f4f1bcd31e0bddf53ad9366df52789c2742c754e7aff9e70834ba099;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24fdef349282db1ef3d7720404f5c56b9f3bd6231a60173bedead4dff786dc639e7af0f2ef3758372cdc84f9d385749a24651c2cf9d781c9954545fc15454b95a736006515062e81;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1eb3eaaa510691856885c8df702bd15bfeb674191d03b4fa1ac576be9264e16a3f75710a00f5cdf9e7579784dc74027d821b1d37cae4b027168d15cc112c648aeb5d806faf7636a3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8047466a6f724e01ac06b0fa6c700d6509fced65146068d1aab95182c923b48ab99ba602950faad77bb904933ac7cfcdba2428f05a43f4d19aef69a556ece24db66d96c1b8fd8a3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a0a706d777ae0d45c7799e010c902a3c73210cfd28c5c66a28586b2e2749ea6de325af8260ba1ffa300eb42811d7d572bed21acf9d1c30d2ec3fcb92443c73111e59b71bd07b4f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda5cfdda0a853030a45510c8fc9b28c2201cf9ae3dbd1bf77f83b903f5918351f8f8e184d9b1d3866d6cf9fd54c38d45a4997e5db55abdb345a3664360f14af7e0c8e06477508eab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha74550fbd3d5ba80c9a655721dd6d7d7936c2d1be36c2942e5f84d3d306cfea9db13201f485410cbc9a0ec5b7a5fd30b7dc1641cacdfdb48f678235aca1c8158110f175468f3d14f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb98d5acef52ad40c0f0e066fded00f5014350d8b4b7b05645dd3416ff653bfc541697c98f221af918d4b1a820a0fb5267d48263a0748ecb4072dca288630323f3fe12eea3b135c86;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4d1bba050d420981469966fac5b6d7e7ba4ba3f8caa1208455f4ff2fa0dfe4edb8677e4f93dea8bcaadd7027ea7d1f045f43d9e241a9cea8e217715c813ae344c847d656bc41e8e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haff6751a12223a1c447e1f95552fbf1a13e178febbf560e3a82edd588954065057070a1a09e0a7f555021a7f4c174ece63e35827cdbb9a1dcff5b869a28cd5b5c20cd317ae8cdf6f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbddb6c27e096725712935e169a857ac78649b6c7e6dbdf6463076e10c6370223bf7459e25c0f43f246c770bdd5f74ce5537a7cc8ec495904cd29f68922dcdc2c0e16148b09cd3a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha66487416c0f2c411b5d2d19591ab04b317098c38608ab2eb50390c37df2b630bba3255d952369023b2b390893f8da2b9eada759107362f971f48fa2bfb6c49b1aa206da8430bfb5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h311f2bfca6b24b269cddc654993025675026e8b2fb1c85c6fe8d05140320f6ee31dfa8f93769bc9a1c0a05f807b76253741fc692b2ea8abdcc13437939dc0b0b26072718b34f5f39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35643a7baf5b7348072db66d47a1108a2b6ad98ccc81296c2528344139627e716a94e8df09632303245ac4431821725e88b2c17b0afe173fda009ba9652611a714f17f01dd6ce065;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1db047e93d8ddd6351df113f3af8e9a18df191dbbe5feba1f4053f94bfa5b86caec919b17f465ba946c4c3783dff1a71dcae979ffccb6895e5f293dc15c33176fd36895e93822aeb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h131377973d28ef0fbc994d42391ed6331ce048caefd8a3d0c2f06ac67b355e783cf1c3424edd82c164343685334a7500eca57d7b7d91970604b77a0c03dd6d43a08e7bf572eae8ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc95f9623d6c8b06c38d1031c68ba6b33f507c6f5cf69d087b618493b1db485db2497d6ed719ca4e7a908dbe3b85a4a85ab3ec8baf77e6ac5c4fbd87593a01266989790b4f09dd92a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf095f6dd1c0be63e9f6b9d9b7e95780c668884606e73ea223446e246942948a560432f7168bca076549b69223379d7792fdad6ef42d9a3d314503b156b462eecc56f631b241b3edd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h137e0a035f168010541e96c241c2d278ef09685959527a01abc88cdb4f6d9605ac1e6b256dcb2d1ffee38fcf0bb0d9a08b62ac45ce92e8931ccf28d2680a5a9f9c60c70d05d81f96;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e88be43087858d19eda332b8cb145b1185e314a8b477490ea9ead2b3e5872f14f6dc6489a052dc449a8735ced0c72191bbbad28829bea8d7fde724a9165e93b95d1bdcb2cbb457a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf42f6ff859455da7116a3924109234fe3abf15111f99b69acfa1744a5ffd08cf3aa2a7046971e546a9ace9392443cf44b74c3094a04cfdd07ac20d44f5a6dc3ef3cce4e6cffbc16e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5f63f775fcae8933f4ccf969c7316cbdc4957b40194bdae45a8bd4c7ad498d56b572ca5ec301792147d229e3cdf9eaa51063dae1369a2131a49cbb22117a26e6a2ed0c497fe29e7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8336843f731ebbedda56d303e815c603f2cdb9e6a2747c91bec7ea31b5b6bd102459d649a1037a577c65c2a6883d1bb6f23a832b1e48e58da3494954c0570d4c57f7262ade19e55a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d4dcd3b495ddad110fa9fd04908a692546e413dde9bb6aafdab2dfe7fb0448cf1c691df838e93721cda16a93f4fb87cf744dbd788dd2750c1eed4d9469b6fc5356a2d07a2514470;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd88ae017dbd9f58679938528d9e5406792a66f7b0876f388f6269e3b05ffa46c9392f4014aaaae5703370f9718507c9f3970871c600620d319c6243603e1414e3cf5c957651ffe8e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7dac997d3fbfd5659924dd39ca9321017023bb3a80388a5b384291ffd0fd8408004e4de07d10b1d23704cd3538579d79dfa9a8a46ebcef55696488a1b49f64a984f2ee6a7f6a031e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb90b04bad9f9a9b0f95d15cf6acbe887e512752bbe2ea854c517cad854915506db3f24356311119b94be95189ac766cda05f7bf0124f972de333b818aef34aa6c1347db0b7672492;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf53a40aa0d38fe2fb275ec03ce11d0d6ea32c1694a5d2ca949856c6df489f0822106e122113291c9bb225ec66064e7ae8b37502c19e7833828d5df709b93826f19db524932f3e5c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7d68472763a9e0ebd4c597fb41ce8e80f99dd7af5968874418a3d06b57b1080b9ef16b8fbc4db81df8d49eb12ffede3708ce52c02b947dfea45066f55b8782e97c77bfcee46a45b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h552bc14fa3ec8b35f1f9c7acce4d9f1d020082e340c87e5e01c173f0538ae71efd1bdba56f6b14fb1ae26f090561238513bdbd24242a29c3068b6e9a7280d36e52080a07b041a434;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8e380a91f16b416aaccc43e2a359f400501233d5b100c6dc53da83beea5c4957cc8df81ff9f3afe4a4aca649e24471f0dbd405632387c95795c539fe7d7aee941b6e9042f862921;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2165078afaffcf8d640a9d0be6fb35dfb14bceee211bb23d24b9836582c70d1fc8037fab997003d4df8977a5e1f8f79151ba748f60af9ceac50b630668b39939c6c9ee818cdebecb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0554daa91283bf01831822d3f068f6b03624d7f408de5595340f13f2fb1019b404d43af2f0f16d5e44acc89ab1e9df0459b2d0bbaaa16fc35b6823ad46c3332b2c74152b4b02a50;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61a2a23ef54e9a0b2a6953f91497d7f0d7f6a0004ff6e8498260edd7f5d27aaa912a7d1f56921138c3d6e026e235e82ddb61c0092ccc70102ba138b13529301938b49681603dbd99;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34029f5ce4f59bd1b5c0969e0adeb587ade15126f28d1abb23f7343358ba397f09b255c55fcf53181a014a713f27e116f4d35e8c45232fb82dbdf1b77a48ca41f8e353b3db7798bf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h308a195fd136b50294ad64dc747a69fbfb014b3233b83313e4586f5350b39c381d94caf875ef6cc76930c24fc21a736901d8c15b64ddc9902d6341da6864d1327d540f1e455daf20;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d2553be41e3e08b592486ee276b7f89426abe085c47409b33d67e317f776178a8d2d2e0311291eb5240bba37d47f1fa8659f4904f41be0a0bf5f845f4beb202fd08a881a08692b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3c4f4608f56cd642f37ae99fbf6e798e3745fb1bdacb7a4b38c9468e14a0cb95972b1ddffc3e31badbd31eb9c26344205f7ec0b47a75c3505664f5349aa0350284b9d6b2f557c11;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb614bc71a9fba07f0ea3d72b26d12d7c4dfa27ae59b53b26ab4dd8b6ff09c130bcbdb79c55ee778cd380ea6665cf59f56881163ce984d96d234923ba64c9415720c6f9ac1dca68f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1ebd217c76953b8eba9dd3cee04f1e4416dc2c5e82d650e1b22afcb000fad03711e2d37cec58f97da570a39b1a1669d845566dc0a3af2ad0da686aaa310905fe3f06901943f9a72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h167a9987b0a35af4c9722884fc33cec624b85b6b13156c2c7872f0c38c996176e74c774495855bb3be95d1ff2a73479b0a7c9c96c89f8f4527b72fe565616cb54a1b62b4788b3799;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51755c37ab96f4db5812b9e3e2f5ff2a11913d96f2f9a74f597dfc743caf0f57d8ad8648d134c5f546015c64f5dd323a76632d6d158e6c7e80bc1fc772a45456f13b9f8cd05c94dc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he91d9d285ee450f776985aa928cb6f77cbd7a9aabf10c7007586987f50a1ccfcea6dbe9697c557d3512642da76944de4723d9b34a33c7e81e9638f66ae32f21b3a21fd05535841ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9043b49b3d181bd7c3b71e2201dcb314af1001644b82456d3a56110e019951f148b44c03ee45e19925ee65c0ff50e4bd45fcc81196a55fd1553374affecb087d616258fbaacb2a0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97155491b9e6ec8153551e1b466766cdaa18ebfd13b8c6c349a4c19ecc9e7f6625ac09aed51756279d9ad0015af0f29edc3dc3364889fd509ebe654b1edd73fef01c17f27f980e6e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2c54259ee3d226222d7082a64f3f1bb37b192f4be92d5780494c563d1f9a35676b6181b61c9ce9c92730f92db9597c66e9c758599dfb01de7cb0524b380291838295caae7318abe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81a79880716856095cf56935cec80bf61e166a05d2e271b00a4c9598f06df53af0e1e6db4a2965d7b4c2a11653c1b0cb733fb52b36ae0a2908fbd7874dd2de2bb0074e580a56c9c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a0934858947ab995571bde7a76ccbeac37b62910c3bc767165b4b8702adc024dd25c1d1097bbefe1191e9bb2aff11136cad01b31e5bd4f10dc271e976a3633748f3ec3bffefefcb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca57652ce2c4a06967a8429f1ffa048c741a4151b97a26754d8c39cc532da0a0ca9d1b71e0b2f9a1832fec4bb58695e387afad4541d900f7332e58c4abf2ad81f7b37af24cbc3646;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7150d7bd0bd8b72cc2fb733b2fdd8605d8dc694e3aa35a9649d01ac7330642b55988587f3109b9a86807dad9610d8a1f8ef96442426e6d70e1b5ed516d07b3a10068508c210243ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b169236baec32ee7fb82c43eb294aeb44d2eb7d16f54fffb43ec1eeb76d1f98dd114943f553ef1505de2a5b512cc7962f8d804782728d83038a4e676582722f1c0e3a697860abea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f83a2b44288d8675e6e38ce85078c37a6b12de1b6690cf7d53359f19ddf7d05379fa419ba4c64f6855ddd6b4b22f6a23dabd22861f4b86f72ed720b89724e8d6c359ac7b9eb8f0a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdcbce86992625d458c54a22909a0a790f99bc2e7e4645051c3f04fcd88a168488f2f0c0505d484a9a7ead507b45dc967eea2368eceda1f430979f2c0dfdf7d2582e43761b8e49ac8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd44e21889a8be006143fd58b229130f4f4398488684cebb8ccbeefdce277ee7ff7f8c4031bfc34d1b746418ba8462cb6b16623df0952c438c0c4a65073e4a2eee0d99ff147a8cc83;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b94bf6ba916e53779ed1732f3c789828b071121661dd91db3fe4f96890c1d9c41afe3b767a7803a8491423d33179e6377b41945bb1ea26ebe4d50e12f59965cf6257906f26d7cf1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8e20970ce7d46072c73d20c681349449b7ac99b435ecabbefe321ba4ae24b743865a2e698a1e5b1990149fdbc578970c820b9b7f615ef5e056ed43336bc6e7ece5a90276ab7b18d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12837afd895b657620b9e3d22719c99b37e97936e56dbe6e3fbe2cd67d75f159401f7b84b768c64826a57f468345c6f81d85037a376136605061b393affacdc642f7d5736f6dd266;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8e1df1e6f002c69d8691d1f0e1e0fb4765892557e6d3765b3bf0063934970d79ef5b972a64028f34e3b89a8a65dd7e604d767bf0c9cd65094afc00f6495530b543bdfb62f4e8192;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35676fb284419abde5936d0c1c465cf8fe8c7b6ebe6bc0a469d046e738d17773b35ea50bcb7bc78b358aebd0f200488a7eaa824dd90d87fc31db1cbec88e26c6efa5500443c0498e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e295aa3231152609041dce6699e6713367e30c7ef8e028af3213911bcc1d09ceb197503c6bb95894f9a0af1d5d2054156e556808bcc41a8a32b11e0c100a6e1a6f3138b5cd5b481;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6864842eea9a8ab26fd56cfb9298a24fe04e30c6eabf39eaa4228acb0ad47b784dbcf5a35945afbb5f6540587d46d62d75f11444cf43096e1a53456296352b75edd5e41e811c2887;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b9cb732344ac526734d6b5ed50ec3adf6d058783dc1ca53476843f70c8f08db05b23aaa9fa5c52e049b7afde6c21a9d94832132651c1f4f3e05bba72b657a6d04b706066d6c679d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7bc3aea333679247b3bc1007825fd5e44e9c444ba17c8a22ce0f9c5698ef939c8319acd1aba72a6ef4106718d0a8b5875b3fe914ac5fc509e79a2eb9248001d697e8440006904849;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc424373e9e706bb4aa95663deffe77c5230db9405802f7d3e88a04cb7249a10e46f7e7e87aa6729c9d33a6c823a4d1e4546af88ffa7e83ad77d7913b260413c06b64904ded70607;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h901ce9ece73656ed84a532f8ef9171cc2290733605cbc2ad16f1a28715c5b0423306c0171b6b253ae05be85d9a03d0de784d8d7ad38d2eb04d96023f6b53062ab491ced5bde6f1b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc85dccb236ac284b10c672a9a98f0e39bf2370fb3c8a2249816d41dd6938e7c81c40923fde167969eacb714e75be66949d17968c195695b5d1d17b77b0e4fe86c01e99a0a9289ae5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49b055b6ae83830fd2b8f0e34cec752011fc0f3c748eb59d4b80a606fcd9c2876e0a0460639117de01f4d7c09954c06dd55e55549e4be79180d2e994ec32124f4f8576713cdc519c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe24a0bc59dcba287f034b205aa98b29da1c7e97ddcc5c8ed73a206c2acaf480885a1db5d7eac83a07035be5785f39c1a5c949616e2a494392ceaa0e7f78cb30767ee21e286a857e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1458cc70c107e07118e7c4de1766f10582be031428c41f26b47db20174f7035075cce970cb2968e39b149af724b77f248f61c4b85b0d2785d529cb5432abd42ba82684343d17292f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd462ea3eb0ce1826df4aabf7f3ae40a070db3d66d8dba1499a652fb3b7dadf3d9cbc0dc3d90c8d138482489dd0ab6acc291f024625ec63f07940f93a43fc10249ad43f13707d7b02;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc10c66ce77148856edcb2af62ffb0a7f605ba3ad8c6ce8a923685e297936427d817e13e063e38e45c968b83297f28494b1c6169a4ea48ac4746205cb88fca31e4a4a5746453a6113;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f19ccb1b0191a74d091cdfa9aae19eee832a436849ed1ae4bc0b9bdd8b31d3f741ea5c81413fa16b7083a75580b93f8f8cd8fe82d5680d55619c5ada5f4dbbe732a08320f7868f3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6bc87a9b6dbc9eba572ec0f7f1baff8575d174fe5da3a9d74f8e6807180ee705d49c68e506767e3731cf00c9b7f8644e9604783acd7187827a0b7de321e820c9c25c4dc909479f8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68703f6170541e10d1fa4d08567dde2e6038a8ca0cf6a55d64bf537f5d2da490e466f392818f0e44ea9d8e938a75e7de84925f55504b3961a9f97832e0038327ec0510f240e474e5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heec68602a36e296c246191f1b92bed541d0699be20721c3fb25754a45622c8475115dcb8a4b4fe83a45c54c8fc497e3dbb4255e2cc4688cb9d84f21c13e90e81d16f7304749531e8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd2af812b33d1fd0f46314518bade7621d277a348e700cb1e335414b90f9077988494d04b0b4a58dc2758ca9c8dca0759d55629ab6d698b4e43a2af3523236da76fd5ee4de89e769;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2adbf9b3f38af1e73f0d580e56d3b2d7c431a66bc74460c099addccc5a875b64cd8eaa7a0475bcafd4950cf9eb46ea0a61d860e92348b5fe91f62c42f5490f419ba81ae6475a0ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb47d3e5c93eafeee34e65c93afb2a2ad206d28f4f5a0ca48ff9ee0a11d113bb752f27c49c89600bb70a6e36d4af1fcf72d21e2d1f6466ce9377aba3a9ee98f47e9794e14c3a42715;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fff26ebc95f2d77a133abb97049cc2ca8cc8844c76a46b32cd2c5a3d100c3fb53eceb28c29c3e9fef8ef79b29f354e8c603d3e6ace3aec5a89bf87b26a7dc30fe7965c5e97ca571;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b3fcd2e57b6092b5adc709683353250a3497d5702017229c34b1bdf23e77204da5cf38ce7ad0138c2850032cebccfb5888f225d86b2c7b82a0b1aa1bad3f451b2384b527fb29ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d47677f07d79befbce021a99b5079403379c7522b15b251a5d1961952fbfef82d306596fa38d9a0859c2f1a4ae2d2525a787ccc5c2bfa0bc7193c222eff90482352a0c8c8d3642a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15a6abe6bac4167945b37c1be5a2b65e6f666695295dc68e9e018c6bc5b707b47ec81ab2318f9433a039961f0ae634985e892b2a4f4f81b2634101be6461854dfa2784dfe16549c1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30940550662b59e38308914b3d131301f9231f1d6f774c512a261acf86a948f3214c0b9e3d6232e3fd1da0c21c3e51958a10530689e0561d7c947fe3cc34003202e9544f5bae65b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2e70b4a2dd16269cba9634b473c4186109fa7bca763bf91b8169e1c1d1f83495a96df178f232383af64ae5fac35a7d02136b11709c93042244cdc39aea07a27c0490c26d7dc7899;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h119205a6a9eb2dabd3220f37fe0ff4bbd31ed9ca5ffb51912e57510677ec9c02aeb3810a72d38c2cabc5aec6b2f983f99e7523c835956a571598074b1ad79ae5fdb0940cf2b6afd5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc31f74641d438c6db3faa06ff3d4cc98120b3c31bf6d9143db6f1c10e75c9373dedbee123caeb39ebc35cc80441d507cd9e3590199735ad5c4e9690d83ced2413802cc2d4a3fd75;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e00999a3907ef8826ab3e17bd1f637a480260b115120afe74bfa5423df4785031f4e289a7c6fd5d106bc6b23a756eeeb44e305689262f48578609b657d013a62aac34564e493f1c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf04e94ec31721b74e8e376ce4094f15144977c037181d50e027fa0267d067cc39f259cef1d072e76070a2ac874b5906d6722374eb88580af8c9994c961d1fa6964a06960a1a24c39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb04ea5660d88a9f528ea96765694b357b8468a54ac1d69e56c544966ba35825031ab493c2b56f324ba66427dfe4bc698693015426dc964f392d3f8c2d1b30b55619bfbb3eeb520b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5243090edd9b9ab9b9c1c0fe6303b4fe0f71c377fb82cab0362685eab3144e4fab4e38006c9b4a6b801dd82d56cb525e02924821a9607f829b10702b33180fc0790669b7fdd243cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e35cfd13295ed39b827157b7a33d71942112f33b9a4adb0aa41dde2213611cc478529c4f1da6bbddb7d52f5b3be24440bdcebafa9222dc1f5a2d8420c1e444cbf6f7d2c252d0a4f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h285da7bd8c04eed11dc701f3610629df67a2c0c9dfd342ab05c1932b4337ee515c371102ea5ab2e1dfe9e27310986a7fe9f3b94c52f1c7f750cc182ecaf5f9c76ca0f661c4da6672;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36486b4c5270ae632159d226ec9ae7e3f8daceebc5602dba2da10f3c7c06010c93cf848b55ab89c20c4f8d60b2b1dddf525d27338fc2a137161a955dd5fd6b7978e618c2c3405ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94d86f2a6f0b16e5e3c8e8e48a3da3531351616afc36cbaa9b85c6546b2b16805f6a2471d27d0d67fde23ac97171375dcf4038fbd3e0d8ebc560011b7e0072bcc4564f176ab843fd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h96d37d8af09f50035888ecb364ad03d6f0bc573632bb503a0d8bf74a5e8fe471d30f5d99c9ace2afb8264180f34ad96f3c7d0438b66f40f76986b07ee7240514899bd411572db149;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f6ff9c8a43e1e8414b80ad668555b41016dc9fe3d1dccd744d5273127dbf86941876d3ebb5745a0c5c9e28bc10530ce2707513aee0e1ea2cbb5cd622dd752e4c54b75cd11e819ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he87780cfbfabea3b4a5dbe171747324075fa42ed7204d0ce428e12145637731ed4f5c51ef7434b16d6f527269d171c51428dc093ef19dd4e1dbe83050956cc8f53aa4e168abb608e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68f1400b032c567ba1faaedc79e995ce9f8ac8a1f2900bbc099fb94668da21904800152da34888ab9643c04ab906f3354d4ac19169ef16ec2ca1802c27d08a37c0acf1eaf6570f5b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b08ab484f76be3a1f398b2ab49992456c8e12f4f71ced84e646e0ddea11489f1c52f905119b8e85ac757b03aca74e61e37212433001b31b8db384189c3d6f7336d11dd25205e454;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88f30daa400f8b8c89b1c50f767c0db2812886bcda563b76e6e68ab699fb5fa01dbacd41be1b8d8200038086623916ce452c6985347d8393feccadc038995ac653dcb01685fe84bb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a12f5f95305aac5c764386e5558bab3a3ba2afc779681766f282416b224136e7b0b7d2ed6daf43195a044ec8b9da87ac68a8d6aa3b62ea70cca1469198305730d76d025f849b160;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6025c91eb6de104a26d081b5d0294fd92f48205142c847d42fd5a6cac8f477b2b61fd46f9ec51970b8b286ea75e5f394caf66b876408091d421a7bd4747bde3e6ffc0fb6735b4437;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12d827dd38b1824c40babf85829d486a3039c391e2c8842284026bf3b75f550597914216731dc91697ca82580de459c10dc49e44636c7e451225c00099106a3b65a79858d7610531;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h323137e647fa2ad5352780df22d237106182dee66113edf91d3c3ce3f422fd16221157b4bd7cdf416ec17e30c287d380f98580873f7108e6332dba2c122f802de3686b5ee6591c79;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd96099ef4f1271efe854ea78165e1c2a73473930378a56f6f1e010a74787de7be6b4ca3318fc0d789d63f89b5e93c6b890921769b653980819fac3b5aa3ca88202bc1311f1dd26da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48c512cc14e496d637d28a2aa5892ac0403367c57f148add1b5236cda077f7463d49be2f5778baf85624db2f3bd5b8552ee406db164f0116c69036470bed9ea81f95576335891d0f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bbea1377a81b6b7eb107015f04d75d77b4ded70583da1adf48221d27ba910c1b8f88bacb60c9c3a6c9035af18ecc53733e95c8ac3baed01ed732e6fd8378230ed39bce822efe0b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd453b48b3c340cd1aa236c45dd1cc0182ab0ecf6741c89c8249fdb06ba5f3cf1d02321b547271a5b23f6c02fbc5cca9b12fbcf79e0de7da4346e8b1d242d5db933e9392a486f37a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45a8ea3a3329bc93e26973efa02b980e1a9a82d8552d5f162a16e9330483f1637ac50501726837d00a73c2b4a340991dede496ea6af9a733d663893d05fa79f2335cd3e6ae71552d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ae9cbd5c24fdc8b16cecfc93685a37ce356fc862a95c7a581c979a7b89816f2b7bd4d06a0770104e3af12e95de1e849eed46dc51962a327ec710c39df3d888bf5dc568549ad79cb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c5b8723643c26739afeed39c75daeda3e027654e1dc4ee0135f10dccd2fa8b46f17a1113c0e0c502d115c49c9e4ac2fc920c02b5d9920612de3bb07a4dac49e769eefa0a175b684;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4bf77888823729cb4baf950c43e05459b26562157f304c2368868296c93d7f18274de4e34f02a249c6d889cabe5d058a425b0214ea9b3a45b7f776824ecab9852e26a0954b0aa71;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb180ef6310eb4a1ea269c494bf67ce40513809b4ad7afeb2c9594ff89506dedf9f43b213b65331d3e039d63795580a62a3fc31c093e0a838a72172a51d23c117c0504b6a04ba50fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f6c564b0d0ae9c4e014945b3a2a28294b4e2c734dea6110a7a470c4bfd37f6b99cdc855adf36755fd37832815da6be4bf423679733041dac48a615e05b27aae8ae8e012b75272db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40602fff1bc3c53a2d9a90b6ae469febaa59a632a9d318a2c08659757286f5d64d8888289aa46afe84ca06e3ee9c4c06c4525008c0a417597b78fb970af8b3d8f580a1f4b14ff56f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9eddb123ce3d1b68083650385c9c4bc7c982921e2ccb8620d58efb1e09fd9c15e420960542a38237c5410cbd196edbae57210fbcf12fd6d951a29b0b86865855d6ebfe896a749118;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1cbd8a2496411a926bf90530f4a01e1bf0689d5ce00728ed9a1c20740ab2135baab39c598f5a05fa603e290cf5b19e8f2bb0c112c41edd533657cf69c263165c8921bf6492da350;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ef3eb2eac9061326329d73028611cbb635b884ea226e3e9b81a1c7478f7e09948afae9dafccc6b278e70a86f5745fdba4f1580c81447ed9719ac1dfcabae72f6063b7d305a2d1d7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h285f0430ac36270a3768c9890fc308bd2448c9e915104cea9f302d33a783bc325712911ecdedfd2f18c0777a99c614c97d2f7755c843540f7d63e78a96ad84c432ff084d52cf443;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1704b7516d4f14659c2422e02430f7d2bfd643bda1ee1b2d6f36bbfa877d7834d05dadc3b7de745e24fa403032f9157797605b8da96d3c534723d425369682246249da2c192c807c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffc98346f41db6c63c315f56d7bea5c14353983878dd08b40b721d6c35bb00af53da982e1bae3c29c33bc07957efa662046b341ef1669bce35ddbae248629d6097691516298b67d3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f69076bfb1db0c716bed3c0abf0cf59943d3290f260d2ec911fcfa32d4870edf1d3cc7c4ba51455c1930e181a6cd30b7ec8ea52048634cae5ea7bea02c0c1bd0ea42da8f9b0c73;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heda1b56764917f37b1e85a7806cf0d2e0cb997206b50eae68e099422fd5e5f8466ed24d973abfbe4ee19579f9efe4e2bfbc3e71074b7c917ed775d02f551de050b0f92e15f7c0e8e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4c0fdd5584cb56476569ed3dc344b69c344f6926417a1a3d5d7e1e111a4f6298b20989e5cd0eaae09b79634b6060b719900d326bd90e1147923448942400a0f07c2be6affacf854;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h216c24803d45115b7e8e7535675c1f3993fac1962efe89a082cf58b7124a7d00ba2b11aa5128a3aeeb2aced14e7ed5aa72479510e9c3b1810c380b1ff80d95ef59bf5000d32d7801;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d33b0deab339e22ac6f4da58280417f502ff723c3fa66dc7fa0cf4f8cbaade398b0405344483369a58673ccf2e8c5af7e8107e71a8e973230af3a917d3fedc73b80e9ba1a9dee39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed714085901340056549a57ca7b44c64471449552742474f02ac2f607cc50673dac7ad2170d7609fb04e8a9c80248c09ade9cab67c4d8cdebe1a941731a42b54de695150b00ce062;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h328070c1554948c6898b024903538c67541e123a1a21043fb0649b8729326304074fc67d92c8c69e08315924dbef1d70532c9609ee7eea190684ba30d48fab737471c45999f8d22b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc34b36a862ec8ca42a53008117d19cfda4a78327e5c2b778b4a62eb8ed2d1363050046e75a880b1fcdba6b552ad0ec42f46998abbd4e3b24b8b83f438deacde784639f31af0501d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33acbd6dd34f97089e4344e619ffa9ec13b265683fc5c71d252463699649a9c12c465b5ab9fbe57a7b8247459bcea097ef0ea2e9c23b36c54fb48e7d07db8079b600552cae3e352b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a6260b2fc3254d3cea90e46302e6f86eb99910202582d4b46762c78f4ff9514883f594ac0110295eb07c1f5c2c9decc0e41f63c92ebf9497182e469661605cf49686efea4b364a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb83beb21f51058cbbab8abaa95270748b563ffbe1a144dfff1b949f65d7f0e9e82a82b4513172813b17099a6cc6edf4f55889c3f8822c12303f950537d934def263b1674e3c2ddb6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86bb4f7786a6313aad03eedf327c76fa2c4464aad7db0bdeef1ec707b44b44765741599d7b977d0a87d8387476a4f9ef5ad509054782aacb75a38d87e8ccd89d2d56fccb04bc0cbd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecbaf6bca5373545a13c1cdf448f980d8b20403199fc79b8f320ef6c1008a5ec081e26f024c44c9667a8a1b893ada876c5cc2c3ea3b866a3ecfd2d0fb2aca4800a87d982c4283986;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2231217047c5569525ea30bb518ad35f584bd3e9bb2efe5b9850e2d6621382320bfbfa5e3caf3fe086a5e3c6f18960e229236b09c5510e473f3e1f80d108607988547502ea4c8c23;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ad7bdf4ab6c5b14bb1381643fbf89346317b7f3d0aab6edfc4000c7756d2c04d8a4ff44b5c86a210531826eb3aab71347ff86a1e3b1a419bc8bbfc0f80c691c12cd5b55eb5fec33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86271cadc1d819f4ee1a3d03d808c76879c49716a7b32143b6166f93e82b1d49e454fae77c1f0ab158d63e53a08a64f551bdbaf2a9ad7c1fd9f5636aff332b82145a751f773c143b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he429ba8a19823a44e75bb2dd4474c26877de4e8e91f220908955e6a1b1e8a98c6d79e34b7fada1f4ad7a29cc94285ea07258c20fcb3f1b02b64d3f372cbb8ff9c4e341caf1c6297e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h201d3c0d5114915cc399fa46d29ff6208e60fcc7f9b1fdb1cc673a379dbe624cbed4bf65b243f753f8e6792331b56e528a820601bbac3cf8f9a97c8f8c9e14f88ec39a2292d16696;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74a0506cc8591fa223785d60617356ebc67f63bf8d0b5bc033084690d9188c62df46d849f4aeba9c5b58bfe63ffc1f6045bfe5e057dfd7fb5de7666142d682b63dc03cb89d2db0fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd953e4ac7112942fbc46a16f0a895e28121aab2b3b5dcd28734a40ff256e54284578f82857fbf5d2d8bbc28334456e3d62c005709d76a51564b84718af91a3149aa8731988cf2fe5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59cfbe792056e17828f2e0f9c6fe62cc708577b66326facdbb053142be2eb0df0c1ecc24f9022957a1d8986fc48c63dba361ec3136b0cd1c07e7fe279f741db8a4be4274a8c4ba2c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hada75555ba7b905f41f4678f4bf82a2514d29e5e87139e1d6b618ca8d0231331388c90f4bdee1a51479e65c27e97b4ac070896a324c58a514442b63b353994dacf289a676a996627;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53bf70b6bc3eb8117799e088538ed8919adde2402d7cca838a338ccd4808d1b5afb3d558a7a135a38624c405e67acf6906d3e9dc744094ee71393e80bbbcb90f84c7b246483da2de;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd720b82ed4bc5a7614c599c9c9464eb617ea4aed2ba757a9250631f4dc71021a3af63ca98588d229364f60a6316db03fcf062a6b042265cb6b7b4646fac169b091b48ae7149d645d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2befcc97585306f743e95e55a25e82c5909994a6e5e6c6b02a3ef0025373dbf83a89d75aff06de88a5e4210c3076df10acae50e25986af23bb931c77ca69e3d7456b48f6cafa01a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb4873b2249c1df8b99030268f4cd2b557dd483ba0c3a62e5f48c15abb22427535c1b12f7c884667f9f1829f95316b93644a0142279157219f827ccb53ec0072e3ddc4ac68612243;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a6999675cd042d979c433e28efb0bad9fa1a94cb88aad01782ee439706c435dfffd9b4457245cff92dc4b5880028e2ad5ff9e071652307c1a9e9879e5469a2858d439b14cc1eef0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e41a6e083e24fde0fb31ef99366f5c6fa66c32f104532416894a95a5c9f15671de3ca15a32b32609b2ab230c8b0f3edb066b085f870d100f14f185e4d6ddefb3529aa36867d11fb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf26e1ff2bf73ff72032af734f1797ca1c4cef9f24eed0a0db3c4555c4518a361d397f40543545b9065e01d4b6844c7c968986280d4b2ebd5dfc4bf6652dc58a7dde21b86bfbd3a3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha15bf6685bafaf6bc00db235efbff6944415df3e355392ee1c412dcd7300eadfccacdda09b3ea65800afc9fbc1e629cb3190f5289d5771673e651b87137730545ad62bfa4b1097d5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2cffab3f822b135b39c7e6214fd15012ab9ad71414096d4b536ce96808cdcd528e4262f367d9fb2bac788a334f4084e56ff0528b9f8e2e9613802e5e7cb373524567ff8d9293a9b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d5e13ce1fcfe5caee6c2b420d31935a2345dbc2233ca198c17003690fe666c9095da73b1840337e389361677c7c366409b83acde0fbdedb683cf8d31cb4eacc5a979cdbbd1d16a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86b8c79923d4498cce021cd1a30fe76b2eb278584beac1dff0944d2a89d23b90c6a747b0d28c650fdd6ec911c61a2427a20a2fc679fc8cf86efaec3a1243f85be3630eff62e08a8b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8199abc7aaed3cc453cb700e243b0840516d1c7579c260a8cccc1a4b692d4279b45d4380b0dcf20580fca66926f00940ccaf341a68000a16138a890001639805bd5b35c49bf3f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe3ece1f8c739b3b0da09ccafe2c4f1bdf5d2f2e6142c190d4d06827cddc99cb028875edbfe86cd31982d0c7865478eb653868c0e926c720cb58f4eea3a47426c4ca3dbcea17d305;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7bcd5e1df9467b787210b2676f60e519fad8d4e40b26292376ce66a49839bc0cd7ec8b57edff36261fc82d352d9946b1bbfb42de5948b8b8bf591d1cc2ea1a7c7dc9361dbeaf04c1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b6a31b26c50e9bac63f354ffe4bfb058901f76a940b57fb26214bdc4ef1214e957f3fc7740ff7d4ea7fa0c7da4a1f35d3a2c8abb53733fe065fd25a6d0ac414e763e58c67023471;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15f17812a9f4ae6524509eae5c12231752bf30e6c5345ff104e76abd04ffc291d7fb9f60fb08ba047f266fa4eacbe9994a3014519a7507f96da44f85341e8d19e553f9c050d5660;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91b679e44321c83f55a13139caed4e34ccb9e290e486968bbaa9abd77307267f36fabab5928db5abcfec97ed11c280259cdbfa1d0a47bb1c693a5897c5c30b7c8f98b1cd497fe258;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50a9cfc7b313ed606602dda82ec9427fbc7fe69218cdd87c51844c7141b502ae2f0197583eb44df0565ca1f1d49936e4ddc27a915b6bfe228f1756d4f08923ea1e5cb72aaa7f1cf1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he379578e0d464851a0b794e59b617c5181bdc64d21e2fce80eb4a52c5ea4d495decb06f5098c341e4f8284cb45eef501d8a5d4ed69fd68c7b2bb7e7415e6f9c52a7835dce8ce8e09;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc19d89d3dd425a3c492144adabbb457bbbcdf1a5075ec93189af08922b7a4dc1b6a8721e08f0b0c575641989157d3857eb5040353bf02b131eedfb8ffb06219237e17af92820d937;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc47372efac6ca61efbf59bcffb8049a32e5afdf1ab255f550cbe0b9ed19dbac5bb9841b0733d686a0e261bbe809c74f257a880965f5ed157aa5b71e8a3409fa4337be71f49426993;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c5ab67e45a6de267a8b38fb2df13015608e2958c5347f830c776625ccfcc8671abc23055213f98fc21bee219ff8c641e7a11c663a6a7775f1ca1560d72b929df304dccb5963cc2a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2026447a9b3809a08049d973a58c8fa42b4d019d01ce2e69e19bb9a8c0a31743a481e07a45f94f2264a81804c52b310522a99c4359125a29da4dd8d7ea7e799631d2463df4eabdd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6f5278c406e13af19184d672fa03629b8c7ff2a7c53a5cae57dae27bab107f915cf57fc5d9f26f27518a735984f118340a6be5629557c0e46b00cb12716198f6a6ab4842950a8dc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8856b86c00f241234140ca78aae7e53bd467e7096003f14fd03423f161916b1cb1a66fc70e4ef6152feea582b7fef364917bd4c7ff65a6e2b355e9b1c07931a7f6638c98444e5703;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75813308fbcc10e82ae2d718dc31b86e28a7c723c227ae615c291b9d544a5176aed5b20f6988e68ecfc162816ff69004776328ff8669b429079ab8af287936706d215ca71dc66671;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e4e36fedcac731f2fa8e12f63343e060a5c391d71f4f1e5cb0b8655c92e46e08f451e91e13e16d45e2ec151b60b28c8db2b2c48dec58abf77db5671676fdb3701603cf401f633cb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5e0bdb3e82d639a007d61ce9073d81bc41551480a8def88c392e9c421d8c34cf9a0e4a09f2228c139f182ab085ff764b8d8e9f496f340f61e2e8a3414a5b1c324cf1f96031f125c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfded48df155616631d35738faff84c39a6a7444d57c7b8338bc14ebf1789d5b047b1ba8c11ecacfb7b2b400a493c4764fbd195309e644576cbbb498567fbcd2846c6f70903976628;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he840516165dbc04efac151658684f5f904bb838880430be0c37335c5ccb96ed0170c912a82a02e7bbb1afaa2db2c451ea4e19c5bf4df9f4a0291df4f75cd6a3f46a81d0569eb0429;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea54c6a54f16f6937989698f2d416ef64a8ea68d6afdfbaeaa06e91efec1f87535acc58d3aa8dce8d34d21c928521115c589a2297e8f9e2a181e8a976be5b84d3f9e64fc7095a06b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98f43d1e2d174f9cd73fb9613f842308403439be24fd8b1fc8737a38145acb1868237d4ab05b7e95f9f1b6652d667f80a7b5ff0b34bbf02f80665db9bcffa107e0b97cf0edbda7d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf874911b05247284f370661e4237f99dee811ef24274737999f543b6f5502558d98b3d7082199c2bbabe1770553bd79e6b425878aaf8b65a78bc886854c444ef87e2ded7b5fd034;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h692842cedf8933733a8ef21176424fe54f3bd4bff9f61c2d7b3cbd4697a92197f9b1eeb78b932cca38e0e6cf3f6f0eebc54ccc126a92cfd41cf09978a9dccfab370c3fa1c4826bf2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddd8ffbd35e21756b99b38870d77b9473f197b89403fe6ed325096fa6c39b3751c1f2469fc3f43f442b88f9fcd9a2dc0157be0803c157718ff6924236101aa4e1661573d58cb3ab4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66714b0f6109fd68423295f93f507023a76a1b2fee33dcf9f06322cea812867ffde1f8a35f9584d5e47d71fe681563568d64a78013615c00300f7a22ca26dda65ed20d66697a5b9f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97999fd02d47650f8c42d2550392598f190e818c2b4eb35025c53b46cfbff6249506fba14574549134e8ae4a33d7b9ad6216c53786a1d24cb018521afa279fccf7fb45b7b98eb83;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa0dd5c09c6ceb6e5f5fc61b79f77bf67fb92249931ff86856635b59f8bb59f42c56561f89f4dc03da8d23915cd7db78cec3d23ec5d170d4b61a2cf2988a73a47cfaf93ad9c88b01;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35d83aa2f1a8e73a67091fdf1c3bbe29c8d6425cbeab0cbcf7f6f3d15814186acd013fcdb8c73902deade304eeb311bb1b11bf19d788c4b56dd3b01a1af5fad3d8daa9e4c7ddc66f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2a7f2b9c8d21a353ccefa1b7ce87ecf56186f83d1a1019207f768fdca230f2982656617be91f5f8e1f5eb02c47c36392963bc0a37e343abeb56ce7e178ba48c6b25e8abcb2343ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74bc9a857d1e4d0038201fbfb3ba88483d88a7bdbe0be125649e224c512ac75d982e2019eb5ed18fba5ca6b971d73ba3abde66cbe8d6718ee7761968941a80e1824295e2550109ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5e1300bd11cf1904fcc3b26f8405082c2b9de7991a47f439f0c8d355de74904e47e1d4f917ebf962f7c838ba6bd959600f4850915fa4242255f2efaafe280513da10188b6efc031;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7ca3f7c30bb2c21e7d465afc9c7e6683eb53425cc37af8ccfc5d5923c122c7c51155aa87ee4ae433f758343b9d61371cad740875fa4e6cdbe07b52af523d05f50e34605f2c29d82;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9da181f8ff8cf3b561bb3122f07e57f54fa73cb52cde3b36422399266973432e3db4be33fc6e6a876189abac54a30c1c4bce45306fe31e86ee137cee23081c5cf4b11b86eef6c31e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc79e9414494d29789dc2462278060381e4fa72b8716c20a77bdf0e072162d86dace6024ec3d76099f6bf63140749ee0bff7794df7a50ee0c231df0aa074e637b7483fac28943bb15;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ac5b7b331e34da57c82615b533d429cb2112cfa13b9b9fc421e2a76d165bb240b80c37fb1d382fc1f3f71f2a0cbf47a2555b35e044e119517e5838c1599f756dea62ec24b65393a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70305de81b1bb6cf0c0ad302edf5249e9685bbeee7e47675f3c03d7615a1345f34e349ef106b110e7d71fde1c9e7ca0576d1de2639780b2a256bcdf933619f2414dba67991221d8f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35f6e64bf4e8d1c6531d40c91a594d0f6926cfef37031445ad0f8d5501649fd69c82e5aa944405878ca8fe776415457cf7b7c4c9ef68fb27259d882118686fab1e8a402eb44e6176;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83b8392a6d1f639da418b9c812db985d5d19feab7308e36d85fb4f49e32a6a9e6c8c1556aa34761214118b3b0598f0c5416597ac780e09ba00b0d4982050285560db7d6dbd9e1c1a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc503f42a6ad8a31287417fbd0b6aeeb8a32e71eec2a11bdfbdd942dd5b1cf599dcefa79acea8ef6acee5e89f144d7d53a56a740fedaf022ee434385bc3226f0214dd9ff28804b00;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cffc4c11db4fb2123c708ad495128578913234e08df6e38c91362d9becce7b93dd4f883f48de9bd7ef1f79c13a32d7bc286544e9cffbfcd78f4eec8500d393e18ce2af7e6518828;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7dfe0fcd3a3f3c56eae1ab28c2fd7bcde876de4177ad8e1f2ca3ada9455f9032879a4cb438da8cd675a9da5074e6cb350327cd17d1dc72bb1ec5044d508b3355d52d98b973361ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1fd5ca0e28c4a962066f0caa400b908cb9d2f0bec583a1dbe01cace59f7ce9b4f4a1e58511eb85be56d0ccbec75320d8c47c0839bca398ad7b1ee2a2aa98a9a82c279e5c45b9141;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e46a5e87a137d5449e804c3b561df1621dabb2db57dcc289df17db330c88e30a76abae56abbe8059ab27ca43d1b7aa2719842e9d8b5a1419ad1a24dfa0527aeaf53c304b40e72c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5d6fb242947523fb2438bde15449e7479913bfa5208ee974f1bf2e94e03fec5636f94a90bb2294d64a622f12b4071b08513e7f2357ddfe61dbbd30b2026ee558e5cc7e3e2c67c59;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haac0964707b25ae71f8c8fae13b37048664a7b65c0c81475dd758de97e68df37d73ef37dccc5069e3fa13602b4fe7a020c43f53a5574b304344b573cdfae0534762016d7e54e3515;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6dbc6798ef8b04560dca909b3e8dc3d165b964e1fd9d170af6b3cbd20e059b3ef8373b16c4b7f6a53c0dce27ae3176a1c9722d41b752ba952eb5e0778de5d595077b7605be6b326b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddff280b6e09c3031996bd0094b057d5c4dab65aea4c4c07254c3354402a104c7abad908fea9b47a0a5a0d0b822e5209e2b2232bfcffb5911a6ce2a1855906d92d8165ddfcec92a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8238ab0b9ad88e69f6f47a4739c4e33bfed067fd7761020b930ca861f0703aed4bbff37021286148293316292c616587d25ea1a27da3a930b10ce549c903d9b05899b2b6a949284;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc93b8dc9435f7bb1c4cec9b5304fd5edfb954486c041a0544639cc942839ffe73dba7608019ea77d376fda7bee18510f3ae27acaefad0d1974e98de07e61491759eae6d4269f27df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3e3752ab61214b8ccb9cde0cee0798bcb3834a64baba62e00accc80ded997f1b2ea6fd29a77cb2e598fdbba30ffb44b684aa11d9048a1d976fb683b0688536c1e8f95c8883eb24c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2ddf88dd0f1b6e74cfcd153e5da77fc8a57305dbddb734c469267ae91a741f7b6225b5e15072d6276bfe28ec4e1d1432639ee94cd29b7eb7cfe71aabfdb07a8e403d8c5a92ef89a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ad4ef3317d1b883253961ec70cf47eede43cdbb3e01ac521ff1070be17ef8307d12072ce970eb99756f742204f346268e969579047a37afb74c16ab0a4d93ac8e132034e008e784;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h196e27091428d99a6e6ebc45c06bb991dd8d6710f86a6372911a0fd63afeb2615e4012906412535f4b89011b93178a56ccac4b09279634f55ad7c2e3366218663eaad1ca04ad5f33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd2c94b549e60fbe2bece11a4a6189dc5c0c5e679f936758e01dee6a9d4b27cc4519c38774a0640bb885119b4a26aed0168126e972ba02e9b3257caabc8360dbff9a8286d0c143c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h901dc455f89527fa93bb85317e5723ffa2b4624f523e0dd4179bd8f59c5efc9c2be7dca56c0fc46e65cb442969ab1bf0f730dbc263ed36b78484b061b7605b9efcae787fbbb7e827;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h755dd08252462a2fcb7bed541619c0da87d74a407094e35117773d87a1b7acf80a8a39745849b19cf7c975784c2deab4fad6b164bde0568121b2478d11b07b9516d18dce1765df90;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b00cd5c42624f1b968aded43253f25b84080b20de1bc8332b2b371ee9f647452d31ff4dab9fe5766e5447f503e541475502f1eb098161c6705747d22d2e65dafa9deb597845353f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4e081c5394dc37bec981efac7f1926605609f9018e3c634b1b8fc4dc3548547897817b24c8928ca24a2033ceb7b89fb87bf4d1dfc7651e95fefdd19b841bb8a19db7b4e25d4dc6b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8997cfc7658e8246dde3ae35131b5aa2b976ec95bf7bb7581ce13f2c0c133cb6ce8cd11609f03e3ddea811a2b26ac0395cf1136ae803c51feb8400adf3fde31b26b9a3d801e10cac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5f8d6aba991f4c6ae1aee0cc2ade99981ee689af992012f34b4182029bcfcbe2f3145c8a3a7d4bb2abed0ce11ee23fde900d55b1525e5a7565ca13bb6c41d8e11157c76f36cd05;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57867d5acfb6225b93ecc1d7bc45001fc03eb6e8b2c40a417461970ae8984467fef042db7cbf071a067b83032773fd095ae975954a429b1f564a881edb403fefa0f67118ae57c483;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e60e388de07052bbd551a9a21438849bd727e9b67cfc0c864ef06f1f388d2a52f8a8cee91800db3480c83a46ddd78365ccba1ebbd796aa0f4ab4f3f2b980e17cb55506f7691204c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f923bf6a74f2d52b46741b967f480fed4051b5582133b41c469df61af5ea7c916e4fec31f05fd91a2a2ecf79f829b9dd029fd58bb8efd94ade8bfa99b7bd0106587854826f3e675;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd0e45e158a229eab6bc928dee03fedd69970a6c34a908f97333f9373386c3cfac54c61893b802008b961dbba616d4119e3ca73f573facd008e16913a5cef2eba985de56250c15;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbfc41952d985de545de12109c2935527006532e451b1b8707d0f1e8d5a2c03b973a2f2aca8b1262abad9bef77d391daaa2e09f91237e3f64b011dc2192f71b251ddf2ce2fa844733;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbad22e6d005cf3465e9d24583062ec8aa61fa0bd6ba5d2c5c7703debad237bbd04d5f123df168b665f7f9e6abbce7888b68820b1b45026a0160f9373e951b265c99ca1abead04d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5d32d46b0031e014c56a558d5101cc5910e5b3ffc2f88b8742d8a5b869d557cf94f360ee35fb0d782d2a01a11695acebc85f7bc5ddec3c680be858ba053cb5a8c5f0ce1eeb46b16;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc26c4d81f2d45a70e9b92e7d735c7ed8d1396a323c165f650fd915fe88fabadc13c172367efa5ab0ce2d068fdaad9e6d09a72cd100d779ec76735e42e6fc0e927ee52314639b451f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3abf573697d3f33b9f5fb585f87be861912fb00548673f74aadd4f9499891bc75b97d884c08eadda2d19be33dc34678df8b755b90ebe5b65445f25b45e05451b4cd13592ce71eaf3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60d33f62925899ded9e11a05c79bdf45c02ae623982ef3607e51e9848f3695ada578c4f6c7482865b2c4a81a3987592a8b83486fa59d2c0930676a2ec1c7a40201122c747119576f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c04d46de0c008654159805b45779369689e131b2218c256bcacf758fe5b24a1d9235241f24ff36c4a4df607dfbc6ed792f26763a494887e9d8b86036d71a1d194d2d20cee711e60;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h363af18b0025f21c65114dcdfe9467717bad0b54f4c75c492ec6a7e8b4a3813f6e36b30bc13307be83a814ffeb14b45ed60337d0dd37971b0678db1491ed5089c93b54d0a987deff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e4aa55688c49adeb0860bb85ec6561f910c520c74fece96cb67d06c2f609ad19dc341b2b4f38814fdb35295c235ac9b7effef7783bd8ddb1c958b4b38c5387e1a2021b9e656a2b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f7378da17f20626a316314d31c768c17f4016acae9880f270184f7bdd475e2c1bc309b9f0d6933a5f775e72a56be7058df73c69917408c222efafd4b37728bec52fc55889522552;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46e9b8bd3bca1192031a424a3726fbf16e3a8173f95fceab64d3e2db6f97ae3862de1943212c7c4889269e5abe945fd9e008f394be4d67b462b5257664a3f81cf6d9ed47cdd40a7b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21612586822d62bc5f372a5af7d456ee3b378d8ec5b1a93ee1cc66ec30f7e0d984aaa321ea47766559965816679efa871b1af209da0b4eb1fdd10bd080683dc1474d1d215ce886f8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74fd1274e809751455ac24ee29972f7d0d29fa4f2c00341e653abb89b3f66ea38bbff5b37aa5852acf38ef1d225d971dee41a603b236d9f3567d0af30182515be76688486cf788cf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4515691d1e4c66ffd78cee96258d8fa15d36de053f29abe0b16e59ba2501aa7c558b7192511f76536faae872aeadc0eff855d73ba9e08cb04f1104e161bf5fdc00afe0da451a6cc7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e953f1b1e2b415cf5e98f51edbde8cfb4fc0fe66d69f98ebcd835ce5d21abd67ebfd4cfadadb3dd6d4072eff690a809309d085f7030a81253286f1e7d7d2036c880fd8e38ee8009;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec27737469d141583f7fa0af2852ef314f4ceb85efb16ee792428ca5741b7146318fa9828d222d90270672b63d8d0f61de98cb42ed695df9e07226bb3c1c1d8518640cf67a4e93e7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h201e50002dbf046649a4a077159cd9ad4c386dcf30f7da086111fa98d6a575a7ca33431cb510906c6433bac938d5da187692c74f58b7b6ff41c4766eba053b72088793b42f003c7a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c498823b5be237eccae45ed2fdf0bb5f3b9effcc10a3e024a38ff7cc69e1540410312a27be54ca4f94d575a05d23d0bba3b0ae61cf42711a83594f93c313ef4138e09f832625f36;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdcc37c047ad24a71a3c2818a3db1ec4d9fd3087b8a733c83f0484255e5787584d691fd898ee513992de1aa20765365f09b2724a77ee55a4b6e08c46d3123d3e5d97d930283e8dbff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6456a89555e7fcb106a2e6a50774461f60053dcf7ccc934e766256ec18a8c9286a89790d494496e2c3976594e64a6a446bbfe784db942af41d13198a1bcc3b6ee5a87d23469a53a5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h698860bc422618eed53a3b12725143f5daeeb8c0b0c8fa5430fe6e8439c37c486145ed57b97c0fea53ad156e0fee2cd32b44ae17e8d53ab680a3f6dc5174368e1bfb341e5cd403b2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafdd56273d61fcaa43eed446e037be8a3d9477ce2ebcc797b585b7c84de993ae4781ec64ed26d86bd6ccbd7097d5c9ac87af47375cd5a663a2c6439fdbfa50ff9e754dd9a7ebe9bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5610fde3798a4053848378c13f4b92059dc79e94187eaf18e605616a18a5d8b0e9417f226191f711f8bd95645d508ca135a76fc2f3104001d106e6346de6c5b2b4b2741f1d5abd13;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41a481f73329086ed4254963c1a26993939ebab86ee0092d6704a29b73e188df098e024afd844d6b5a5940a55260f918721d3812b2a2465b56a2b0b8b448e5b7fc9aa05a9533dfcd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h692cb145b702fa37cd1e90c1a033ddc55d62eb3e0eb672259e0914c062fdae0110b02b52a64ed419129242adbfca938e8c21780d4b860cf61d1425bc7a6578fde476362746a5e407;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59413b7cc9fe219452cd914b21dc69da149b02b654b6c4ec82acf0babb306a2bb865b908d8044ab2d6806995e4419fa00a61a933203607ee9636e005b5d8b5721cbdf690866d95ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf40a178633b9fee87376ff9398f330bf870681be1ba0a82f221a6426288113cd02872e1f71846d7455e2b33950b4dba5e6dfc923b0ad0cc0624f1016def5b06dd8d64dd02af4486d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ed9b359a9114457f0c3fc45e3da0c3734ef0d18f94eb92b41706c3e439b6b37b070993b012dccb8c73ea75f8203d2cee42663e2c3b6a61bdd8bdde25cf0570c74f9aac5368dfae8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71c13bac67fdffce6e261c6b250d8c0ade471a1944c902b19067b9807e957cf8e8765658c1a2446292037e17501967c2451598d0f86a8b5291b9d96153a851593b41560bcc4f767e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11f6c2c1be901c337ccb323a2d30e5bad635d885e9b63f1e855a7a6326da3b08776659112088abce1b58a57ba0a715fc46a9bd8d04668b63a971f2beb7b8bd794e97f67b2de525ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71849e7b0bf7cbebe0233b3ee46ab26d2f8c87d41ed7299e3c5d5f4d4d3e1adb0845d0d4ff3100ad7ca90385203f1457ff3a48e136b85ab48658a0a5a44ee6ddc49e8625b1522c38;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86741f3ed2e3ca9671052084fe2014922332313d35f1c4935653d20ea22be4cc66ec08eb65a4dc3ebb36f8f01d1fdeda88b2b2564554fa48bac73e8b1bfd86d1650bd1ac1968c1bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d149ff129edb5570618ffc078f4558e2863c9f7f5a6989de35d471df4328a4aac09f994819102fac1d7e77062f5448fc4f039cc5f3a02f83b8b0b0c5b631d913631004f90b5bbce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f6c07a7fde9db975051b2864676af5ac3a2d667f44fc6b3f917e5ab6d6eec9814ece32c0f66336caefbdbc6ab5c24463bc898f0e0172c797f14f23f3d9ac057497f9e3670911ea2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h962f470df893cb9df32a17d334c336752f7bcea84ff08751ee356334499bf63574f62527e43caf90af46dcc8037ba41e2bde389b488fc9ed9c8a7a41422b7dbdc89b59d6fb72b4d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60ebf35f20118537d20a6d75becacc451f87f9856a609294849ac2f11134e4c413fe84f1473f137a414efe9ee47014e824ab42bd7cd716d566bfdf4bdbd56014da429ae49360acc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb17784784c0a0b80a6e3a3e30aa53a1d47a63498d8860e39cc2519dee391375a75e826356c964ffa9e802bcf1f151233b71946b26a7b2994969fdb317caece4cabaeca2058ce917;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef3ed367eb76e6e5b8be693c198072cc1b18d2dd543a1cec9386524e33ddb62835eddff04ff07b343804b903d24ef9ffdc37d3a04d1b53805d848ebd9d75002c4202f676e648e11a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69546890a357dae375ea413b9ca4cb512dfce84ae7703310050958be46d614657b63d60fa8b8a8bc6992a8af205b0a3c178d31b70e9c6c5d46f61b65f13a27fa7eb42fc60b8fd69d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d0d8d792d072eb599b726f0ae3d685a67effe1d35c5a20e03f6f17c8aed370986968538ddd527d9b96b1b424e07049d20d978d6cec5d8f0df836177acf95cbb3cdb4accae7250c1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b6a750bd371e31e371f4a4e37c4ab92d3879b46b5e78f8eb0d1db6bb550176cb2d93bd40b2bc8b0d6b1b806e0b92e144fa08f20a439392c63573b138b45f59695740b8248681839;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e6f0f2eba19d4babba329cc46ce20c64d3f3e7221b8d85ae9807c0ac1213daa4189f39d52d56e192c0c473c309ecd06a7110f53b1ff1b8f906f27d0011951e082fe3fc645ce5680;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde79c5b7384d36035719978652b7ec528714f3325a7ec0dfcb66989125c5b936e1833d06d21bb0d271b326b524cbf837f7e4b07655584cce0037c51ada453985fe17a64d009844be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ddcac2f6aa1237092db909e15839fafb6bc39d11ac69b9fa2a7519935b9f1e640e66f06b2a13d3c80cb7ec4801b711e1a93f993371f001667f4f1dea85be347551199fadc8cfbb8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd97bc0a87f4ef95fef3d5368b6db53a7676a35bd010f08af7558feed37810fefc8b0e612c177af148710f9763faf79b75373fc593ad965524c67c3c1e7e925edd15288139445c2d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha761700a110621006e9d9a5f6d6928c8343ca61a974ede6f71f3f24b842c685c73e9a54d582f0fcca3bc252ce2b3afc90b80d2b8b4b12cab90dc5288df19a50204c31fb50ccce2ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h384c69b20175cf0c460f424fb0f8c54d28ddf3aa0ffdecfdd37a2ce5a2e7de16b8353dbca8dcedd7c68c50d125c729579210df5ce547ee69fd7f458185dcbf25fe6549c061da83ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d7ad576b63ba570f3b609c1433bcf0d0e0dab94c6e7a9ed228713f9b203e9a976559bca339b591717535eb1193f6eb16a73beb0aaa72b454b782e57b339860866e017c0655ee8be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8f390addeb2a3396623f1edf8c70857fddf32606de4b945f113a817174f5af339be21b674b97a84521d1ccd0cc074f52d915304d5884de5946c835e270ae2d1d6a402aefd0542ef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b4051c45e9028aa9354865b791319a2e8d705d4c4f38163ad3b7085e5e2d967c2aa696e1809136926af0ae2c037949d2555a9c9b4742aa7f9bdd77c8451a80d11e61d1f3dbbd30b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0352350aea3f9cbfbd05ded2a341a1935ccf51b7ed68aa18b8a716c9f3c37d06261e87a93b21a5fdd1240f05a5505a9476a93cfa593123b4c43731a68151bd72c531f37e0e42093;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d0e0a86ff9c3b6f1c5ebf5bf63a9e5d6b71777b639b53f697dd0c8b431bd5071ffb31235a0be5eb670a230af12c8d742dfa57a6ca9dde2812e7472b0a8dbea6ef58302c4959613c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe07f81bfe9de615f8f883b9634ad086edf42f65081cda48861505aef6819aee1f3cedba3921fcd6067f17814a5b050cc3a1e1652c87407902469e0c860507830d17123dda4d0bb7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67a406e61d0b43aa98f752b2a93fffe2a6617e424925bf995f35d0d1be9456b08927fb4dea3f7d784edd2dd812a46ee309eb0c790de11b852122e741dd7a30540e10c573f31687a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f3dc14d0810816976d41bc04f45c5f8b5d1352a57ac874f9c913a7e18a4e9dbf0357357e75fc0bef76f85e33359b1ea04f13ecc80a82550330906eb48f6e03ab57d07e95b37481c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habfe8be53346c672a0b363ee7ad37a7f5a75adfd6c34eb3a2b618b4a366db84a2609f536866fc7af71feca1e6a28a9123b30cfb0f25b668431be23444c34940ef4ba662612291b37;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22fde268b82572152e7e1c91fb5dc390f9105a0abb2f8a4b3dcc5ca8a1a118524c7db85a630358f62504924562090ad75d84b58980a1ac40ad7682b24ca57da7bd9bd81b01b2999b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9123f79d7d08e421202a817f8708dcb81d9b62cc75e596173528b8df74daca0e86873da567c78736ec5d1edbece8b05bf290b6a607582170b16e4dbe39d522d661d968e04ee2771c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdfdf665add9fa6468063f7956294cb859252b3358044b53ef6841b2b9b48848f2e4bf7974ff51af6b92743431eda18401e3f6191467aaf76e701963a66e9c3f6d53bc88183ca90c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97ed2af74be3dcbf8b13e16dff4dfc7d26c31bdec0f8d4315c6c774624dfcd345f04e335cd884f79d21bba03b18e7f4c96e0dd819afd94b6cb693ea18af16bbf74927b9d1f19dc1d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h288c323c0ad825c35a62ac302e813f8582a382987f5bf6f0e946a2bc411ddfd4ea9c75cc7b3d5f0d7d081122d5f896911d0dd3449aa68d78329d166c78fc9f3af81e4c0666625b2b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d86c7baae1d773e13ec0b0d5016abe2da2a2ad7144b907855a8e80261a6ffa3ae5f15ddd4e5becb52455fe5251e110eb5e4347d78a505719b873b7282e6beafff53465628b4e8d4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha583e682080752c3f4826c150c1336411a64c78b68fc8488f8a50f69ce77cb99ef2b0d5ff104cfd5fe6070a24c2cddc52a029be07495cd4a55e0ce066e4ee6710c9b5b452a85d4a5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69ee5db5566fcd18ed93e40b10af7be815bb8badd65b6636948f01ebfd65d1303dd2408c24c8b2471e2d1213604d7823f12a420d0a5f111c9d548fc4e06e77d928ebb011e6be4053;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h261fbfd3529297508f8e9cb91ba03f75b6d0a16af6b128168d5cb221917d2a62c01139087c5907522d84bad640d5c6cd2f1e8b7c2bf893ce542c5d003e626dd69f7896523541fef7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27a38111e565a2bbde80a9b9e0fe84c7f13893c133470baecfd9c7949d4fac487b6b39d10a56d7d19be10adb01208e6e7334a60754ce0303c9691ba2db90ebd8326c642ae5ab8db0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13eb9f9e4ad91f74c6512ab613e6961dd30df5c2db72130c0d1a72d227e0310cbe1d14c590e431c19a87ece12f2a004929878f48994a6cbffa14d3f41edd7aa1a47be5f3ceb464da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3be71aa8c5aacff3ab2c095a449adaaee8728275de751b60dff1ca94c9e39943fef1ac9b0243d512effeef3b8aff7729b1eaa760d5741c0cbce1674efe7b1229ce0e9978f4b0566;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e4f698e25893905793895657e80bf911dc85fa33150b3b9dad76500278140052ea2d05e51c977446e254e8d3899d62e666e45dcfd06e311eae4ac30f6c025c8994de8d0dd5e9a22;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a37e9cd8ed05b2883cfe1d1f52d5884d4c892f1a615d425d36efad84d67faf32f682b25a9546c61b00a089a52286a3257a317465aa6c541183c202714b938b252755e3bd8a5c16c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4dfdbdc08bdd808713bd3a4c1a6d209fdc926c26a3dea6d804e1f1414aab807ca02b0f6339a79a142cab5e309d2d31bb849b972330e863613a37ad5c3777264f83f6af97844ce84e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52d88ac45db6e86e51c3db24956f9f560cee607040157379342c60d1f305db5d7bc26936fb8ac4017859aa07f631236d599e50335bb83914284ec9847cdf2438bfb7569ec7fbd5e8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb059f6279368ecb7b61f99028431fb43901073249876ef1d76100c4ca02df6c33459171f2ce23540997d5bd34840b671f2701b33423a3b7bc2aec71aa57da2b1116adb49a9c581d5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4deb574777e0f81b97136242c03110d5273a29fb553f1547e80c6db61baa8463e1f98918dd9d39ce8900e71e44612c3dc275e054423324b7510a980c9cfc8ddb53626d6f895bfa4f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f4ac6ac8d78615a2c7027b590306182abb342d5a839d3af2456bf255dfad4b5f878aa6e2944257b431d1a276051e5272e8621a5bc527c824ef8394edc78d14131c0898794a65a1f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h804aa50cc92a2778dcbdb79f27403c75b978cec17785109aad1ab4f0d9aa2fc0483bdaac23f0b4c7a84f1ff84e30f2ff2cb3fb181c7423a86453c14aadc72494a263f179dc5b94b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60a1424483f2ec62ab16c0c3cd9f2167c301b820dd60f39a227cc84d59bcfc2172622df4610bf50b31c7b598e9806361e479f13432a1a7f9f5a1f1c8cf8512c85ec970b8c521bd58;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88707a40ff397af6def988d59c08db77135a61b0faae2163fbeb5d0c84c186e7283ea305f286dc3189b076539e86817cd9c93fdcc9514aa44f9819203b5ba142ea28e9e2a7d77b63;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c1bdfce39caca2ed59d219f3b209afc104b1025dc999cd69ba6a4e694857728b04841a09eaa442fff8d52de6ffaad8db2611618ee94c273a3766152b48d2eef6e184f5c34aff28a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h452b30d8194d89538678dcf9846fc8ffa298c8240e175b2d81c707ca4b0e6aed7a9cc98fcf3647639394b5f67d248892cb35b60e7c19b3cef4f1412caaa61c660cbeada816b07382;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68ddbf5083dc2f3ef9516863838d5cf6bd31f7a7a2f39fef8a8e96e2bcbb8d6cb48804499514400ddf574311420c7fffae3d6553f2f9ef03b30aa8a3c2efb11215580dde42e2fcb3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0b555b860012d4090e62773f3a71a52824c4714e3e4db3fe4a84205e1d8fb1ceca2329b422f9128cd873c0d9c4b419bad8fa621bfca182261ed8b003e2b7e39a046df1389750c37;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59ca195fe042a3f1b2e3256dce4561bf9ab2127ac7a018f5ff32bef70141eeedb7f43deaefb9bb77ecf6a38b02e7f86e49c63de1dbf1cc3f89ceccbe1cb56a56b2af6847341a614e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc65c472f6f224adb5ab1816a497299d72878b342ffdaf5d887c93e5505dd08a3bc4d37fa4e1b0c20fcc259d34957f7304519e3124c424d0f620b321b56c1456260a86ca3c886b218;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h111d8c15d9a8ff8eac26886ca18d71d9ccf55d06468de204c425f16808724216a9475660b1fa46b8da8ffaa06f39c683de2de92162e3cc6d298e7e50f6e4b4f38be4306b8960de8a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he00347bfee8d6f78fef1fd59370123d4a824fd4e83bb97e6766299d799ba2e6f1acb6137996f7f569f7a09f47bbcdb11350949a28480037a3a22789adc5b409925cf22b96fd8dab7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h972f81ed24d7215181174a1e92056c0f12f1508ba13587ac847e1834b91059a3aa992c0be7913e536c8a4aed3b5cccf45b147ec44d9993936406feae6a7137c5b504409c14567e0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf804113c5e3dfa4cd61c653b28ac1aef33755c021cb2d86983ab54a4ca16f0d69355d3addf568ced154944159b915a97e667f5bcc10aae20accdfd49e77ba3a3972b7a0f7f96f8ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e74bbb27eac650b719fed80fb3f29655e9949f4639cb367796480c7bc47b719976330da93a2bb8b53e507d2ee617de87205a2fe42a766b804ecd5ee04d78112389402081b0a357d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h768e287e39bdfd94ee8aec6ade3e2608c937344b4d0840bc3f1d2f4759c96987af5d987ae8079a8048aa3821499fe65dfd8aa9cec252e22efda7678df96be775938bd04069d5f8d0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb88d379d9710b7fc5f1a1297e1b34907b28dcc413490fffda55db98e985ff746fb4943828f7ef5841c506df913b0b58024dfb74cf5c4bb1985759dcda397150b5ae9f2c063a63527;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54e318fb1ea05e5bf5a47ef31504c0fbb0461e9df3b2d7eba63f9b59d34e4c9b6698a51ddeb5c6e7ee053e0c47646419de8541a34d51a08f6ad6634cce6a98d069f050da3cc7622c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0e324cd8356eb23544bdf5ff3391893fffc3208588ea9e689f4f5496f084150b10bc74c8c59ed9d720b741073f2040ee59255b9479ec183bdb823d5318222da90e9e27ae536ca78;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b50e66fe87f21faaca5631ea00712d279b8d5a0755ee1626ff9d34ba6d9f03220b737fe8e319f76a01702e8b530626ab3b4e58dd7e9fb07c6669c56e7ed8ad72c42e33e2f910ea2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5682b065f1c770295ddd54e14c1f2b32ade06d28bd0cab9875a22e5ba8ea51099aa74fcee4e77bad0d16e779917e8cb94cfadf82f8c927319d2a0c3a95fc980c0709be37649711ba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d98a2cb1075f30862ed867e0bfa798850e151fa15d5188b8a19d9472a7b35af00c6bb4de40cb78addba13686c2e8b60514b9580266108398c649584528138a27372fd79e4ee5d1a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93d1a6a2645d8f93c8e3c5fd349e882dcb5f4ef026f5d2be9333833bb106f1c4ddbec798472a030b10a7ee3edc8f8653bc67aa27dbb145350e6c3684de93c65afb7651aff81de7e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h505872d3104ff1e80b5f15b7896c61561f01546929e917442d451ef4ab6e0d3e189dca410a5202930493f2228a9d3bb087b6fd0bd7703c8e4b68d5a5f1cbb5a6c215f481c4c630b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd64de4674ef83b29270c07e1319b2be6735600c7da3920283916dcc04bfc8412fa2bf6de31add3fb46782805fecd10444e3a6f3bc7a81aead96930b9a9087074bcea527cb2b257d4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h540d254897d974b920b38d05388c3a6e1e6335a8224ef0bffd96500e03002d8b938efbe1222bb45212aaa1b70906ebb03a44e6018a52dc877a86a685c1dc2fc34cd8fb1490a10166;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b462d12020b604598d1c350a60347022b07e439b08ea0ac833e54f3105b43dadd7c57357a9a9245ddd3b2ded0034aa78607f5748add7f188109efdb37f46eba3a21f63e88e6f9a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c5219d7efeea43aafa7dea49af5e9c46ef69817344b5ef24fda4687ac4e6dfe0bd98367d3682c730415ba8515a11b4adbd1b3d9ea22323876f2b02d0c86c1fa613e03bdbda37d3c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8cd9e2dc9d16af213f146770c50bc46a34f86114ed2be7887c4b6dc64e62ed5ccc680585fbd8e91d408b58b8cdfc33da3d2a0b1545bd76eef467c2404f662eb6e638f9a66b0324e3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce32999933ae98c3e0dee75b8eb088e817e89dee60808e1903a5ed12d59ac07c3e3931e4be67979d09611baed578d5df519a9be53c7b29c442759c538425492a836214aad0583304;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef18233bae2a6c6a733a5645aa6fe968145a9833c7c1ba5b57445645b64520438aa87a64994afad1a9432a36019d61846baa166d2d9e8ce8fdef821e51f13768186f5fc369f0d054;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61d729c6c91ccce5fe90432c6eeb07ee6086457fc48d5e594f8dd5520ae63c17b4a4d3220fd1d54221a17c5f820899b96fcc46f11a376ba4674de3b087e7a5e3220f48ae2912f5fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2f37e7df8db2b222db15b67f30f8a5dda8efca0010c2d2bba5857c961a1dc2ac7e4db0bb9a711caf0a99701bdda67d15c30e6f3906084a57392da4ef9ef124e1a0dcd6fffafad8a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b18f7f154c651a6034057717722069d9e0dd186a8811d447f4a46351e85a09a209ac0c31d82cfb4308a01de6ba66732a50352b8283bc3f4aa4a8fdbdec61a96f6c66cb45cc03651;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h888574c1a51d1f08d03d52664a1c59ce2f9f278fca67a65c0805c37861a6036c1b7127c0da583b501a0771aa3f500656423b247bc6d05850d118ba7e2c6926d2deff2a72075df183;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha47d94dbcaddef847b783a470d25cf35037851182101226ea48009ed7994208fd6ff2d12ecbacc9cb11709d3968366c212607036ad49a3bea98bf8ff5ddd0f5b07ef041677348de9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h821ba420ee07d9ae7a4b6bc63df078366379fcbf4dd4f0eb3f5fdf92afcef4f8406648c353780cb165be756c6b579e5252f750caf342c1be06a03a337ca3e2440ab6126d53dab219;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8015eaf73d054365329d2126309d77f339828e1c7af460a69d5ccb20f6be4e2c8e59f14d03bfc44cb2f250f627e02b559d6fdd7d760721cd31d82a3e96217fb96efaf9b2dd104db2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h608d702175917e67f5bb6717b5c0213b2c1657f68ac672d06d0ab5f9432215371af94bae811ae5fe7cb91cf67da144bd4109673b1bae12af67509f4ac4ac9537a242133cca4235e5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ec9f48cbee73a8b63e85928b175b8dfc7579b20f6c1d0e2432b17224bac8fbef056cde0a4929861c9ffe2c124eaf00d6411eb235d7ebed218db17a0dd7daf1f6907a1120f43a658;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63f859827ec2b4d962ab6a7afd91726c540d6ee145dc15bbfba89962fca849526119fdb678be8badc1a3f8da9ba5c7e34e1b5871373335ed23cf335f2d832d63fdbaa6014bb63fbd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7b4b4cb979e9be954ab84b5a36c8e6f0a0276f2ce1acd5184d40fff07f2e6b979292ed914acc760890ca9c44bcceadf171de075277bf1161bc90fd50f7290f021a07ae1b4a10aee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42e1ad4803199f15db0d3483d145810665ee8dbc0fffa728fca9a895e44bdf41ca539f368139369d49a76674089655fda167ce4d7f2bb1ab4fcdd0ed16007c7658b84a8561067f94;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h840b4a3ff24d2fe77e9a25abfaecfe7da5cbb17218c3fb1cc730497db284800046707ca1312da1afadd962ef6a442e254a75a5d789fe81905699c9bff2659f5f25efaad62122c260;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6ae1e3813ff0320483270bc3dab05f0372cece9e0857de3dd1aaa23e5b47ee93bcb1a85317dc64b4e7a3cef96329b69fb2e47b008e7cdb6fe7368a719c55e30743d1759fca3c8ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha54fb01b998b50196699195b7b90ae6e464ec26eae8820589a2b756d2401f0264cdefd43604dd5bd909caf1fc21746063a9e34841a12d17da779e0eae351501a63783c5cee0b92da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6624cbc0ceb2bb2fa554fa4fc1f5d81a0fcad50c9575133b15cecd125838e92f5b29b88534c28fb6cabf8f909c359287ec0d91d3968d1d133623d17291f28812aaea6bde7a69cbfe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24870772178af86abc22327e2adde37c7453bd5ae65c63c80e491f8a917fd6598b404cb02a017b9d32864c540fbba7bb2bdd929cad7d13a036aef08703fe8f7e5fc5651b9f708330;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7292bf45524e220e195f8ddb33188cca27c2614eb84eee1750afbc383b1171f589fc87ad3e40efbbe8feb877a66f309bd15c0a3f653baadbfb638eec6f1aac6fcfdc4151c06c9f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3d6bfa06a4470c00b876dcece9e5c90a2f5464e0753fa355b8a0eac04dfb7d49a1124c164d896bcf0896a10e2d2e5649f1905932580724358c164eab16556f19488585c4b9f90e6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99426e830f3971a20e0744b4221a9c4569519b1fef38d77fe6d8fa7f7141b7c4038f35464841fd78984b05145234403d564f8283cc6cb09cdf8e47178c83eab9ebb5cb5c22dd44ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fba9790d24cc71130a1dfb6a422e6e295cb736f26f3c3447318847d9a73facbe0061c77cd116e5ab1fc5af4b28fe9ebda835f9203d92a3da5161b119094b0e389fd265548df2878;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b0f28339a9a22a1302cdf5b28afaaace92e72a18caf4f5f7ebd9c8345b2e0aa093f2aae92e9c0e0e18648d81176aab4e85a5ea7a7d81a522ac0869583ee812c9238a4d25a74cd3e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7cea7a67af052142004637446203edef0e57e16078bfb1fe45f5efe7e23546ade21061de946d44ab0adbef3d0689a4f7750ab18e306499d63404d34390da010f22efb24b2a9f4b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfbe2fdfdbf81e1a416ef48d4d23cc10f8147807746d3dfe852d9d469c0fc4246c53760e65de391c9178a0886f34cbc19d95f893049a9f0e6eb6934b069673bf5a6f32e6c87ab6c72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ea996c1c55d26070a374782a417fe7e31dd5e31c9d6b760256e84913829f66bfa747e2244192e3726a721f06b29741773d833d5d76433edf6f63afaf7f0b2962e9115c454c00f81;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4426878f4be0def403b68c4777f35d7e88524d1dfa464d69c50793fa8a9e0401ac30172b94872f1c7ba2a84352aa9a103444de6b5e2905e4aa6f79c47ff28d3bf2c9d52b2a793a91;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc238b8ead8ede1eff35009e60f4facb20aa9eef010d36a7491763a9c8e27671caefa0118800cc82f4464196e1249ee15fd24551b6220ae46aa017d6b15c97fb14e740774c6a86445;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5d032efab00f177e47cdb9c5e88490b3ea2f8200e59404ab455ebaec2680690f96cb9b93af388bfff7f349509721bdde1c818b05bdd0fc9c5dca0a7dd5755ebd4c0c50f6c8f01f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heeff39d5371648127cda43d19a7be122a4a8aab0c7f7a801a323e3ccc4887e0c94db45ca9598dfcd410eeda3e8864ecaf325951ae1a5f8571a59b77f7a4b1c117d125ef053e7b67f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddeb15068026d1cd12b59f0c699d5c341aefc35cec8a6c7d92ad362556bf27371b2b2dbab7d5a9976064e993011e075b8e284f4a1fd1fc18be0f408a2afc1a0d81eaa2f46c93b21a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c0d748cd4e5b70252a958ea3c9343780b1a4919924b2460e1b720463d692f1c5d040ed7174e3c11a3f5e7ff734354d3cff1371bc82a4737069bdb471c05bbc7e46583a28c0c0adf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d51060f59a29acdeb302de08cb76996cf212ed5ea6fbba0d915bb67478fa7769371966f41e8431322f87ff24355d6be7560f11db10d8fc376f201506e083d50d23d855161273fee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6c54f7779b217fd5444a9b33905790e5ce2347486ad5c39d892a02089702427d00f26690b967fb9bcd64e20d35a2b71b9ae220be39c32762a800f31e4dc01d077d9865d990c82f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c18db512b01d07c32963fded1579bd2277eb324d4672c7baea823f1efb8fc6c5e7ac4464019c13172eab33b9a70c127f41a1d949e13a03c310bcc9257e761271017b4df8a8966d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20d2a4acaa8fceb70f6b2b706e6d3867b9f0cbc65da7bb1dbcb29ff7e187c168393e956303a5deb67919d10536b72284fb83b91871323defe52aeee6254a835046c369c20add4120;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc65d6aca255cb4ba33e8e344a9280cacbc2a02ff4c7dcfb2ce894fd1ec0785fd2fb598290e8527983b4d013fa912d620860e8aabc8e315b5a70bd08df648571e2dbc4f417da3d16f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4fed9dc632a990ce64a94859642645bdf2aff26051c8add6d31fedea9b7e4ffbfaf913593e42aa285f7fa9a6ae3fa709fddf0c6bf5ee0c34a8b0c585dcf8f6f8f69b7f5ac06d2e00;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a4c8b99869920833d52f692c7d78c58c834f185f77e580eed3eafc83f644e739a3c0c866b279033c41e7fa25c2b4aa73a36138f0afaaa3ca417b5c1ed7f669cb85241f2cce51022;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf597b362be99cb5e509b9fb6f720f1d6c5d98037502812a3feedb3076e668961511c8ac09a727c339dd75b68c7f10a0921525dfd39545f7467862ff25732e84aa422b08ecb219ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc44be40c63697e9e6ce27eae12877b59a33d5e34c6402c70b811a2a78f452ed974774417bd44fad43a6d86615da215b2ae7db438a7e7fe6d2de171fd81cc8ed6ab5f49de7286fc1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42923b4904ca9a1bb67803bf39ea5f7cc7ae553792f9409c6c6dcbff8153ab343b3ad7e1f8d7e93d6540f5e21064b0a0bd7ba7b9d612a7a04b286df2fb71b17320d71c0f2c25324c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba94c3b3c968fb9726a044dbd0fb668516f7f4ecfc428bb312e856d8938e3ebaa6fb9810accf658d319af7572896ffde45e3c1abc43f8cd10cf7ad4fd0a48a58dc3c3fac18fd8446;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91f650828af1f42ca848b31f3815342bc7ccc56f0995be6213ce408efd79939a4b1489e480f64fd209ea12a1bb1dbd38ea8e9874ab00975a7c9ce0d61ad2d0ddff31ff1e2b6648da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h184f7544ecc184191912ecec03af9436c69acce2554a7eb1606b1672bc5aa981bdd3165dbdddccd0601c5a7bfcef508da19b0f57e37bfdcdece47b5f62185e454996a3fd71a48796;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a047bffe12fc5bae6459a909780897686e208af8b3cab0431c8048e83c7d3e79877d1a1962b22210e08949fb987631f8b4e5f2ada026dd5c8c54bf89db849b6303d944b2a8fbc0f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf14fd2425e20d3c55bced13e00274191d496589dbfe5fcbdcfd647736bb69b0fb7b99c09484d8ec0fab09ea3fe4197c2cb92fd32513894a8084c2b7b91cd61a1d106b85f7bcb756;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h574c3a05556f7855261a9c88f7802b74a652a4452ef159cf2dbdc5bf5cbdf1468b597a4f58f114335ba231ff18fe0d9cf92533c7631c4e5b6d76b90e50e7165abcf84e46bcc93e3e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee7307d7fdd241e531136b9d0f66d61a5433fc1ade55db46b6970b1cafca00cd9678d5e398099d1eaee9e5091bf3649de25e60ce497bda4c3977bf16e34163a2f51c6c7af3542dde;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd10928cfb3354c373c6e69fe7752c84e141e78df77a554d83414107fc3979fe9e5ddf8229851a3b09e2c0e63894cc38b857d6d329a1fdbfed45cb9eb0f6980963c51a4e94b84693;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15b7ed56f7959ac8c018533dd17266d7ede8f27bf167ba0af1e8abeba55f9be0203feef77f8ec753f3f765d5cb1818dec7a210218a8963cce0ab3088e4a62b5add1ece2ae135115c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2cf2438e772d2e37d25160bf5dc0c591c6278451bec307a2cc6bdaa45b674b879669679bd11216653b73324d58e4392ab1a690309cd4025e609035f05896740bac6a36a676d5e7a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9f5b9a552302eeca136e9e0db00a1ce182609fcb9c4843a30f107c41eaca3195a1ddd746866b2a3163e9fcdf7124d54bc6970b86c73a16491697119a3d4256d1c9e60190dab9bb7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c1485f287d47d80663f42ee251f716b934a679047eebd67d18cc49effd82edfc1799ec252caf1cbfdcad6a864b96fc51b7998f684eefb05a858440608b325cdabd34241bd77df14;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5ac1778a6f508706918bd429d4510fc4256ce056ea3a9b9530606d56a2e34bb3d0cf72b88174bab67285413da47c1b999377a053137ccc610cb31bdcf1555c984093807c7511f5b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd2b2ff3e7932a49d8bca4cf1ea9a3d695e13776900fcef2f078db15651b6ab989fc0ee076fa0a16432bb020a2bf1754e16c76cae4e67feb3e153d898bafa4e4f7c7853ad6f380ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12554e14ff2e98baa5f4a2a1f68144aaac40f22bc2cef00d1a60296639bf4902914389890492b283958a18f0dae772dfaedfd1f00e4a6d6f0572c4d627d1686f59503cb70dae5aa1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e4c8ca2af8deae759ca7d5d57c10ff019390712388bed64648fa99ac929c40b42bc82d2eec17044cad3696da438a3c5be90d8fdd012353f358201ec9b74e4cdb1b8031297fd86c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9128405878e0c92ac6cbec8a62458c994f6e5c665652abf90ef6e74f66e656398cbc546e8cb5f36063e76d3e44d336c6b9aae0a031e0e12a65d855970e615cd43e0d6a64d881606;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e16fac13f2e799fc643a659e207c07eb67d236e5266ebf1057d410df64a8a20c3414645e1ae9c40c559489ea9352dbf586463de582d376439023ba8adc8fd64f4a2ed03b3360be1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc569b57c00b0e942649b2e735005651cebbc2b9fea7692752a9487f84a607b4f3ef0fc00c3b5a3df78065fd524788dcf55b36cdfb06c98d6a59fad888b147266b2a6075895ce57c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef40a4c4417fe6ca973aefca794a6715627ea9e5f379a861d71ff029a68bde6041bd88379287ddfc081edc7b64ecf18d8cd6680403fa27c7ac0374cb0d9404947cbc918a8d2f5c40;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c87b4cb376c1d9727e7f2a15f62b1e8bd3996c2d53a4b9c39d4d5d5392260d79210c5ae3242f29925708dbc37537132ec95818fa6780549dfb0b497ddc29f51eef3a12a613d7f85;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha941e6600600f5039a9875d319ebbef5c9f8c67ffe5155838bee301141bc2000bfef1b987dcda465cf0e81f476b73cda8d83854ca4a048ba96a587000394fe090c9fce1f3cf5ade2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a9373dad1d6b11374f202eb7048e5853e8a494c3992af5a0aa863059eae9d8f0b6ec794dc22eb12e2841de24897a8d5b3612c7fc0a42f06e2af8277ee8700920055c7f82306978a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8cc1bc65d6d2512742d8b5e0fb8740886cd30abba5521861fc97f7ed0e9f3c5204b10bed64ac4da09b96493bf6794bf6709698790a3382d09422a6ec14959b31db9f0e7915159ba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd73513623d03f8c47ce95a2276d6fde979b30494b2b00cffee37c7b0e105a704da6663011a3f684ce2b454c1a700e58cb846ee9b0067381742024d7c089241a1b7c3dd92f960161;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8192674bd48908708b7599dd8e4c82895a74f923bacab8f84829836dd0e0760d6272be3950f6a2927d65757e1c4ae31e475080dd12f133969fdcddf79fac64d12caa04b3ff3b084f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h323bb7dfa2f4f5112060eec8bdd6208162f8ac8ed6212bb44121355fcda2bc1580dd4818e2db13b798c94163dff08792c42c6edb1d3b06253a9184b53747112fa838b9a5475ff4c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1977a644745b38adc517b3d6e92103c5bc6e5947b5167ce18e3dcd3b5a539f71a0c35d2a21ef5dce51ed40b32006c5f3eca60db3450d46a28aa1b41819eb5683d4284798764aca6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdfad2e03f95b518048cdbd0251313e403df1982bad0f7ec044e0f231330c9329a02dcdcad153a01493064bcbc5259d57a54ba9123953a5cbf97fa661606c3a5ed36710903bdd7adb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8f627eca076ac971a2b85fd2692c972ece67c87dbd31ae23a7764c3aeaa22a5f6962e7598ad0317650984f67e8affd4d8d0f537d70213acf52e4ccab541fa3a364c809fa3e22876;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h185624c4edb85b0983fcab6537f5070573d8afb2048c0a117cabc8db6c69977bb370a7ac88b60ca957c25dcbc76281ba45d99bb4888acbdccdf4a6edd99507ef8cd2a5c2a9685780;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbaab17ef090626a67d15526578e7a2755b79a3d8354ca770f977ebe5ae6c5f2794c65acd7b0bced0844627a9a966536589e0612e2371fd98a153e40d3ef6c17b0e5f8442ec410fe4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c5ad218b4c2a1f006e1a117c63f1ecba20a28551ca3ff9614f69a3ca027637cc2344aed577480daa5fb51d9a7e4b0f0c77f425db803b8efd57ede97fca1003535125fcfbbabf3fb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7d4123007429997ff709ed6d2b5a12b6a321c7660b3eefa0bb01b60f429b1f1e42dde9d6f7a10c5d83963aafc40892c014dd437caad9abc30d6ace067c559082b583e7946e90512;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73685b54d666247dbb497759ab3f2a66dc2b17f450d8820fe5d0e38d517afea7f04c6f8c25b7ce5b07c39891fb6d18f485c059cde53736c968d008b38f35ac57e126b97bc2bc4603;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h545dde3b728a7dccc1427309e459e4d1e03e627eda07f05ed32a9fbd544938c99f49af68ec8402a1846a98c15119e65bf188fd2c9744d1233d043a0d020e5c3277902a545be7286b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84fc2dbb2db25a59c2cd5b018c8b9fbc86df914adae9c191c917d5fe4cc22a022a48711c14658e55948ee30cd26bb77ce9dc939138e22b59d907fa2e5bfd7b14ecbca912c9b78660;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61fc0d916df2f76ee5eb40fb89758379bc776724127e3a845da2bba0120189393cb55b9cd852514f36a19c5057062698f68bad01818109d0e4dbe8ad183904493117e4f58f0229b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8fbda0284b9c9fc7f77cad8e4eb2a4bb02183ea235551c1222804ba76b99c15075e572f335985a90b418da2c9964373822f0bc92b63303b34072b4fef57586c873727811fa788ffa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf077ab7027967fb7f6d2edb3559b504764e0639543f5e1ca534ce1a2ec62d813e45fca1c82d94b3a64e1fdcbb1cf9984fdb90be80d194c30d6e24cd094ca737338ea41a871cff42;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e4543763efdae794c0d8523f1d3fe04a4d2851bf5400fe85a982d2a55aee7ce986d27639aef18f786a4a9599d1c3c8ee75b9d91e9735e674d5ec1cd92834a48ab3db8b6274b4869;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b6548dafe7359131a04525deff1713e04b024e2e7bf127b3a1a4773b70f2ae85f6b8ddb845249a2eaa5e190a8e10cb7328b98ce7b9be48a9f2c1653c7d056aee0db9bba8f7b0e89;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7aa4f68e6a57a78b6384fecca8037c9eeae9477210be4d3669d2632ac527bbcb7fd7ac0d93f6e39f3c82b5d2b32746b49150c7facd4d9857d976a919c0d673ee02d4244377d8f46;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f52ef829f3b9337102a74825889964a8864b7e2754741ec1bdcb6c4036a151670e6dce90cbd7b1a566d09aeb3063d2a972fce401adf14428480641f7b3d1d40c91b3f64e1996672;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had50a0004d2b65d4d05e1e1d5836dcc0777f721e52a2b16e572d3cd67f7cd5599933b1cd8b5d2340b0a87b9ee0875556c149a3d43fe2f2dbcad2b89c2cea8309a384843172109225;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc204ede510707650c10b1afd9235a19e1981197418d2901815465a3f691cfb32c1d19e5d14d7960b9eeffca0ba5ef6d898d2353d6a753d141da0df20e0d0a0c600371d5ecf3df567;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9af8896a10c6143a721bc0034a5c1623554cdeb8da6b9a4b8f0644eebe37fec857b50d4c6a7e081ec88641bf983f80df35a487add13f955e6f586a43bee66b70793a5e9609d32979;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b3a36fa1360debd7ca890656b7bfa8097cbe1a3f37f2ce8027ed961ce96f9b2458d428bad3b636b2e16df0d5dd1a37fd2352635f7004a68dceef7ef95dbfad62aae3fc471571628;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c30c68789d513a0a68226b2f6452d70bc44727f934f979c4ed8bc8e1f4dfd1b7f442262e677b609ea1560f36ad19e1e1c3b939cb9760dc4e71d1466725d6842061347a865928d41;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h995214d278394118f079cd5b2b13c5ead3c14cdc377ea4fa6fb104f1c12adb9df14b9c2a3b760a71b365150823efcd5a0231e756726a7750c05c69c3495c81d2ada267aaaf6d7bf1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he426599f0df70ea9bfbfd39ed4bbb5a3624e96977521b29521c8e3f882684872c3d460dd24354308a290b3ba19155b711e123d609dfc704aae132c2c9088df5d1465d57b61c996a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hccf4b353327162aef25bee30dde5c17d07e57f89ce30fc70fe898f3e0baf6f8e1186bd96559e9ced3eba694e0eda2ad999a8e572daa462d2070fd2967a4b207f021108d7438db5d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62382291015d8c85dd2b6013b4ab08928cda1d0f44aa69c9766dd6cc49297a1819f17291aa4c5713840d3150967c455e1389cb354dd78f9a712c43245db89b805e709ac695e219a7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4dd05f154cdc9e18327852782f2fbd90a99c56aea769cbf7b63d3a3a6e6c3639ccf2a3d392df41b0c180f65ecdc6a46d1385eb34db6e79c42e3fbe773fd7f00767da35a0d2bb0fa9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92f5fecf5ba2144d239d826853badf1f94b3ccef8e21c4dad76ef7e5214b1fb631baefd2b2968523081fc390ebce73d71987dfbf8608de2179fd55c460d5d10eb527b501418f9687;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60938080078987b3feb5a56e2984fdc27c7356eff9787d0eb7505c3a543ca24847b973ca6829a013b27ab4ddeed09868c1e7d4270a9f8fe60184ace2bdb634cf325f57b31fd54541;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33aa4b773b60f832372475f82a2874353a30109c7aaf79d305d91d9ffd7df54a0776de61011b82712f6db977468a1dd0164641e30ef63a46be0eedb8c6b108f58f8c2502ef66dc01;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd05babe06a9aa9ee7683190c2b12d940c2a6d350334c807674b4beca48516add0c9799239e96cb49947a3d512cf90a7d5677f70779fae2b204414aa89c397c155d2175bff00faba9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23e893d6a0ec715f688023fca2a1e1276b114949ca023a3a3eef499aeb2c76881e1f49a92604ca8e2e541bba9033d9d69420c12f88ae708bc7c5aa38129bbc8a4dc0bb11f7948d95;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd20ab64bd91d7c6e8ff92d795bc4f6a0b31e02c6ae8f8ca80e143ae602805703634027761c970acf29ef1308a8becb5deb6ed33c3b409c2ce5cf5fcd5ad77daff481bcdd460ce0d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e4989839e2d004e5f4b92f1537e204f13b0229452efb3ab43eb8ebf4306ec765af4f844290163cc4d49e35fd5037325b0c9b922dfb35b0b7e1a638c5b95d3ed0d517a78701c8a8e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdad5fe9f7b6ed1757a3f328f3cf0d115fb4f1ae4e26741470517ac1a51dc483634c3710bcc161c73093e2c8b2aa58619821214ffb717a525c88a8a0559889397d055de7a9e651007;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9811fd8fba8fb3b33a1f12de08c047759d37567ae0fe9f31b18a294f8a5ed2604d27168b3bb6abd2b1e279544d08edbeab8ddff6d4c26c2edb079b16db4f97295fa1d64ae3ec2868;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc414fa0eed00edd6fcaf8d2d512362d404d79b827e1fba036077c40bd93712b034276e4384af789a060f238d9d1870779ed088208edb4ad94ffffef6b7f21e2e13b03473f0bcdffe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc36090414b25738c3de54800f87fce35f19cf90229d81cd3a5533e32852a80b651eaf5045241643d1a15530ac5fbb740fb42194c1a3500ebd5e22a3581b1905679096e6efe529464;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h436bb67ad4dbc71862405b5c00635fe97e70f2df21cab6b1b8a6842541b406dddded454d6f600fc926c598040bbc391c1816414cc0306019f8e248a4700d15b84c279cc0edd0da4e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ff7894dafbb221fd2a15e01a5ba85b81f3f28ad97d85a354b788bbc91f7962b7b7311cf2d68ca555591f4d69739523b862d8c2c03ef8a9a0c0d255161a91110df7b7da955ba8b38;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7c09ceb998750d40c276e0155f426e9e2bf37ed4dea603d557588886d7b6043adae81928ef559c2092fcdc24fc2ff215e5fedbb5f9ec08fcc25272816ae0a969a1bcdff30aa09b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2933515732b25ea5bd4e764c7e5e69c1e3421208994dea5f6a92755adb6533f9fcb26a7259a52bae5b9f1f982a6df1d5eff288f66840e2a2394485d2aa81586b96449d639433d0bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2918dcb7bbf1b29782673b5a2c654dca7b348240b4edcc29d68433f42d7ca515623f51a9bac54fd2dc865a871f241e7128a10e9caa46c4e1c091d0d579ffdf7081975ca876a91a20;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d1a1a1425870e5e546a7106f845da336d37005a9132f4a9387d349a3cb4b6a58984432bdc07140acd00f257daecfe8267d3ee430a9cec3073ce272c46d0cdcc2ad36bb89bc12826;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c2175d5724376d74682936164cdfd02fdd055a6cb5d2eaba6b274fcc5de08f1307d1cbc06a0c90726ea9668ac8a681978959c6876124632c2083a7ca40a6fad79dae66c56de4214;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h134c0d3086068305ec1daf8a973406431f4f632b6e62dc9d4580f2f53c969bdefac26024e9dd3f6d03e37a7cc9c47f1f5276eee5db001dae4d6eda94739bdc50e198aec2300d52df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4dffb65c54b202a5135d491ef3ed1dd11fdefea0215ddafc6ab120424faad8feab0b9fea8c8f21e4a5b35c4807f70db89e1bf1127923f77d5744de129a952ee151412238bea542f8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc88abf75e2a4ae890d8b8eef5c63e24528e19137042d2fb81fc31fe3052e705ec62cdeef950c1af70525acb63ca4f9eb553783cc0797d600a0c255a3bb135b59ac4236e8c29b53af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77db38cd9982c4d3926f04d430c174029ebfa8e75735ec7cc743a4faf313d793c6731362c40d2953cdae21682db11b89c3a2a543a877fd1b72613101611f3f85e9e4a5320646bcb2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h906434cb7a7bdcac98b74a98430b32216e186cc3e2568be7dfd5ba41cb5da3905d7ee9d39376d9127060851bbe31f331a266a962e07dd266bc871688d51b9fef9c899c533d1d9e90;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6d650f38cec17c18b66409c65e6d739a36ac4d1445152d422795627af76eff5f001882c284fc86f7d1d9fe7a23cf68ac813d7d6fa3e8e0f2ab713c5925b6d00d64ea4b831b207e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78cadf62c78e4274c2e929a777f77bbec9b71deecee0d1d97f8af21d84931da2fd20cd49dd76e38ab7521331bdd5667988fbe11cf94c4d4576dd450e98db6c2d92b46e75497c0c64;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1521fa518c946c776b01552f2854e982b400b17df8ae0b3859ccb063cad33c064e172a11447cc6f2016b766a088f2d034d7e774cb32c449071edf112e48b71a2f07e3033336c9dce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h689e9d0c7886568a843c319f3f7a0186845c07dc9315dbbf59dc09f15e23bf1a3c325b6c00c3382f5911f8d5bbd5db4f630fb4884e08dc2b56c6ae58497149022d732c69b8a1a0b2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb550e6e1244db3caeebfbf928ad131692eb196bc1d96e36b627e81aa8b93682649c8daa50f5988656997f4286862b02c7a28baaddc8fb3ab76dfe1efe709b886e6164f5066df2bd4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4e32d08decc3c19a07e25779b5a84b0a2a1f576bd0d9d30c3a1ac3cd6910620a4fc21d5741be92c1a55877223cb5d8f58a738be7e0d4c108076b58581961e648e13f1d57d8fb77f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9ef31481ce5a88445437ef4864381567fbc015be30ea999f42361ea08cd11e310627adebe334735f1b517fe08ba28785e8c29389b3e640e4c70f65526c682d6a75346a255f40015;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51f0b024eacb36473a0a4c2c03ef07484d36e3e29b54f336b9a97d0904f0bf489f3110dbcdb289970f1311c2b81444d32b73b121e9e39b7a9e289eb9d8c07d16ae7bc623c69e0ba9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf202ab76627956b9823da7d67a5dcb5ebccd677ff71123665cf009a8be7af454414b33f17fe0704d56d41dbfb8b4b47b52de52c3e4faee1e7a8c42042f4191eddc3e6c9982b0a04;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2695a907de5fecfc0733b526df048635ca4db73fdf14e3099d0bd2ebc825fe929fde1b0ae6af83fe7b2dd909c5b12911e9365b804ba885dce2007c2c6ed245fac8336c84d2066cf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46562b795707dbcaa289075a4aad26d46f32b8338b0a211a7130e1ea0acd8030fd99a70c9f2faabcceffcccb0db6b45bc1ae823a75b4e0fc3f511526c773d48235db320086939739;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3322b8f992cfbdeb9fed416b5054e52aa1c4056f51c55780d77b4eb9abe8377f1f38b35d921068cb6fc41cc499f402afcac1c4511f0d98c11bb6da26ba1312d2222c5b47f49475b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2bef4f1e99c5335fd77ef56a28ce99ed00d57815e25f9c9dd245957659d1aaa595cc16f86019b3acac2b7abfdc3a3f22ec743821041571b61a47f4c233e38a2ba65799b1442edd38;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab85251b87089442fa4983a09b47a13fd542861e8427a9a28fc096ebaf8a78ea6b962b5201a9d953a9073dc54425c23fd9e0ccdbfe2bf70e9357e4732abe48580db17d75840d9b20;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd652ccaa3225cde6986218958852e78eb0fab7446b5b29deab9822054c00686a589e804701b78cc3d3ec95cbf242ec0754efed4b9c0a37d50f0795977fb610f37031e44efd8e3e79;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5606ef60216a4677c7da4207bd78bf11e8f757be80c8258b7db91a838173312243bbeed2aedf7ded48cfeec52245d94f3ef6ab6e7ae350e5198d8a5890be474ee7f2bd3aef0af4ac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h658c015780ff8e3d66cb3119a470cd039f3a5ce8b3ccafe031ed25421935469865bd167a9aa01658254c932e63ac4b13d722377c6c43285786bade48696ba3deaca2892614c2ae71;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92df866d06c9276f58ae1662f6506c47eb508822e34a6989b581818a119c808a0fd43b5e391d39c22e95ecf6b34ab7775c33a849f556470b4b77cf243ebe8246bb5daecd1dc75c6f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb446590b743732930b3f3594322cc9d29412231c88272c1b46aab5bedc237e154d6b24718c64dd353301abbd21618ab39870bc24a09b51e1705ee6e57c92b21082167276849443cf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c0295b1a7d23ec12ca9ec84735649c13ceb3b343a9c678ecf42f3dea79bf5c5aee6b67f32bfca490291fe04791087197d5ae9ad07545946da2266ad884344f9a8c6b3bc88240055;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a0e36ebe1267d307bcf161b880971a5082987a86413c6d6e2f91f0b57d48de10d4fa703af5cf692cc52d59c3ea5b7064245acfbb65f628225969e4798d5b98ae4d1c7d1af46859;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h724622398719d11cef922754a2db85ac15a796bc34f50626474a9931e45f25192624e93d6874015e5862293efe4fd41936334d58bfbe4de9611d8e67924606d5a6c728395f8b73c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he155cb81ba1ed999099efb9f65102f358a3b35fc167291d3cfa3f50625db6fa447e7ee089bec54a7b59e011feb7f8e94ac58a4f7c1961a8fd6bf5dc77339b16f1c83079829f8cd3c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9d52d9f45ccca97b43c080877914dfdce414dcbb79492ed32f5b2e6e200f46d03b3e9cbb33ce7f263b9353e9461f864ace1b57305f1bf242fe38709c09e443e50ffd7a72612cad3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h804999ecc6ade2968b701744b0ab9dae1b712e1f938725054cce2ba02c68e21aa7e970ca03fd8ab2724c06ccf8b662f5d70f3efefdd7aa5064210d9fb4026eb4b101ed9a761ed4e5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c3a6715d733b1e719400f74f664361057020edf76f8b656ff7c331c43a122a1e3b974525324f4d7836b16a4b61adb7bb655c1616225caceafddc310428e8f77129e93ddcb037d07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc26f2d6fe0c14fac9456d3bee3d61fb71e0542ea319ead97a137fdb0f41d509451f3dd862b6d6bf57d646a54ea7da33327ce6aaa929bcd4956a65e6df0bf29e3663a480882fdb025;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83a7509cfb7d279b16d2eaa7f44ddc499d48b7b5e591eb64f6f890f076b07679e34f7e8095aa010b21d4b03a5a169fc1804a6e40f028008222f51e0046fb6bdf421be657a0401c9a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h999123cd22f978fbab3b46f804edfe8bce4ee451b28d2de76b2cad1189defa99a12ddf99f1589c2360ceebf0dff6f714137aa4e88f31fa9fbf5cbe1b12901a283bd6e99ec9f7a33c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7e867f8e201b137a468f5c32535e8bb3f9cd6844d764cf78e01fff733088df069872cc7305e92821b7fc96c0acf1f7b004d91d614665b78960d6e019f5d31683eb2bcdbaf54a7ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h214823d200bd5490b952b943563dd5b51f25acad0b4a9300f7de10e6158f014f45df00f42cfdfbc48da0d61801e4442d1a4f8ef4d8132893585c97c4ba84064bf53c3cc7e8613cc2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbee2db2df14e5fa5f11c22f8d31983f8607fb266df98f5a802e21775a324cd0488b5a6e4913f3214b824b036a5cc601119e234c0cf561a925f3e9f3ada1355ad782f5e11af8c95c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d95cd3b057989372152fbb4f1bfa76e3c3245aed5547e1267980a915000adba8e558481a5b3e7fa9ee87de211fd76d293b8a5f37973c9bbbf2937ed5a3c4ee52e2102e92091f9b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h598433fc04dd0f251708ebde99b885bbe662f0647b3dac3e93c1d1ce7496322d348028b6629699d6506e2d4b7dde880bbecab8b07cce302fb27c13e4e219d41ac4a32436bf8de54c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he83fead891bb435f346cbb2cdf9b9084593b068c9d7d1ec3b97cd3850ea80b39aadc48a44200992fcc351e0c045e0037784a68edad16c4f94ac8b63f1a5a86e3f72c2c29a6026226;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e07af30f949ff6856c962328853cdec6b5aa05c5727237b126c3896c94c2f910c940043a8438889f82bfc1b3d6642681ef8d8958f0744bcbbb813e7a46d70126ae13b4d3f1c6b41;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3617b60c1cd622df2f0f47b425db54387a10312a95ada305fab461c1dc94c99d68d56930dec619a036044be0482c2a690fb4abe76c4e7d5074663de42065d7c0a48789db688d6fb5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38342f569a496408b1f1fd09ad833c71808a7ebcfad9b77675a96c63f9ed96672dcf35d412ea109b81812ff01b450404e4d4f1367439e0a7d24c04279fddc3ea240bb9d2acf6c393;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea3ee5df196034f8b07590173a63f742a916c23f3c47790958f760bf1fd540ec338b4abf0a983c611ac73bd04c12f8d4c361dbd2d2434dd5e15400b99a7fbbfc8fbc116e24f03057;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb55caf890e9beddf616dc7f7339b6877eb6dedf72845a80a526a24bf13b774324296b25ac51314026a55e7f0a2ece0ab348d43cb5cd87eaa4733e2617906a45ba45580e9f55b976;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e60e5cb4f18d10327a47686d0aab8790c2e1a254cef2657099d591db2723682d7c9babd5f4888113a089a7aef7751a31d9c5443fa153709d67bcddb329a00b6f916cd527483329f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6101d306f6d4d502c95366405b3766cbd9014c1d788b158cf2822cb94cc338d2af192d2af399f299aae4511c5764b843d620e318c2bd8bcdbc4c4d626c1ee674967dd8db6e5fd9ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf28e12a576aae3af791e3dbed456ba98e48d5f5c4e572fd622c386b73bd1faad18543ba1d869c22741a84fdc091d5de11908a34ca8629e90fea53ebcb0a16e10abe366d4b4720361;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8dcc55966b357df44c357ee0fdbdc13c81426772c537b271a4c966f2956c253683970c034d37c4ea9bfd35f92379b2ada326bdf51006333b093f4748ed7bcb01d62ee23fc425bf9d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d7bdcb8331d73f4a4e904a7b50ba7b62497385352c045e3208e846e69d58e667c6526dc7a8b102455883915c484c5a9bea92a4dde82927f66b617a0637351764e95fb26b66d7e2e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a7ebf64440e59d9f12facb0edda680c8af1ccb66484d5d80e7e10112d8cdb4ba80b86a79568e96a07af1940ceb400898b237a5d35734abea36578810e409607f0f068c9f5d08892;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc65dbe8587fac31859b4017cd0416b7257e6178374b16a40e54bed5fb866cfeeba50051b2365af76860861373cd23a4a15fcb8d50d3a49c82328b2375cf0ed53fd8c2cf06e20ecac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f3ef952bbed5b139ada1623784639a2a20c8b51f6fe78c384cd6e7340dd137f53de1a987a0703d2c72f7df3c5e8a99bb8da23d2833c39e1017ca2cac439e2e6252a49b145382060;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h632e6f4ce4f76772787d3c903ec89f319e3ef700d922eb8a94d700d00be0fe7cdbed44e2c4600b9d8a774b6320aaf8992afcba6d6e9dfcc37251814e0d34835f035dd51e910c86c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb375c8a7512fc4d92a8e371a0e7788cca26af9f737781615910fe186ec80d6d30558bd08e46583642b5988243d1d9065e6bcd44528f3599101eaf1d23477b989e1754bc12ed8da8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86750746117bea0c92a151995e4ac630918c7a8f85d86954018c8af0eab6e855ae3d1710329557f01039e08727cb8ead6d8fb7d89f932246cca486f7e61ca81bb0f2b78ac30cc3f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93c83e0b4e6b0a3be235aa2267fa2f2e33cc1744a66aade52dc45c73f440d1b9eaf794c2aebc5dbdefbe5420e2e3734f51d7ff9380499e86cbeebb203ba68f497a6f0ac0c51f6653;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a4498876c7bb6d05869a3c9bc893685ce80a42252a78aa48eec3d96d8a45cc631730f30f4e4587c0f31a6f552349a3a5f82670c1a23ece548dd5920a989ba46db1ecca3467366bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc143fe83e3c1a3a0bf12ab2b83c31470578435883e66aaf71f417a5a280e5047850427920e1146929aa6094c404a8e30c461b2a9ea40b61f80332ffb949f10a375973dd74b529766;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3785f5623894b49338993626f2444b33040e3c700f4aeeb0b2a19db9e214138277a73bdcbfdf1e762bd05e71beab020ff74b99bd501abc17a882e1f8e2c5214a5c8fdfb702defbc5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha80829ee7d2a9b6f2f602c969e109a4da4d7b08dca39afaeec4d4046c31d390d2db04b4b04197c52163f40c2143d350be0a1613e64cd38e15e1137a0c3cebf3f9ec2bb0eb9c76e6c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8fa9e45acfaeeb6c8fc35c0a9805be5cb0fcfc6f851ead1f3adcab96f5c54e1bb659391eb1d8b188ce6a8a9e26e9bcd8e9ad272c986c246af65acebfcfa2117ecdc44e96ba8c7775;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd8d5c80cc58ec95bc79167db779ebb22e49096d91992af76d90ed436656badcd67c3e0da8eaf9f2f1bf5d9f625decc231884d909becc7b5ee9488876c4855fc80988e5cda724328;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h478803510d0d9c08562a17739d4480d07bc32143c6f70315cedca0815114bc86100e7d0673b61b6daf12b06431bec3204987978091e3502849946cbe1f89c7f0c9cd5fa88a013982;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefbcfca7bdbd62721e9b2e65cbe07d3e0599fcdf756fc2042e00c48250dd4efc881183417fc90e9d36b253ae44e2a8149f1ee40b4a55b70b10cea06ae0265e7213b0fafdfa94c57a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h628efce36c31c8f776520b6360c5d14679ec2ab4f4fbf23a03325d87966297feb6effd2b3e2a7fece25a9ecce1a89363d72133a1daf04570c4e9848cf2fc062dced622ab2987cf36;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha18199039a5365b1bd3eb244e29289e53d540bba31dcf67f036e477af4f471743efea4a5f1a025577e35cc9c2c79d07793cf3d659647994e4a47071feb1dc045056e4a3932f3b69;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e7d41646a467be06885b9a5a97b29a40126c6d373a5f06dc2344faf510a5fa59a4e0c6b4fd3198d23cd9e02a2578f2b57c0d299c7c560bc6f404c25533ac5fc238a0fc35cb63d78;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80c5852959a4bd782995136ac816b81f51608840ac8b2960d8c5d7864ceb3dc44ae123437fc937f0d2d6ad03321b8d5e9234d92498563db01e140920534b1d5daf6e46d17a9ea626;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8a4b520f1b2e4c0ee849f1ad8e70ce343c8c952276ecacda0e0c95cdb75ccff4f034b87df065a00aca838cba1a20e6212bd79e45a566025d2ff71d77ef6aba5b39a015c1f12aacf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h237c3b02b47d0064a8fc4d81cde45e55301d1b1f81a0327a75cac75e4c36455e2f5c5f1bd3b7900a4f24a846f5413cb45544eb5ff80215ea714eacc1a4c7ca8152f12611a0c95d39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32f732b74e224c3286248c50730a4b4ec55307849210d16fed2aec3e67c4d796541475e11d385f8eed09002713d976d6b1260473fbb7787a49c649d9956550adfeb65b47d98ad1c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h157b48601c96d4c88a1ff665ac678589d8a8fae596a590e3423e7551ab7212efd97da46087506227cccde91aa1cb8e0275a9f0419e72ab0e4f649b5d03f536d2bf1daaa052c6ee63;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87c4f049a008b0c127782b4bbb6374a30e974869f7ea097d950c15d6fa19b0664d53fe53e7f53fb14af640d25f9c0a9ab78f950b0e5211dca2edcf8be0fd1f5d2fef49d40dff6d50;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9caa18a4a582c63e847a42baea817ebd4dd5492a7cbab8756c1beba08e293e1c86ad7c7c9ba0e073431b4d6bf8d05549b9600985a28d907f8a730437897817d5381407b5b33d26a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h37c88ae5069e84c0a13c3ef14ffd4cf1e58506e0c4139c74e0abe257611ed6f8097e4f1f41d418b7237a321da1b5fce1117bca8ebfcadd3c6ca1e4ac41007e3b0fac796b7a5fe8f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cf9531d2f5f5c4dcf5f42349e825f302e470496af226f36e2ff9634fe92f88a8c43137f7afc901d33caa72df8b7fcb68e7e5c40aa5d414f6f8436e34e04d7fbc59290af6104b0dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28a58884960621332ddbdb0fa3beeadd31869ff106e517c96edcb46cd6fecc5fc37fa030e304fcd48055afe7ece2cf13c25bed080f42a1d5b1d01ae3cabc03fbf5e41294e76d17d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e07415dcb31d8319e76de59ae80c553941d808db96b8fe5eb9a6933fc3a33d6756b32b169439c89b4ead30290e2c266ef66f7c291bc60c20e5599655fca732c6553fa87353e33f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22f27e34cb13cc619eb972c41bdc628d46a22bdf36abe922d7d2ea079e005b323dbf3f3c17d5b720a361111fea37acfd5fcb393d80bc6beed5a7dcd28b9338a7a306de5e104b3d49;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3263b2463cf83e43f981e763318396b0db9cc07323f42910fde9c2ba2d1f69645c2db18a679aac613c795b2ecd87737d67af9984609697baeb82c83a0bf4c5ee60ae99b77f3a5134;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h171622420745f6bdf2bc7d1928656f25db1a40a7998fd8a99d2c5a9c277697c8c57b06bdffee4570c7adb875b9798a5879a143e458cdd21626a3ed9435dd9e2c5600ea9ca9a16fd5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbae9c8a42c5266c1128d221e5d46e2811a83029943a35e4c7432ae413edb8bc3aa3cf2a0ab1f995b1984bd9237a295d68e5abd21326b33037bccc8cf4eacd2abf0a02a4086918151;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha79073be6336c492e01440042109716fbc5575820e79837ab4aa9d66bd9e33d3b311316222b5f4b9ed48e2c2e1259362d531bc02638f60ba9dd1f06a8b95cb061e4bf359b9562fb4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc6d288473bef74079376147b55586f465ef445c6447b46efd228ab1073a754e7b6902d0e527d62678e32b58c59dae285de12f4571f2411f1209b4898a7653965133afb981be16b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81bdef4bfee71196d232cd8ee016641d767b740083b7312c63a228042da418e971af517109e61035ede7d560f7ecdc7e8ec8ecc5fdc5e29d628110f122e3a18e386bdafbb2b59bb5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h796de8c58edd8247d19806049f6dd666aa5987a0d6f9a1fc0ef24f44f2e0fba940a456fdede6853342e3fe33eeffba31a861dd324fc04b6ae49f8998d453ce418155a7564ddbb437;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h751d174c81c92ca76c60d3f8ff49f396d9a4def13fff0e4bf7c13bf8b98e05852945beb72172bb1dd656311754dce9e127ccf883af4b98183de431b55b8b0a7bde15bc36d7ea0a12;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd3fde3547a68bba2c87638be093d83b86e394aca3ce9b310cf27c4caafbabda4166a3e310f853fd2f4442adddb996cf75cdc08c1209370448e2cc17b693ccfb77e8148c9621b34c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6d3bf9ca798c1f073447277b1ba6347e899513dfd8b50b477b11a0987825da6e7c00e180c2dd8a83ff8370f4520fff97323058b09587ce4a1d8ccc33d59096c62ac21ebbdac7dc0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6af652d2e50098614876567551a764a035eda2741a0b2cd9dc2cb302e09bcedb0e24824b667d9544e8f6961a855cba736f92195637a6c39a7c22c99366a7a29cf73128fa56555e6c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee412996abf81e9ea40c69fc28fe6d6ae7b0df4479aa07a0c4fa663f16112a479f8b943edf410843e895f08bee5e69bdf2914bb4928fb18df210a02fe4b28a6be4571d22246d5b5b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22093ba54fd21acf1fa7e6196bbd108492be23105df91d103dcf80295930c8a2e26b19c6dbd78482e889ac0febe8b7e210bd8174f4898b54c27cc8fe117744ce9873e45ff606d04b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43f27d5a0edf5f562b7662166be13ac315075bfefd8cbb77f1b81bfb2f61dc989b432e3830f09768c69900619476fa974d079dc7af4e21f343407cdf4b973742a0169d589b5bf291;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf042bca75dcbe62cf5f049c69787ab3898096048a303c31c4aec7dc79b706524a0d633fbf8a96533306cd555bb1f6c6fd747bd8559d68f9e2d3b24397ea97fffaa1f872940a92676;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d4d8e64ea5b44dffb7ed4b138c5030ebf33820ca3b4dba7c2d9a1805cc3732df5fca6227a4ede1c086e7e97070439fc29f68146f442b977e9aa65cc4867e638250f8c15b01e1311;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7a758c27503a6141798b82017865d2f0ea7cb316e757aed9af9e6495e2955365766ead9a0c6521df0d9927db240d7622101b69c72a0aab702f9a383bf3d62fd17d6fd18782359d6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b34e6e5980fc6e0ef4ea8ecc8c8d800d5d4e518079644d829866097fe416227362b97e1e3fd5977cebe1b38824a37ffedce6c811ee52d22c62a6ce074abf7a7acf4fc4d128fc900;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8aa2d4d61c9eca97d74b58c25dc010164ecafc3602fb295bd76a1968c2157fcc8f763f147b6867b025f4e16be02dd8b2f9aecdb63122c1c02ba59fe80c9f7a01947afc76bec01f22;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he18652690f1649b3bdb675545a0edd80aa75d95a63ff3b043187b9e4461aaf95d59a572f8f16a84ac3855e3b1fdeff0b9ce00360ffbb540a6c30c9815e05c14129c3f4008404c14;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdf08a6d4882ef72d9857eaf181eb75b834adde28a97358e1b34bc256e7e4ba89c0663c8a2ab2aaf9acaeb92ed975b1feb25fe2f663c5b974fc1d08538f15c1e2c2ff79cb95f4701;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1fc12342c3ba3e33839508aaf4f3aa55b1fcd7ca765f2f1a52b08dcded7072ca7f415eb9fad0b1490104217eeeaf132c9acc46c718f7b06f1e1922ec42efdefd75f0a7a8f4b4b55a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ab52a2da2921b7a84d1a1d33e3a68d7d71835012517bcbfc8d0d9eb9602c44f8bc45e530d44f8549bb4f06d94a80f5c1c02867dfff73d6f1494c546c837d174b8e22ecb5a44b00f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7917b887298cda12de85946a0b9117717a8f359a199143f5d012c14fea49cc610f64d1df62311eab554285062f2a447a36cec8213f7209218b55ec72219c934590fe32df697dcef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55415556d6180da30cb6e38a43e300ae3be1ec4b588a860b5d3af15ce2e474d195e0bbbc7ac95a201b6a80ca98c3c2f070f0e25381efc30bcd6da6655d13290f24d0a20f821fae07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5d8dd81376f50024a1b231b3699b2ed23315bd15bdbde60aac195d17d9a787d0ef0df6bf31bdd5c0c7de7969e8b6be9cbd3927f409a2fe6e2fed2562fbd79c55ad42ff3f4fa5cdf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b8b551225dbf63f8c5f4225c9264f8bdcaacf284af03f97bcc82ade00c1ab727072859be4ea407629daee59db366c2f3d23e2b44ce04c76fb41990489a1e2b5daa15e75db32eb6e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71b1cb81bfa1898b4c7e0cd50a43e8423e7737b649ce3b592b8c072d122977b35fd553dba162226d76d0172d8f81aa92e1ec89318d16fd5cff663e9b4bfbde87175b090fe2788a0f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93bdd32412060e4bed33aa77dde46a096057e6fe6d41c778dae0f57ea38a38c555038be5bd34c20be9172cfdbcf510b097c5bc37a6a33b5458d0df6900eb8f2668cfddbdea8d78ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68ed33a9db18c39559731ee48f141cd06f05d1624c9f3febae2424bba742f65b2b3fcd44bf6e12d7fc25fb3485f1122bec606a38dc028c7daff651789171f5ea07b330225e5e2e54;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he19b177e8b4dcfe851c14b599a24eaef4434a24ece75731ea5d8318af1a5bbe08d47f7e82b1d04edb2da565e324b677edf76e21b463bcd7d00d2ed789fdba510d04113615a2aeef4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ae27372ae23fca59a4f91f4137a445d8598a9e2886eb8ceb916a8b133e8ec8d31b8f3a366ee0791bca80106affef01319c44b9f7ea2280b70aac27d2ad5c396a81fc566e1f18772;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecd1f03d458c31b6fd2409c7f6b597a7fb799a721f4d8e22303d2347864284108a97de0ee9be2fcb703ab97ec91203ea3a56c50f2eb61d6727ae07d9aec1fc18c6fbe328396405;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb823e29fec40911f3aaaa1b63c1ac8500c81371c5cbe5f1566c92add00fdd393dc24e3f0ff0b6209a131417b3d02c4b0dfaf8e0cefcc744056abc3c475d70c31bbcb520ff08de82;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf392ba354ee9021aebadeacf6ca4abc642439fb5f01b8e6c778fe253c45321cfbc4009e1950bc2e3305f191fbb92f9a9bd81f211fd39ba4cc8ac9ed3988a1bcacbb9dc5870f3747;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h996cf75d36683886aca3f613dbabd7b54673ebbb2a10aaeae24692bfd4eac71c94756f5c5f22ac7f7c33cb190e1c056f159de3db9a0d52ccd4da3b815d1b691e9c4f0322dc008a25;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67ae71916ba52ded41f77647861fb144d9b06fc643c4d08acaacecef0012804c053b1d4e8fe929c3a5b2fbf0e42d2ad249e83f09738629f44487dbd795f4a3e48b33dfd43fa038e2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f784108cd3a5acf2bd72308d55bb06b8ac1f1aeef6262068b21759d76422ecf0aefb9d35ed595015116593bae1e33faeb5ecb98fe80a47df3477e302b2b886ee783a6101ce4097b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba46665f4cf6d7d921e9e035c44e85462ea8ff3b1e51120727be2fe2cf3be1696762fe2eed25a8022f46c3e20eb6af3575f314c4424eceae9b7cc21303fbecf4e551356effec5f71;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he921b47f9b50d264ab10dbeb7a111caede4cf0c2acf3c800e2c79d043274f1547b66dbd122398b993b87e645fbd0ded2b9a55871d32283b75e720c67f3be089a6656a52b9ecb74b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbbe194101e99eb84d37cf5db915bb28724556e2c7651d675208b99a8be6450e8fdd4745d27a67bd61ec110b8c4aaec770db14dc456efb4ca19e6ece331fce47e9453eed12e60fb4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72e6852edf3f4da43f38d2c58ac96a180a740f1dd7979d54fddc588b663111017cff1db8f485df0d716caeb12e0c8b61c48340303991e0660ac57ecf822e0c7b80167338012eefb9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cdf9ea2a8dd08b6cc0e925c2cfcbbe4dc3f688985961c256a811f29a58f30b9700bdebe996421579f40a897037340cb9ab4f8b180fadc3cc845ee48c7f17f81edffbd547f4f2102;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90cdc83736691f7acd0a526a37c25513a3110e9d0dd8704977fc0b087d8f3a923f4d4a46ad46acabc176bd5ba9ec296b3af28ccfc4f455d29aee01d1949165a08f5e5e0a833a05a0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ff438a73f1c970178897d78d4f9837d0a5c0168e1aefb9d9faae65796dfa305c350045bb37f39726d5fdeafedbb200a58b089ca5b7515961ce4964c09df204f94a4679ee948d87c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca5e6ac007cb24aaba8834b51ec578085ede4e0e26546625970b722dc2eebc1b91c06ccf51117f60becfa4e779f378f27e4fbcee36cb9b2aaea6695ff1d8994d61c810f87b1b68ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8da3bcc72a4e58a6e1c0b8ca7447122813b0677ab5bcdf39fb07a469545e501db0c506b5e6c7ea558289e86fa153baa4dc2fc92e4571348112c69a9a53ec6fec8a1fb1e6ff301bd5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6a650adb5bb4fa4d9bd1e53181dc621df00cddcad4b186a62c51a2c51ac6737da475f80e5d267e65a3083c73febbd857920e0747f3293cfc0dfdf391afc37b17c27ee95d3332cbd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cf8e2dd6b7a558d85201fd3638a5c6b8a6bb74179409af697066594811c5f04eac81bb081f745a754a78c773e33afcef43cde1df880bfba545af3037ae02e8a2f4ef077a1498e87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6afcf2a881a7c3d632b4207a4e47a12ff4c8fa7b405ab394de223cce4075608baaf8d580de947de70e24a573b561d06245026ce13d0520048abaf15aa48e588048aea5322338f005;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9ac756747c0e152786132284ecd900bbde11032267544b183796f3fc51c49454000468da3c69fd4582ac1767c9078f4457ffd51810d4581587cfc0467c7cdd0c1945e8187757bd3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9cebe4570c6c846c8d9591f8e6f31e2bc25c0d4b82f92e985882dbe336d9af915739fc2cdb78264b2a90cab3e55efff8bbabb38b9ef283549a037b47fc45bc583cce2036a6797205;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f460b2e6705a5b13b8e9cb3120f9e41e1c099ce9709f3890f8e40900bcc93da027ecb61c9497c2c0d33d30d242ca038a98fab5a996fa0b36b73c6a1d0751d50b0b7841c2b70dfbb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd36b700e0a8bf3fca4e1b929652dbad70b4d3ebfc1ae40b08dfc921a446243a305e173becc2e13ad4b1a10c3c4230199874cd38553e12f962f199dc6217e096ce4a003315bf7b9cf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ae00a58f0bfb6cb6b5abe49219306a1b914973854b05a75aff8c58cc9c1aa84cdae087d074e7c2c8205ee309d0eee3987b3dae79f41b8d7554b0dcf5c682ca357dd9af5c58f6044;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ba1d18ce6ab62455797e1fbd06c141fd418d22370ad917065dab2c7982c4734e62909a4d92c9602edd956dcb898012b6f69f0f55c5dd4d1182ea9935d73804ab3ffe134cc63e19a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbcca93f5b4ac743a656c9f2bf921c269914b316ca59ac159239a01c5a69f6a55f9e16a375c9c7d9e0c484b792d69fa64e4df1f76f001b94aac6e105c6eceadeb689f0e47844bd12;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4756623a874462e0a1b347e235f7f21931ce98b95f04ef85087de19a2ca6ce474d3a8fbd662b5ad7901440600b0ee9fc2c201d2305de07409b27bd6530de5de7c832365c83dee3c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b124599652adb06d265a8681a4fc281356bfd6381cfe88e4017002bf80e96f8f378653a63f7571af860ced4c0270b88bed6fc1a21e13a6e3aac33bc6ae7c4f544842c2e64fce14f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7ea3122144ae274cd1cb487a992f1b74c818bbe1520d7ed93ade744e47b3b81846fb9fee6ab5578c0cd8f12215b509eadcc6f88bbfd3ab5cfb9eb72a51ba5bf470f7a3d5deb2ebe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77756911949c76548f8ae49ce8f2e7d85863bfdc5188ce10f2fa4f7a52cd925f459dd5353ded4f578bc03164a3252953318f4946cf32889c4ded453a78cec55f3d6eb31362ff8ee1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2fd156291941f97a9a0c11dbb32b145b5cd072266c46cfc9ad855a8062d8855d0ac2fd73a84c3b938c4f7e1f6bceba0a960565519165b606ebe5d5956c3bfd2673be3d3df98ab77f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e62d160128a0c403c4d91dc0c42dc8b3a8d7c71461273f3401a1fb4642cf019e11b8de1a60cb9d6b6b8699f2743bf1dc598a07d7265ea74daedac02d4e75b0d90d683d6a6e25e7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6d792c0ff89903f68b0a2c6df1c64eac113dce298e6d2f96ab6bf3d518e4c4ec2f5311e33b2b253bd587d28f2a3ea1b20070e930265c26dfb9d6d8bf9360312d0e10fd06f063946;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15378ce453dc9ede6b2c14a42b93ebd7c0f237df51af718a947f41487a7f53c7a2a30322cf837ce3403ef70df3d1385a20d0f837d6d7133a7a85e90852e49ee15f2989b33c719385;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51c775b63c62935eb377c094faeb9c4b388c2a1e8204f89d7eb7e50a0f41d25115f67adcdd02b0924581725df71366e6bd4594c327dcd6ce55dcf1f67af193d09d7ad307e221a539;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3591570ae625ff7a72e52718f7de2ac048db496d7366422e9f3093972bece3263b46696838d36e82712bcb415dc5bcc5848a00c42202d5accc47901ddaf325cd9407193e28a7e5ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8de3c347d220a6623bec7ec0d21bed864eadc6905878c6e70f010d2bfbf5b922e1a1746b2ff57709ed1333cbbc0bfc5996643a4e92d4bb2b4a33867918f62b9074f7a59150445ddb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71a35c97384f6f314d195687d5c19abcccf39ccc09e807042d6f2b217872e169d87f9b158b70a1a9641ea0c56029d54b8e9778c95d18a6956dd77405f9bf5901bbfdab7e6498f6bf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8dbdf1c0d014e667b87400ea48336569cd67c4439d54318c621676f21ae62923c9a9f56ac17c3cc7305ca917842c82730157ee74346215b1ed863713ffb63f59498cfa175d880871;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70e2f96fca30b4e2fdd9f6bdebc6386fef525f56ecf5415a61bd292d3e187f58015634a364485189f285a1dfd68dac8a73b254810e793261bc0e55ecede301e7cb6b5360f42c6085;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a9bdb4eddaf836de8424bd9b755e5034666c4a264f67e15ecf80e794708487a447896ff393a6aa1c6d450477da338123d38500f4072c94f7abda49283effc04d67c23b82c690b22;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95395ef335614519eb6823eec9314d1b017347bb9e2323c3d27e94772263e62d819f645a24446e1011a0b70d2f91b4d19972d29fc3f10764ec458c2acc46cfb7084a7bd82d8a9b75;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3094ff2943fb8555bde6d1fb2817c3015aa229c7a000b8e080ba6c070a2949009e5043c5c6b936fde680377d5b5e45a733106c2a3df1c3344cdb7b8cd81210e27090b27afa01d4a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbab21607b574fca8a5a91b245055e4c3f805d86c33865c52048e6d4386cc24b4cc0e4442a84e252e2290c9c0c6cf1e203b9251cb61c4e0ff309cf96534ab1230b2731ffc85f565a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he43eadca4cbf00add458fa091f9eab3a908e143a99d0ed9fce39fbf054e150427e5368ae84f23f8ed687526080ab606a4e6023f3a3fb6efc87ade253473102d14491e8941a30d987;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h906475c8245fdfd3312ae446d1197f95a6a2339af794a6a4a8e80fd5f2574f5652eeaaca7ad52905d0c0850efc81400bb10c5645493c343d7d8d02f7fb84973d78a3790705581295;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf2f2072693920da07997fecaf993cfc35fd093e59888d1422464ffde8b8d95c4eb50a1258886c4eda226b817ea28299d18fcec76dce7e4c0af199d0ce95fcfd154e65e903515f71;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8209c75831b9aa13a7ba5208e8eb296b1054d2e8c699305ddbb59e3d331179ab94ae2ab321419997b723febf9db78c34b839956c92be6667a460dd57c4bc0504c980653f22bf59a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heef6bbc632fa03e590850f9c381367a783b0547d3fd5c1f7ba870a5ba35e20cde60380402d9d48eec2f644fd212f455ca03ffa237ba5e36febc112143c75153f62e49cdd5a3e6580;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf044888b02b26d4ac3d6363bf2a3a6dcc883d652c7d33b8b1deff1a418208719218ecf1f430185c31a966b26e2cf0120b4b8751b578e4f3d85267130345d845866d70cc9c17c10a4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h395e6d0a2ea2633ab03872499ea33fda32d5007517e0de3665dbc63927954c85befbe5d5c2b351804bd3bcd551d8d24846b2d4dcca271ee1b5246bbd71e727133aa6f37d048e6972;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h738d5a6ae11b37c3ea96fed7986e173b3772034a2601e55cc250100d2a30b80e289ed3d8c3126491052340f099c9900c95cff08136464609b98a8d3f430f964f02416564816a3dd3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64061d2decd5dc401ee9a042dbd799065768cb1dfc91e0c606ec65ad646a2d74a093bdd4aaf42cd709ced9025f0d8e79aa92340036cf825adc0056d9133e08d09d48f28c3d86691f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h742083be7af3a2dad9e98a0c72b720db85f3ed8cd9d52c29ad30238c3f48a7da97fc5227bbcc5c0465e0cfb147bfb5a0aafaa4b06e44f6108fc1008de5cf323c22b16209c30a3596;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbd6caee855f9f356ccc20785bd51715f28acc69cb4bac041d3962c193812c36e70516b39e0ed9c1c2679e211b93067de653d5f40f0f15ae7ec9959202247e5eb0684f62d3b5d347;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedc153ee2e9fdc15163fec11248c6c41904a8db584bba58c571683667e63c56fbb13be1639bb675551f396b93a49af71cf0dd67115472d3e4ee3ee07c3afd9c9ae13e82547ace792;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcf97f287852a993ff4db4fe549aa6158c9e5bb4fb60e5c005d59942154971c2a18f83084b9b758afde3594e60bc6e87fb6778636b45d643ec6aa9e5871dcfa2ad5c9d1abab6c308;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16fe50576307a7c171df3ba2d5f99656a024fee8602cefff223b89c43525121f7e75664b531021200e759c80208c690e93b797d9aa1257b0829c334fca0fca61276657ba84862273;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d60a39e18c4e5854a94c3ea752f92f894cc21c3b951b5f867738908771f65cc76c2d3cf6173cabdaf135767c69e222b0a9ba0815f65bbf779b4348b75659ed505b9d69ff47ba19f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10fd11243580256063f925faa84285c7bce8b35fe78cd38d43f88de217425210b4785941ffeabf9185d21699fc7591787f314e9504c7f30d53b76e90b26121d7cb6c07867c9e1951;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5623b98e2ef34374f08473552f0cfd242fe6bf72695c448d6e7af2841f1ff6a9ac344ee9298a3cb2912dd35dc9c9271bbb03db20b5780336874aafa68f302d593d02d874a65037d6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb403e12892d981430b3bb7e4e4c2e36dff3b56cc5f1c512c0d2d418e3f5199774fa41b889a42f0f0de6b16751b7eb2532ceee2e8cb3b5e4d655455c5d4d21803577c68efe971cfc2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h848d362b3ed78e3359f57da0f46697552d8a0624c33311595495a6eb7da858a173e33b35a45ce7090a366881427238cf07572682697e589970ad22d2d406213fb4bd464e099dd53d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0b8862b4870c63b96246120d28489e8834ae7ab317b547bfb93efec9a04eccaba5006f73ae1f583ffa35b31ca4bb83262d2815b3509c787cb40b6b3cb5a6b67d2d6a240b41be66f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c975fdb1bf80383f718d1440b1c1ce8a66e7f57b707475e9ae1dd1a5cd180caf9a282ff7742825f82ac8cf67d742af8b505845bfaa24a44f6022e3283ac3f4f05d90afbb0dcb6d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb6eff8a24b7199ecfff2d3b009529a4f45dbe627e27216c571ae76f6fab67657289fafce8fdc2ca7dfd534df0af805a2e4270b8e5f3733bf32b8d6ee4e53f7ea089e6b7885b24fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb6ca9472ff7ac11b83266ac45f8557701772fdaf6d64b83a7f05e2acacbaa40069015b20d70bebab25609d8390982485169131d4ee3ddb885edf5ed29f519ff69e3380f46e154c3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a88745048f10b4a91a8ba20a2ac5a53076755947d5a9e3ef5d240ce9d1d5c4f52099e2b4fbd4c24e0effb5846d33340d3f1d1d1746b8d123e0ffe45b67d0a93dfb3fdca13cf567c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ad57c048155984680f95991f2d4c5459b3c5f96c2824a69f7a305ba4005d71dd9885743daa3fda78ed13491abb4a78adc7167e6af7d082f929951b0c6426ef6a3f193b2c566d8ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a0af5eb1ddfe572b4917674ac78ad730a25c0eaaef3245408b9277efdf79d6b47a87474da48aaee54935801060f0f26d4f0479db01ee04c980967d5fabcd4bdb42290f1ed44fa2f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8be11e1a3353599b8bfd5d23227e278f433e7f8d9217dde5710d091608bb4a1572a5a163c909b9c87c0d6cae74919e9f395040e3af5bad0ed74f4a295b0b40a6cc8f49a46b822a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ea008a8fbafbf5435bfb88d437a8c47f1d28e412adc2ad707f11811131a8992f4b2b987c061b83ffd8a9f5df814b1d907b74d150f2b26a3d0cc417fafe83f66174962fec06a9a29;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e0ab7cda5834426fb81413b3267a3b816748c0912bca5f12d2838d151bde8250ff9a761d2e94d21d3195ea9f6bd644110b851a064167e34a4826fe844ea1f056fb9b953942c3e2f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h267997e89cacfc8608ba1539f0a2c240e17d77a65f1922bb459e900cf7745bc68ef484960ed0d63d19bad0d474853ae90e49017b7efc615f5cdee40dd2e134205924248fb26e7010;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h392e7819ca8a63868278d25b9085c163dba84631940f328cfa1213d08e388fcbf041d19067aa447c08f19386b30295437f0d42ffe6cb584c0dbb3efa498857c7db043a4c36300c25;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3346949d74330c38e9dc11fb503b053aa76aba8a186a2dc586ba6f2618b3c35f2a0d0515f1a21fe3cd5a14fb120f98fb97043da415635cdf68b9821b41cd11e3c80d9c4d6c9dcca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd83e78ad46768deb988af5765092fbb9dc1bf3dae02f0ed3e56e9c5a8c4b701e96dd45261fc42b1392b0366188e23f7cef8b061ac15931da378b0b00989881ac43d67c4c879064b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb907a5d81c270ddfa976bedd3d8c033542be995bf857b010d502c209c70e10b41c864bcfa45200aa370463316431f1c7773fe3a88c31a3e81c79358f4a94fc968f292e91e4fb0130;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd86927b14a0f9ffc1b5b661106040807aa02876be330f075a87e24b2b9ff7f5732117f021aae6c90c9227bde2a6fc1c37d11d811a85685ba57fdccc57b7eaae3077c5859a10f85ca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7dab72e082d518d661e7d07475337720286c594b08b3928b1648b3181cf2c3f4da4543aad0ab7dc877f4474fcc5ff539d453ce97547b9c10ebf613119f88e0270403ca10ddc5279;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23d9625e157cd742c25c7d9b48e48d832c32276211ad9de4bcae5d395824c128da90d456b7522d7452631f1d95dd4c855cdbb1f2c5434a6c4dcb18681cbe8463df6acb3f45a2178;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h652f42bde5f5849cc63f655727387f7ee0a819d973227f172bf33e6c50f7a852f290123fa1b6704ef7fccc61e528a3411c4032a9fa98446408b2f796a2d1ff22f57555333b039c3d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d9ee373fc29949d2cedd8590418a87ff95f079e87442f6c360ba541515f1525e1d6d2461257bf6f910fc5bbd22fae317957c70964e129a47bb6333ad91880d1c5996f1a79bdf102;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf27b5274dc3face0ee0caf2c52c2cc70271c21fb19a4462c35fc508c6791bd2c4950fda247fa22143fd9520057016dc320dbf3dd0be2de3a7df9b46b4f6af740a323fad682730d8f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64780180e32513bd2848cdec4059493a29105378aa30ffe7d968c0dc2a0c118b35879471affdd11fa5291eea923f09aa8a1d2a6184a4a3393ede1b44bfcdfcec140092eec9e77c5c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h658d9eba9adc0ec62d8efbd2a07d4c0055af3023df6830c73c83cbc949821e8955a79242f830ae58fd331b1c1f066be7ad6aef89e46d0c7485eced32778cd7156d935d3be5b787eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a60fd8471da455b6865a1e9f7cf7d6bd00fa3bde4c5d1840e8ce3bec49f43fe7b575a7594c09a0e6d8ada1cd140f7755696585e44ff8ec0c23676cfb11e71aa68a406a8c4cafc7b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he89cb63115de941cefa0de8f1d47d3882f1f88d7abff5c70d708da18378266682b4f9e5f80702cd21fa4d01f616a109724b6b48ff093abd7b5d2443379501e8071469dfdbc96b06a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ce5348222025b1e1203b70d83e93b5f1a813d0f7cac171cf5012a69543450a59f7a02747b6914393e181cc83ebe904bd95c2fbcae8e1cd53ef5f6935122e72ffe8132f2a1c90e15;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b90d056dea2855ccebd399bfac74bc14356766455484a0729902ae2581384b795865f64a891850badf1d39ab0ab14f860f388f9abfb1144c8d3b522557dd7d233a0597166c91340;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha655a9a0e51e81a4970e459a774daa7e2041b2607287690df7cf55aabe4e82f9c0fc11fcf61c31f8169b702f895712b38dbaf29e6e8a88a5e63df72998010730f6bda6a7c7320691;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf04935c2fd9245746db2d3ed527054fac73871c0f1627d5c81ba78760a84591f84058f3dca72d30604eb5db6dbf2519cbbafbae410f9d19c4d4d112d335c5c9de9cb975797489ee7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85f14ae3adcec5a86021ce0aff6db8f3ef36707b867b654434d2b742c5b957a6a322088cef4176fc1c2901bd79145d7764b33683fd58b0cec741a0e21930034d4782edc1a91ba166;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fedebb20a59781475061af2357a03e9f169ee1b7ae4ca0cc43fda7c1e108293d590d5982b0066f4e1178e8ce279c05ff455fe9dcfd92720f1342a18fca4c4c2f71930ab4fc6230e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6e91dcf97297f9020a30b1efde10c0f787e11454d7262abd718d56631f3462824115607848cf8d47f6d4091270dba1f529968f6f09f66c0cbf366beb0f7515c6e52c47326bb63e3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdd4946add0d3cb6210c31f2b4076a3e050983ae5ee984c4520a68e1563b69e0bbbd9d4d145e238405d3aa737d7645137b86fd6cab8e557b15191b447a410d562abfa7f48a2353d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4bf7954a5354dad58da8c9c3c8ef4257bc8610c232ff28bd87742341a492401b0fd24a56aac3d374ab459a4d3188bfe14bf1fa7806a607038afc36249f1dbedf1161efeec65bc072;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc70344b9a6da7b0e0f30f2f5fe7350a719e75cfe223332c8248f668f120c7526b50003154a92483dbf0a515a9d00176e1c86d3ad85c9e6a73d5920157e5cc7a7f70d1bdb5851c736;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b8fbab58a630b2f197c6bf8a1f43e125394f2a69cd87a32f752bbd9e8e2d8f384fda012bd804b59da7f09f8db87fd4bb8f3cb7c3ffdf03f1129feb4c2c81f34e0575cca9cfc7c52;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42b392d632ad5ba9dedce31be4e36b0375fa9880c74a6229a313299536a032ec8d0e8a34efd760190232659e1b135766f8c4c0b9539159021e78cf26fed8fa7f23218f58c1e3bea2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16bccf42c2de77d5c5cc09eb95f5ac7dc8e8d3463cc5c89fd978c158763849118b3e92053d38b6f2e60e0ef82827a87e7becc825efecac42bb1208e969d8e5a92f5da1bf95fa356b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26121796b50b4a7410b9952444e336decaf1166a3df5b0c5effe38552f96e5644393ec7bd54c5e71674c32127104c88a4b1cfee5d86d0c6210ba64e536df3aa3288dcaa546691c64;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5489cdb16ecc443f7783bc77316311d30f199e49045f541dc2121b07c6288c3e6f5e276e62679b3de5ce14c5ea2935840c43f2a312769b4d7647f9f04835a19c67b01a55f2fda68c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3833c1b7d09002fb4edabfcd403ac096e6d237608308ca46fb6f0a14f82c40f4b410100c87a6bab151b86ad66177794c8217107de83f5a5bf8fec8fca7fe50d8b080d8e7a3b0fe01;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefc663bd7e60b768974ca3b562ea62cbc25122bcb4ef0f0bdcc567a53690c06bfdba8fb8461953e8d804e83df90d57fad3427683c5fe96d5754e9e90f14ee225f9d4eca8bd4ac84d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9ded979a0f50b825baae909fd01b2f5f3f7b7db3f81131871cad70f85c4e4b2f91c005d31078cedced05ec53497f7aaf95615a20c1a603f21d41db43bbcf0a5fd14aeb911abc5c1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11d6e74a53835c71c1a510a1443e5c4d1f2bf85c966ef5c2572230255044af22dfd384909b61a1fcb29d34c4241e1c9cfd4e33c36de59a87fa70d81c503020782dbdcce8f417d3c1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h334ef9f7b3016c2766995bbe77c174fb9e0ea171ac7b3a191d5f7faa10df7f0d490f0e89592949a3779cd2278323aa5bfde51515aa7594516d40631b686e19585651da1e6ae2a840;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2801bbbbc250a97fdb2058ced436bf99efbfced6bf12cd518edc787a6291c091cce96c4216af8c68ef725dc1739d2200d0cd5a75d8ea128fc0760a46c9007a7a444f56ba4ab4643b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb75b05fdb749c3ff6d5e5fea9e4fad9febc983668648720509b50340e33bf2dc43e9c216385cdd743d4d6cc55701da326cc4ad7164cd87e8edd466aee008a4f4160ecd0e6f29f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he25943e3e1345632bfb6037bde7d4e5d1d34b758a4887382bf8042c9419f4a68020c142cad4229d5d6e0feafcbee1ec5ac57da9be1429450a3f54473d1605bbbbf6c7069144d6825;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb963ec3ab5eddd5b4ed77cb8b5b631fe2daf46540033934087f99b39fcc6f2ff99e87716607c39b0379bf8c80f1257d09fce7af96502bcc89e102ffee9c181281f658a9432c9edba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda7fa312fbd9047b1f4cc46e053d69deb39cb89c626c4764b5fe9c57e3514330012a18713145400608bacfffcbbdee6518125ac2cca6884bd0140e23b0ff7463232592ff00de8a4a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h956b3998621f20a04ee31f0d95e419ed71568add51022c2f482b45561882802a916c39fb1cb6df8af68569e585905a250a9f6266e6310a087758e190e7bba155edacad90852a2a58;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53a1e50b4ef95e769e269f2e5360d7ba35ef753256af07e68cf57c89fd8e7b475f4fc52ae2adb7bb00974ace1f3d2b49f5fb25f6af0a6e32b764af781378535609160a1d8cd97723;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76ad222f1abea8828627e8ea0bac3e6524276f81a2b32a6f6e5be7f941c6dc6c5f0cdbe78691e0c769aadac9fc6c081fd70fb78cf76bb3a1f13759cc0aec459b1e3ea6d0169b29f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36d6fbce3c49b50b26b92ebfda2ec900ada7ab5cc72460c70a69efb3b6f12bf1fc728bede8ad34a52f86662d767e0b23469cdbe22501e649a7537d7cec9ba5dbcbb1e06b483cce16;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd08eb49e3d683264d40a37a3fcccaacb9da72f5f10df815ab2c07951f69cfd02ea33f1d527b9b746bedf913df969b4dc99cd44cd7fb32e336e45d831ebe18dcf2e255a6e72486b06;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84ba5fcb3f4a0626358445ba1d9230d753ffc4b2f2d6ba0d96e5b99729b05a7c5c99134f7df4bdea822bdc8e7fb54d82cd1ae726587664734ac29fc7a41bef3ac90cb6ab0b664a87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3b6d2dbf3efbdfc8c0537ba8195f0d1b9efef95c5bc0b6cf12b8eb0cb2e0763da87b5b26d01892c8f1f80daf0d3de6a2465683ffe9952bea1e2212e3b650d4d574c13608e406b73;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h489f99579f44b9318000d7072ff97cf9bcdc3bd1065cd23c36bf67c8ab8f05bf870e009a175db04bb1a31e934bd2df56194001086b1fca33b57ac9858aa78160d82b552a13e84a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf28efadc80ed60d34ea33443e0b6684f54ae9b7f8325c34e0096813cfabbfc9bcfc229f2cd29524850d1de8ce7130aed65ce15bf512007de2669d896a16963a5d6ede23d2ba3ff02;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h380bef335ad052ab19590ab91c9ab811516c57431a2c936d088a44dc84842c8c96d98e112f3bcb3d9200cde0e034b7a14d925c3bcbd5b41f774e1256363cb6ac624226aa4f45226d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc872d04db9d40faf65a16eb9f0591faa26f8b2a567c01fea268e0100fe48a020bbf3f054068883620ce6f2ba2cecdbb1a85b7be40cddf1d09e6799c38b36463906112370e6d63a3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9fdbcce082aaae393e580a50120fa8865c9771de246a678690ef27236334fa5326358286233bf02f647001a33e70b8d01895ea1a9724410b76f9dc23ae81dac826dbfe83f4afba34;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b5ed8559b8413c1eda2501df7ecba16b163634873e8e5d4c8ea38732f2d041c0571d06067183fc4ce3a300c6bb95d4dc9362c6af26463626844829488efb48380f63add976dafb8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e4aa6c8ba988a76cc26162ca7a182874a025751717b98f58601f1cc21559064838b4ad4daa429fba8eb15ec61dd5e0830743ca3cd59ead1a3a8ee7e1c51cd878983f0d8fbeebf7d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h679779e2d561c1bbbf97c6cd3f92ab60704c8fdcfe3d59ceee53adfdf828a7346594df97b9691d5b2d8c0733ab370183fd4614022b5ac9d7ebe90f072052289b9c01f226d3c4ed46;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd94501aa21d511f8659c3cbe8b163a26824f2fd97a81a5d9550c8e2165fa85ce4c9137dc3f67f285aa84b5b9ed251176285dd74f6f7ca00d3911c2b6972af7cfb514b78ac4fcd44;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e4b919cdbe13d8a6f27bfb1472a0c2f533a2a9ea17f9ae214f62de3d3644430f7556a4aa6cd17f1504dd9d268e255e526fef4e992b3de31d1666235902d72299ae0444da43ff32e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46613dd8eb7830e0be7e44bdab722f31b086d5bdf3a7e207b87972db96a8f6f5564fd64fd658a6c0715ea7b7a694c61a8c00af90f1d49131de1e86bfa5399014418a7235c8a439ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c6d983652d54075f06ed0a564c9b4f171484c931a8d0006bb124986e205a63a74a8e609c9454ae7664e366266a1cb5d333ca0027964570429d2c3b79115e89a998ddc4e0d494790;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4004d446b400f90c2ce13bb39ccccd0ff813766365b2e5d1c93d402df9729a765fab658e42c974b54c310f9f482841280c5665bf27d7d5c86e8fda63e52f2f365da969dd6ed29358;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7bf68f9e22fe7cd527714de7cce64499303f6e7494f6b2f590f098649be2bb97e490b1263a71a7b47e03f0eea4454d19a6f14fc19bbebedd5fbeaa3d73e7ac66a498a151fdfdea9c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h981d7f7d795777ea11e800f5e12cfc2acd26f9bad79029eb8d4dd36d1a983a13dbae65eeb1af46a1b8d7afcef0655689600ece4c80f8c94d9e4e52e42934a3425e6c1dfc4ec2c47f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48adb852cb5b372f68314f0a3108e76098d87e224487f843de5856d9b22cabde840360577e741af744b5c9e8ec2728d73c1626477f5caeab6b60e9147aac9d81646ca1b85bfe31b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76991e80dfa831e4884a4e24c56ade555102ea1ca62a603d47cea8d9e800c7a5366939268e4d341d90285b6b3b18f4aa2ef20d1f992433aaa35abeec529a0d8f6a8e83d9429442cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he61e0d2901ad6c5dffcf535ba5d69b568f56acf0a214ba7f984612d292302936e2021e4c038ad8c24f39b50d91b847ab17382c80bd9a225239fe730ff61eb6baca941d3e57b1ed8f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he982987328052cc764607ba09db8eb838ce6b5b397a6b756b3cf3e61e16b859208c9110b6ad0baa57e06d70aaceff6842fb9cd66f2b999ee93e96cc7de44c7347e61c1738d056a46;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fd590a16a973911114b196d247b1cb894d01b05de12523094392d71374a83d129df27dde84054284b4e704db5f558cc866ad981bfb8b52a9b13470f5cbf842befe9d90acf22404a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d26278ce60b570ab26c46f71890333e6dfc614cc07ab1eaa4b588953224de239ab452c9ab884b978c4ed85552638d5e42409c75d211a7dd46945a13db06a47bf694fcac1f71a3ac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11b038bc856b008641d5396c3530362841a0d13bb2f0fa4896bf913487a67fd8b797f5d186fbad508cb13c3de0b962b9f4f70f63cd45d74437d5d174b62554be9c980b8853f5b87b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ec71b53ec5a0eaaed2c3a3c60c918d3c59ad7f3ec81ce27aa4dc61ab82953e96a88ccfbde27d0a26dfee2e61fec94d30ee4f6e49c1b33daaff6a67334bdd9d3211d03fcb89c3563;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c67e758bb5fac006c05ca2c3b9fcc06c22395e17d39bd3b1c0717de6c6071ea969d2ce15c1a56cb03d62f3ba5aa9c019e6ebd35eccafe4477a04e844fa5b47c979f99b28b1b2323;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3be99c94c3c284c9ce13183b0beae72d8ac9ecd4b9854a598e73d7da2c9c5821f5e2f20b17d2e504c7cfa0a33256f35111ea65aa07699f2f061fe1ce87d193eecfdfa3a95f14cdd9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9546aea1a5cdcdd5f760c7c3803907fe63a865bac300faa45d062abb21ecd101547eb0f5fb8da6e6bf06b718aebe9b83a9dae0812f2099debbfdf520a4556cef5000a03650c43859;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf3e3a65ae22faee2c74333013ac85a5ca9a5089e5558ed7d78d2926f30eaf20972795f17cad929641b0a667f109d8b63320d42af27c783e23b753f42867525250c727eb9d212aaa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5018d4f9be03faaa867c657518d059b0d0fc52551242be55fbe2cd408ec6c49e8a599abc82de505293419c06aeb165e6aa4b2c70dc8798e0e2fa1f72538f66e4135ef9a5e4c316f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e7477ab4c75e116daf4b5638ad49f2943c5b1ab2e911df2208f8f8bd85773f1062e450212a70714cc430aa422c01fb553fa04e006ff588b66c9d464adb191a2bc96710afadb9c97;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdab6ec9834261eb0a8b44ae06b736139c6383228bceb9c31057655984acb2d7e3d407e63ab491520ce9ae516f446b89d3c84d8da81d7700bc4422c4ff3c20d73e16d860c942dcba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h114a2c416cf3998becf83b53bde3d6866c1868c58510e2a5b07715b50c3995de0bd3b001c5257c4a6e92665661e5c09b60f9b88f8236c7a3d55ecdffa9f6aad29fdbe849ad5a2b23;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd79aa5ac2e3aba5ed881a69fb55b9bfe545f1f840fcc1a74d35b18ffaae58cb174a8b20b1b2d1c5453ddd5e35d2a7a3f221a8e1a7be1548f8ccca3831512060f24df0c9443193c84;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15170029629d321c6119be5ae2115ecc85cb7fcf141da9ac5c268e6db4b2abb8302fdf93c84c15918a9dc584817c6de3b2a2e695ef9439caa612903b99c4a3a640946393f4ab4a0b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1cfab5fe7ac23f399b73a060a1919a22412100f3e4260a67325724dab959405c88c353355c85c14c749b20fdbe01cff4f03630dd84c6e64d3a87ee7357812690af5c32dbd38dfdd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd43d7bf39fb337adf4a484da0ccaee09f45d96fe29fc76abd1b77c2771cb74763ab770ea0e145f9c5f9483c912ff96d5827a37081ef82a5a5a0a96965977d32b02409c3f2e54f129;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cb125742176b4ad20da6a6803c77fa268d82136d28341ee572bc9e0e6949f7002d2f4ff494ee9b41964c4f7963e37fab0b3c489a21025064fbf56d2e45d45cca20d64da94c3dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba2a15ec9bc9a8bc733e92a09deb69adc90e1d6a0a0f12b5d91b9ebe74ed1ee2646add741b3f3f7f03216ea7103c174f525be7c789423f1f7846af1889468e460c9a74c5e5045fb5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0d56c811626bdd9fc29687ba0985a6405ca970b1894eb647bff7ab173840fa81a7df6ccaed7a410be97a1bfcf51595606f93095c8af7d617014ba9ceaa25039dfd73ef2542460;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bff14c20ee58fa760e8200183d74c80e3ec80ffc1e920d5a3ef8cc0fd407051d3962cb77e16f1a241e0635883d5b57d2a4a569fd5dc3d0c1bc06ce0b54d4e1acb170282d00195b6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7b3d11b2451d1af58b29150e108e972748ac99b5e5b3ef53349084b9ef5f3a05ee2e7268699bc348670f01acb6ce6805583d2f99dcea35262f5221ea55b44343a93849d6bbb037f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78d5428c0f0d4cdb3c6da8990f77a7ce30a13de6a9cf011b3b9b0c97a6e0035518b3156bb0264b86a23c3bc9c9994b99fd7916f9c34d50f93130b364dfb9d83d99de37309b575412;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6411c06c493f7ab73cb6dd059417ec8abe2e0932b9d0139748f45e9578d6079abee1524e452aeb1cdbc97df0d93b3af9690066d840ec8afdb360bd4b795c8cb0ff90435b28382a4a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27cb46847666e044e87ec54addaf9f3a5f64641477327e853e159516e4d23c80b1a65281d230276c543737b6a8e3b201e878fe64c1bbecb61e2b01d3cd90fe1f1b8f89b118910c8a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f07d173808bfa41fdc2232dd185f70a9ccc227e76255e5772b7454d1d8f06b38608891afdc5cffc04d5e691b7e674340bc8762e6af5a0a2aa0f040bd675fdc6c3640e0a792d516c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9b17bcaee2fff2e7495d4ff1eddb573463d6181e0a50b2efeed419674a815af1b4450975c3f45dbe131e69167dd2be8477b480fd29cf4cd493952844120f4e972d92a1c87d5ea31;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf3e7e4d3af4dccebd68d552f71cab8de7d72fffd5b5abc2bef85874dfff386fb1474357b9c5b26a39614d8f4a0593e9eb40a5bd0ca60cf2929ece4ff4388fb05f173bfbfe2f60e1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f1ff2a4fb69ae909ed1c89e80b3ea52400c3cb45e1d2e747ef0cbc4ad5016a639dec720fde208a8c34a398f8114f6dad414b8a724001b3c6500742106646d1b60396131235ef2e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d0269e3e34a9a78e8ac3be2a9a0bed0ccd1f3c8b71929ee187bebcc5e6f5d9c9076af7a8a4001f5933fb717502ad7237795807cd90a9cd77cc65f279d9b2eb26a11edcd0a056ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb024494c362b987cd3dc75d69d0116d41a19c75c0221a24b249aba2f89659d2cf334ff59c86f7cecb063c09f84cfe01cb94e043b3a5cf4c72b05f0dc6b516d50b0510ff91dff9224;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef63d9bec0e4863b3b7f5c5b388d2674c13d7af865f35f051beeb673c74d0c81a85869888443f3d1713861272619320f8309945ba2fd47e49b96ebb2adaf997683113338324b2cf9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13175a40437fbfd3f2a075c84a8738b72d0a172ce71e796b3e73ab75fdc40d07b82df08ea63782e8d45329e96d2fe661e2e9cb49c87bda695a9f891a5dbccd6d6b820a83accbf3dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe2d121fe4d0193e64d5967bb4a6c3c9523c971849b701fc5a67426389717dc1c5920ca9b6e213dbf55846bae72ad20eb4ba9003807246a808c9e9ce0f809e84b39488d8c5da93ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha49de7939c48a25ef1775032d3bd7c0616a446efdde1ca1c4a3ac86c214874a87651863ae3ddb2535f959ece349de653cb279c2f3558ae41d00e373b9d55e5848399d2a8bd010e62;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h867033fc5cc571c186bc3ace3bae14c1da7893c527f6185e611c7dc21081c1390c7b36d04734b011c02da89ef0f88b2f5cfd68c799dc0a72e4dc71893fd9707d03599bbb1157a1be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd9cac0b6e6e65e681b3f693298dfb91e6cb1f154c24c6c9a81487e0dbc520d2a197bdee87e59e4656e320c5ce15d895262abf4e937bbd5b4683c4335dd1a49b44045132bdf32cbb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d1b61b9896a3c71585cdd7b0758b16aea1be441902b29e179bcb7fd6bfcffbdb31b608646a7625a7acfd887a3e501810cde73dcbf158229038ccfaad4be377d3355d3880f7caa02;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5eee63da811f029643ae3f8b824b9b18cc9c27fc5890be1d21b0c45ef00688932a6de8e9351ca427c331126f678c0dd5fa53d2249b0d3f573685f6887499c3cf4e5725059dc75920;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9a5f428b46c8cae99bb0135b910016aa77e2b6505df71dd7f17e041c9291bf360feaec0a7931d0c56c5609d89c99b466feadca702995311e0b78efa449c243fed184ba395c3939b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ab1e49efc2fd7353e27cccf38808dd2c6ef8072ba3e43eee81fc3d7c4a9ec33cbf68390aec955a57536d281570f4c6f44eef7c1196e3ed2d6432deef0c970ec73fd26ebefcdb5d9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3425a37dfb770905bc00dcc5fdf7ddc4253578e7fe7acccfb9b638360d434442790c427b12da505550759ef9106dbc95c3a82e3fd6df1c0b66f1bcc2294205931d75a2c438c1f6bb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68e71b8c414fc5e91434590cfe43942a0e8058a5134b7be1a225a7ddd1236e3fe0975dbc4113276cfcb57964acc124ee4ad925d9805694a823f7fe95dc40db5a60dae56fcfaed391;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hacb422c5bd887ac2b80898d50a8962c76f70b4c2d3f43af1a23443d6dd5015558b3167629c291a0ca71c701e8957ed075d3ec13dbdac337e2a0ae264f013e6f0957aa3e185b84d2b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb65b3a821b706f42f11ca0fb6a5c34154d53920b9dee68358668fcade5b250721dacc9770722fe529b52599ab642456345e8849798d107564b3b908482e88f0aae8edeafc20a964f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c349931c1a7406ce0700175d6d269fe028359e5ddff81ffd54e0b40bc70f350b904575ac57dede28d4b4f6aa42a40ab31fbe61258a3adc0f9369d0079000b709cb48e7b27e2ae4d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca08910627b053c87527c7571973101180b31d6bb2cfdbf1391d9abb20a3678d74b2d006d09266b3abbfd2d1aa5374c9010d93c8435bc3a41fe597a7602e576e2764b58c5180c2d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd59935c3299e14e5cc5649401a3dee32efdef4d45b5ad73c6291ad18ad65c63bf1d3a7ed5cd60ed7cd17717cbfb1e88e019bdaf312fe52e07aab2895ddfeb4b393751cc12c2307;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h773d106e30b3ef7dc178349973c28e2e4fa6abb8d3f36aa7e5eb8f1ddab8b678c27fa5720c0e4fce6f8bf175631bcbf7a3d39f393ee4d70138b46218d1a4384b878b817c8379f92a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8de1b021e93e421b0d26cff977ab7a41ab6fdccc155e02fbf3fffc498b1c4af39caba4e63179a0d205e72eaf9f48cc31f604ce1c4a866a984b99d95cd358fcf4628eac75b4eccac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f9dd5be2bc8316b08d0083ed6042134f228e3c924b0f64e366c768821a7bfd911353e8d0671c2d853bd3848419d50aab12cd08aa1861add5c4178583748a06133cadd3d97da964b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda7db104af61cfd509f922737ef7e898a49ebbb199e91747060613cf450d1e130b3b5e9a478041ee4ab8928c023b51cafb566e1e05f1fba31b8c57e9ab5c11a87f4db65c2ec8f3ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4700b6975547d7239650b5ac1e546a81a44bb73e3f82d7be11286b30cb2d8238faa04db28822f5e206700954e51b3816c8b620b2c82f736d00afa217b3b51277afa9cae8e2e2f72a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56e65a778a25e3f6cae55478e461127f5ec0bd8fe0ea51cb92137036bc472d37ef5369f6c0fad222f2fe54489d41a93d68bba462d25cdbfe311cbc073ce49a2cc75305d377abaf1e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6f0c4bd15644ee4a1a3a50d7c5c06667144f46f443e050dbc1a9a3c4dcf5067a9331631a2404022eac62017f4c5d8765cd987b03b4308ffd4b972b3c3f7cd92406d7454939f1408;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d7e333c735b6a7dcb840403a9bdbbb74c6264f3a170f8f850ab5632dec92bc026ce84980234f12172a459eecefc752f6fcd7b06942faadbb0af79fcdc111e25768d6fd3d6f8cd60;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb16d08229603907ae4d448bd91dcf776b77db5ecf9cde84e34bbce5e71ccf2bca438d32f7188f0219ac2898fc8b80d9347e6933f9ae33c73502db3a07b76825818cf05b670de576a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51952c4c7a9a2d74f7eadb7655fb67aa2aa9b00a1d85f6022a0304ae76ca0e7982b990e47de22b7ddcbe6c7b389941503f0af2e9c5bc9efe8881222440aeccef6acf3210f1c3b079;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h413f0b6dc20472d10faea85fd07b34e75a695caa010c56451e607df297611a49359d0ed4f22a73eebf2ef9d285d7709ec186204ba1b348e2fcecb0380882cbe804600ba85b62ed32;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb272fc347187999f0d7939694d4ec8c1f47013dd66c675cb9769d614cee67b81c637f26d2f3cc11dcde19c1c2fb4b7464a676c6a372e8186700128274e1fb0cbb7daa12ad94d5e96;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h953f61a32a50cabf78e3d389872cf8c3f63c90490ff5b1d1e6008bbac37dad36576d5941e96998952924908e01e193a7a1e1f5cd06c30b3ebba32a108de60825c6b627f7ddce28b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he193d30cc9eaf723cd6b3cbcaded7d61f6ab52ce3568165e404052b7c24837e4730fb29d9ede2cf1f71355fed93895068dce1ad30c8dc84537dfd500f224992ea98d1be8d0183cce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h795b6b3702c2d126bef58b0446d0c13a3241f9c4129f753ce6b0299a7553d791e4c4a88705f378ffd59d6995c5573d344ccb8398faae4dfdbd991ecf1b0272b7170564bd835c0f37;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95e6a8c0aa875360f5114dfd9556582ef77edd824585836514041364265ec8c4a88ca7e8f603a788a3a659fa3a053357def0e5181718c4852450abda88b0be85014e9dd7f93a4d07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd9918e3d29c88d4b08f564c18bfbdfc92b9f186b8d97ed66e53ff8df8ef7615208fcb31383f64fb64886ba37eefbd5186958dee7f00ea3ba30f14d7a9e61c48212e82203df6e8e3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52986d0f0fbc780338a8c17da7a698b588dfbd7ab5d6bb03bf6f6e9bb480cb3ecfaa7dcc6f24e573af6b97370cccd2aba9db44f61db6b5c456a4acde44a5d4fb74158e3cefd20f53;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haeb63af5ed6bffddf72713247904d09330d113bec76e9407fd1541e106985399530c2e4e2c04055a18b2a3ec61c4fc2892d0820ae88ccdf1bd0566f4c31697484ce615923e2729ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had4490746952814c7c0148933ece1758864a101e18dbd34a1f9966c0b197e8951abdad3a4557d849b45830b1e3c63e3c49c6adbb4c1199a413ab6715e4802140c922d8cb1886377f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha049f49e6d1e0f37220cb2fcdbbbfaeac44c004b4d9596be59699a12cd76a598528156cb1d0a937dd4812bd7a85bcc4cc6a35533391d15df526503522f74921750e1f342ef0b7982;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67aa2639819d6b1964589b8a7d0cab6f2810d1bc133a265b1951793b2539b1f3ab8a8893ff0075ce3a90fb775218642a5b503fce9607b928d8a7ba0b5e82fbbf9d58fd3cd3616105;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae3a69fb6be9775f2f33761f43b9309337fcc3c3b1f4e27e422f3e2af3266d79c56044473fbd2d5327071f8431b85d69fec756e5e77b01b9b9d63662ebe1485dcc1bdd09d99dd3ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee1fb818b33113c608010c8a54f5ffa13eda426f7be3f59a58f16e66858b814ddb1c84ded223ecf1c61aecd2458add1e784e0a1c66913b4927f7acbc3900fe0e014663092d3a27bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0f9dddd054ec9d9c21c8764ed3f0225f5727a85f78c84bcec22fb2e03032e53cf9124c387ab4b1ccb1da5c4c19613b1e09b6c0a3b627d6cb295e5efb8a9b65a074499908fcee77b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c7bed7ce28965e7661838e1c1efe9846dbffa419b2ef58ef796c97134d301aa2671f36ccc278a7845a81405a25d6879a4c17946426634e9669561e71823657480115b7825233797;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h814f7e7dd4b930074bef5b195e6110a8c860b98d0f0f9642822c38804d77fa560515052426e04ab1d14a42276c908131cc7da97c008b5efa2859ace0452853c6caada217844584b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ad993fb3b4698851c4ebdbec2eebe298007312562103381f5ce20a9cca422d62cdd1d641fa5f4a22fea768ff03073e15d882002ebcaea621c1da3c055a5b760a344a0ec73c7cc41;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c9f6699e13f0aecf2f73f53a133d25966ab0ec27276a220f24f91c89f2a76b4e35d78c454c23bd2a9824cdcf7dc900a05325640366c3c03732fd8166cdd98bda12b6a536902ce72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71b35d49beef3219f6ae0d4ec58533a966ac2d0fcdbad4732b9f2e4cf57d8c284cfa4c2e1f9059edaef0e5ef36f1c8001d884a6ae60ffa408f0bd93d8f5f2b20ee5e03fc9fb8e0f8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2760a4916ef7d26befa180cb7d2ca93e5546f928a1655dd1aa6f090fb9b25235be285114b45b4af5344c4d814506bb067f6e9433a0b430fd5695584217a93b3ee03f6325f52956c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fc885223e8b50da7fdb471fb03707975479031f95c5b398012ce30a4ca2b085f34f482923c682c96a175495bf0251810a6319be1888fd97f9062825411ce04a3a05810877d12fa9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25e0762313c28d0ec5d90fdfa67d05d8288934ef0f37522f4009c8705f9cdee30c3d34110e0031a9daedc5f6daa349a04cb535a127b0506e55d69787ac2e572b1464fc0a6a96934f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafd46ed3452325375bb77b043b84b6565835f4ba80c2096dfda2740d0c248fa4c8852170810c5a7f6df4915c204f9c3361236a915ab5cd3b5197b8679c5ba2490ec116892f172ff8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98c0635ddf43d2a6cdb14ce073423f87dae4900078503fb6e0d9ddf4448bef909ba74d9ba47f4ee2226bb02a0514b66f79e67acbd86652f8b43aeb3f81e1a2c9ece0c66dc8b6aa14;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef8b4564db72bc9782b206c1df08860d598b9ff0e11ef26dc8b6468c18c0d4a992552a362fe76561a61bcba9208cb69f256fc2f40dfb031ce7efa6df5a42d9400c73096344af242d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h436fc232756529c9d4f50278e0d4ba887f3d07085da735f59dcba090eb662c391fc82f609074ed20ad0ea36ef9557f6d7a6e979b6c67e4876dbf9f5e6045d00a27f2b78685eef0dc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h360773672006949d31dc8d5ab633e8236b12ba77751c5769a795c44704b7b3e17836ac04556dbc6a59c0c497e6ecb064d8ab4f5634ed41b75c742645840bffef54d1dd8afc85b0d9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb089cd7502e7d6cb82adeb11a7d11ef365bfb127a5cc1df29f4dd1f40febde8ffc4f84bb123e9ea02226920d2b46d502c386e7ec7b02e830819d9706133b284b44d046d330057d24;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8b2a680a626a8a88f7237c28d63ff06aacb6fd4ba608413485cbf3e363791aeb0927f6c26e04daf79f577c517465b2d10f3b628c577d762ff3c981966d1f2fd6d89c2915173937b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9a1dae433c4fd927d4e92afd2694c156e09ce9eda5991a972f098fb378d99e7df5b8ff92898d7582e480316150a40f34c001d9a249aa344ff35116d8a2232080fe2cd11d18068c1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ebc2e43a41080ae751127c306264ef0bdcf0c3235c3e768e6610625c58c855c04cba0fc7f0f33c2b80e609ed1554d64f565e0d66de01a0ce3872a0c3ba9d2e8521d8b9b80b720b6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9f03c6e6462b886541dfc67389850f73ef49b1aa52d2c43492f2a06c93075a4c36edda585fa1dc141b5509b14a426ae91e25f026a53e562f9fa2543c9bd8d3aa7820bfd20925b07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50a01b2f72551bc76d07fd2cbbb066c15edc05368229c0c5e7f0482e91af5ba489c1b5fc380f3c61d1bbb6a466150d25ab829dffec4bc053a68a9ccabd8dc9be10e01e63b7e58a75;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c7a7c626e10c1fc5b82845f5f48096243f73af34c273456a4e96afb123e681ba2903a8c7c274f77bf4c8a8079d7bff720adeedf00f6a6d501b0093dd9fe55329033004e563e545a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52bfed312055a821d69312b1dca0149ad42ae479540357642a177223ad6b42be3c621011fba43300bb59b47c94c7a73b995d9f6de878290de52edb126e48a6882ef8ebc712f8c8e7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb334b117b5262e3a5f75bf5b31f2b1f2c6d24a143f7b2ed0e8f4de1b985318079f82b924ac3601679de288c38a742aea7241e803fb5b2b7ff712378d996adc387a3b4e2953ee4b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a5dfe7bf9798fc10f7b6c43fba53e647a9d15e2e620f67705a31a9d696db4b2d3d439c8fb7519174a3a1e192e69ba481afc65e3d5aa033d88fe11f864b755a0fc3971fdab0191ac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9904e6d2768b51e0e91029fe55cd9311c8f3ae06d2bf629bccf1ddfb1f28d54b910cbd7f13ff8e64f4a84781c918e7fa7600bc78d9e75fe1245bbe09b8c18feeaa038d4c3203065;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4bd6fd119f75d8a665cadda7faa0102bd9a5461f346c2ffafad6edad625c54cf7796c9457a96155afe85e3328e4f44f3b316d856680137815a7c52b1087512f8bd3f8882f2ea85dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47c96acb672e4379bf06160e30c487895d10108b27a466d24968badc20efe9ca74013c0ef69b43a89d9991fe4752b80ee8c25dbacad75718bf4451940307db4d65d5a0ef5b9bb999;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf194413c93c070d67ce96c82ef08bd63bef25f6d846be1ab04095fe9002a6b4914c01dcb3d97d59da5cdc94a5790ca404cca205e7c5da9bac5c7e4440feba5ca4bd1d3262c4c00f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h466401c2ca54aefa813138689dd42726ecf7ba16adf96f8aef28b00c7247f9c4d4c8764a68b2d61e334be025d78b3e367093fcae49334894759b05c6e54034db7fcbb0a33061cb1d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h998d10d424fb16033005439cdbf34cb5eb9eb7d7d6bbf5f4c1c807d77681d4e336d182e62c6abb0c96bc0a9bd4ab4451ff48cf2d325d294332dd57bbf8d6467335cf3a2d04f6dd9e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bd0a9fe41931ebea972b1ed6b3bf621efe0039ba10b5da41f527d3fb274e9877418060553d1290387c6e4e04771c3a8385bb5979b84491d420b971589b596a62755cfac715cc3bf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h769ccd9e2fc446a1b5e9348affaad9136ed6668ac1eaa5f966a48d64ba310ee5fed1cd0e26802485e7e5ec4682d33abc30376e589184caaae8ff7f0bfa27d2a46b9b87c9cf431d5e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b114dd5e8d5c6ca79bf30c6f95f113c254c9f72d72433b52d27bd0a7d467a2e3c9520b6ba804325fca6f3c1d2d0e0ab54b453c62cbef26319a7c4de196c726a0fa32fe8f5c03b7b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd028c29df81786ea5f3ef82da0a01133ef07216a8dcab5aaabc503415376e57c8f26f460db9d495ca922dd79fc54b0cc7804478cc578a4bdd9e495c953cf55da95a35f90a2513c9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d2d4abfa0601a7058163425a803b92d7cc4dc8fb83f074a6cbf9fea51c5d5c58ab97f6a4880ae54beb1bb53970c19bd04eb71559b8663a1588f159ea7eec2b655127631772441e3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf5df27f3e069f80ad03753bbeb502861ecedaf9747ff778c81425d73a3e4f3ba2f9a506ee8898da972b89b18e678b1c8fa07a303c084cf31d902e8e0492642a44f5741dbea33a0a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb618f3c7283eb7124c421d4e5791773fcb7782afc8c79ffaa8b9b12cf057ece23a8cf64e4dbdc29e6a40981019cb39069be24006ffd430dc44cb66af87a1239c02f35ffc53c27eef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h946a931ff568e8cc1ce6ece97ff33c73d95d3f370f1ff5239cf24daa1be4cbfcc15369c16c510ac06cb656dd56a98503be95a4fb15f217563991e7b4ba1cad7b5cb4538ef91b7801;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf76ead2c1a017cdbb6f0bef93e2fa1f64ef1df10654441bd636d67d06ae14f80fad4e235a474f58821c49e72fa78c1545d254422fe0ceb1d68c6824f42024ab9c60faf02fe5ee5dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9545f9c91a6d74ac6416745c2b9467a20b30eba6591f3b7ff94b9ae7f069e8349b86e8d3f1ff06fd67903ab9a540deb8b83a487f477d067b2d4a8eccbbdfb7d898f7530f863a1b8c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he532c4ee0ec9cfb51d7d43199ef5900ce726686b521b79d7ad518101c9a10cc74fe4b94c9a368aeb8c11dd48d1c8740877f476c0879c9fc8200645cf1d3359cac2097e5f588fbe47;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbd41343b71d132aac7497eb3a36691f5342e240cc85b85f2490412012b9d1b485b9c5610370511d09c859cfaf13b5938ab31d30f593e9cabd8b535345b0067fd4c52eb637486b3b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26fd71e072bec0ad6dda5a76bcd61d940e8e24b9ea24323019e868f01f1191c708059d23efcf393b3d29be1475ca2973c1e871d4279ce9773eb5378282793c6ab39dfc5ef9f15400;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafb5fa7b38fca271c68ad8c84018808c9a55fc63c38074f0e1bca190aebda731a2bb2d66c9ac37ec7eef2af253ae98a1d81a32980c67894711f56f2f005a81a52db648cb2bb3261;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e8ffc61ef9eb9af35973608c3b412f3528224cd5e7dca6ec8de29fa5a4b71d74d91c60ccfd5b94f8bb804d76474408fc166a245d2435e4477753ef18dc5e85ca9f7e851ad9a8c72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6094cfed2b9bbfb6335bd779ac960e55fadd919bd2a25205608207fdc1d9bd7e606ec3b56596d2b9930c55067e59ab278d8eb4a3c11e61d2f1bcc6e56c10e413976197c8671e9765;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heda897c9f92d9f0165399ea47af67a805214afe5eaa5ef3e41e9330254103e8818245eac0966a88ae2c1508126cbafffcc2c0d505055bd60889d88328c0d79149b638873750eba01;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h793a7a355494ee6d953a255b25edf394fbdb97db2e66217b83c084f57b0bb7115abae466a7620c1d555a935d37c64617deb3d1c1ce659d9de9fe7b11ffbf8ff733a2579976823b81;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb018f3cb2d7acf45fea08af8f52c0674850dd0a7a92dce5bb9f6ea9c43f17eaed06c5f01771d2d4d620b411a165fae74c80bb4725c9e1348525ea9fc472be410887968c419acb6e7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa92dda1696a82d224a63ad2c726f6297aad684658f9041b9eedd2eb548af4aa6344abfce02dfa1f067f6063d721dc9ef7a4f6cd1de69d050c75b8753e04200987ee8600e751f67c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd039c3982e0df5816184793b1d0bfae117d6253ce4868b83528869ccf03f1003af1c36f36e3e455eced1a5e994212e82395ed809ecdd5c0e400ee597bfc32ece3d0fb4fc1ea9cf95;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5e8b1bc44829712a5fecf9fa6cb42fb78d8256ba9bcaac11643c2a8ad55ad809cd81d4a1d8dd9e386c7d32a3fa0472bc60927b0c3eeba18a565e16c31f764d2d41161ec69040e77;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25f9df993d999c3d685bf1d3cbdb63b85133607254908d333c8f80ffdc93d6c94f6f4f076f5aaddfb3b0b230d2e5414dedfa32f2d684559630df310e6b30e65b5c564390e4b268db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b6af924b1756939d9a35f4cb530098edec2ab910a46d00af76f4fa2d1fe706eee2d80b2f25870e941487b37746da1fd3fbfa47c8a6d699aa13d82ca528811a7baf21df8a87d708a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a7fd6fd02c2f0a21786fb725e4d7bbf8a40d6703ff915c00dc46eb5aa670e0954dfb5147a7edc3d549ecd7dbbbefe17a901c487fe4b66f47142a9e021c288bcb7de3206d96af807;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e8015866bc5ffb513619e6a4ed498cc99ba2d4a601fea1a01c1a469ea87688b34b1143b7fb160bf0360079b0f64e85defbd984e0730c183ec8560ee827e2865d20fc3f5b64ee4f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3fd0cf0e783272d6fc651115db5c92c88966d2504b67542fd372e743bd4b8617b6816402910b7b867adf9b0bb0db080fd4e8859bdaab00eb767960e85eab8d2457f169b0187920cb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf408f1c78ccbb4a48f575626c562c95abf0a1ddf5515fe077654acf329f49beb003a315ece828724bbc2ee0c9966166a3e90397fb0d59e09ccc6849d484623f2636350bdb3e8bffe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89906f00932b13f3890155bccb17065cee40750f154ead956a64c0abd39400300f501211595f6b7f2afd916ff0e9138777bcb91eecace2573ff46b650854401f40ed9502726aa490;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9561a4a405e008573357f102e44b4f8cf9bfa859d47445e14da6e2d1220cd32d051aac963ed68099c623a0fd05d5424d30bdc00f9dd63e8688beb9b05df8f6f4c3212f41ade03994;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h323a1bc61036c0d461a8a31174d454e14f50e0e8634f7214fb4bca25c849ed993bc18c89783726fdf19408fbbb2dd4e643c2135e563c459ad6d7897f92afd1a4275bc08ff637361c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc92d6505978d6b758a08bda224ee581ec7678511b88ed64b8db4f682b0d9c77dba2f90654e382a23b739346be28e83a2e1365202c429ae3b25f48740aa4d0bb35c5e715eac6ac9ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7345fdd94322de5e37c7f6898b423f0067c9e0492c720af2d9df3b763417fbca6c9d1705d30f10b3b35f5e740a069e57b5f048518aa47ec5d2ad9a43b7bb882379671cb2d5e1457;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f2e424f07ec46bec429bf223b8c4af29cb42a80db5d65b5cd1c64f3d7bc8dda7fc78106efde41225a18ec48fb7338c9da15ebb22c2d82f99361525b44aa47ebdbf466f2821c9b15;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85fd2059fd9219a76776cb2d2d6660e3a773ffe8df1aee69d3030f4cc2ded1a216e063b13b021f8e6ed4ee4c251b9b50dfb674ebfa713dfc7cf62e0aa08b52553eb069bfee1479bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab89079705b39d92d5e4b953ddda8451a0cd555b668d1eb30eec4e92877faeb0f184601ed4346071c8993bbfca741fe115b97569bed0d251df5c8f071353ded52a7ce4387e43d866;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ab0c3a504dd9e384635c20468145d6d0a4b473fdc30914363d90d0b85c288550cc2fe5df4360cf330b4b7544717b7cb6da79da8c1ff6953b6629aa99e971a427f1ce2079d0efdbb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2d261dd553bdef38d2db5a93d668711f2edc89c18b6bc514bda5a9c9732cfc5f606b6f4615fc47aee34ac5295776e6bdd76da1d570a967aee85036f08f727dced02f04ea62d4c2a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c1c7fa984aecb7158ce3ffe976d5ff28ebf9803cde5fc6698562ec14bffcf0c9d6ccbad97d4ef4a9c8f244c94622c5f07309d40e22ecf0e7cfce5f53a1f213b2aa490e93cebd68;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce7e06c901fa9a2e8c4a5657ae0df0c7b6f5c97e1ccfd8bf8a80b4af5750f36625b7c1cc8b4c52b441df97203ce99f384c4b28db5269fc961638412fc7067571af86b7ad4e55c92e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89acc37dc7dcf2488ab6acd0fe3a5ab25155229415293ab2804796909149a695f0bd80cedce78acee81e975962460df79f36ceb8ea1b7915938001fd91d8e94d7e21caa5a518db6f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e6ceda362ce51af19cc567b5b637586328b32002d4641b45e580db31889487d883a6e6fc215a7848f6e3a3e194e073b9f2cbe3e8681ed8e2bfca85a595c34e0ae4d20c2e710c1fe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1dcb8916f045f061d27715a1b8a1a82cefca0cb59d8cf3bafc2b70a326d045f70cc5ba602eb6f35f1df9ef76f955bb07d93968097a988342e18b94dc7b0791aa7e68e0b42dea1340;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd04aaaf32d746aad022d518bcfe28cd45b5bbd127689875af9da91293e9274386052e718c2c671140a62bdf04c364f33cb709b14fe5cad09afee937227f6b6a5e22336c4d0dbddcd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a67acc1d1fdbcf7e8d03d908d334cfdaff61307340c458d7de474e1608286a6ae8b842a2b66e21b15faa08d1b18b026dd92cb70318135ed18a120806d496da19b446c3128c1d962;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57fbf893ebec342406533d4c97069346348fa69f2ea910089771facd38cefceb34c676c814c62dc2eb13fe3e1bd97db248005e0bd169133d122b9f5c7ba2f9f755efaab714d4fc4e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffd39bc301a73865a3dedcf3b10c3a68bb290c40939d1e088ca8034a23a7edbb46eec86ff852d2f0f0ba411f1fbe01208f6fc5c0b969a93f64c1e33fdf7481ebfbb3e0ac8faea9bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f78672570a08d0ae7d31217d1695ef4e96ba8b6f2fa12a3f1f4d36ce8f6a9283db3e8ad00e51f9db3cf0fb6816fb44195112411f7c302a99af9d6b76f02bfa442c823945100d45f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e99edac8feb795fc29dbb11d4301f6654d9e746b9252d53c3296663d9a6985ac6f239d26835c02eb4b63afa31e0b420d13af971bd0e8f8f2c8dca28328732588e670f8203339da3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5a6142a6583f2e075a92b36cb4402e71c227e3f66005351acd9a5cb8369cabe9001a5f31ab1981c3dc90ba0d5dcc033853cdfe492234f18a32ce3b601fdf6930a7aacf4dfa5d39d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbef4a54275cd4d91e053c2e5e7b5937551432df7b3acd5cd2e288b2f0f877fbff97cdf1c5c3bcc7a7bf2ccca6d83d5527d1291c16a289b68d31beabf84ca3ff1bc9b13258e6b95af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a647374ddc7af24074373c70150fa71c3c191e69843a5c7f042a40eb33ea80dfa1ebce5ec1e8e318b546ee38834155aa39bc0d8afa0cf21c42250ca67675c2fef20c9d5516a1f44;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8893b12d4a49b58b531d09af1dede3434167112e3e7b727a45505189d0f33367057d441a1da942c5ad33edd2a22cd0cac5d4a7c44b8c2e1ca134be88f80394e18cca41b3ba17cdab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88b8d2e986061427220d59da7b12e40fe36379fa1c5c3d977675624088567775733b8135e38eb27ed5f05d09d4d856980d5af48f5eee2961a60c2d99243ac7b46f71010df7d48a1c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfaf84c3d4c77f0902ce5549aa733fba6899a8b07c2103b601e26b5cfceb366a3c5ef9febfbe0ad53d8293a22f1657b85da9cf96e5b1043e9fac664e2783860864d44122b5dfdab17;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h855096460041532683a5af26fff5c87b601582a6ea41f098e09e0581c796cfa6ebddfd007135e0317b9d4555aeac954bc442dfcd9c4fb3891ea6e36e937b52629761421b63a20026;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61189b5b85a20dd055830db3b7c1e4941a269aa4d07ba07c9ff6920acde7b4611c50413c8a9d0524e457d690e594a9980f4ab94d199b177e451cb2fd9d114d37cfb1889b61cb5d68;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1c24c3a27a23bf3dd138109dd0b7f84d61e119037d556dbb362a7d8e83b6012b00ac2a37ecce3fd482e9de02be1856640ff5ac9b6068546af6e3b16bd7b0dfc52b8cfbb2d7fceb0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h158a248035090303852f1273271a8ff55c9d1239827c1653a8d087c5995b5d71530e4f28f2034b7d03485f806c7df5e622a89b110f3046a66957172249a770e319d0cc5c1141b0a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6351b5f3c5665edc333c5a665fa1d4a694cc66a56a358465a322b67327f86b9ac9e00db70e9c860d91830429b715f2caa9dfbdfff5701960c59f996dcf353c9a0f6e25253a515dd7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70be7171c280bcc7d000831f8904128ef9cd59eee31e5bc2b5eb8ff8671557f07f8e95f24de8773951f6b81bfbc2e2f45fc9421a977b63babaabd4c91123b8d3c418f5a8089277f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he68ccf9d33a61380f57dd93965e53d16301f7f49d4f5de09526462d2c9e433632c5c2695558373c2455278bb2612c9930080637f631a32bd74d2135c5254c8ee338ebba3ae752af3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9f4d17d38256ce36dd0dd4a836104ecab07a3fe804ee119f67a1e19571237d3f67bf421def402aee3be349d20035085f08c032c1c75415e7a24a74837851c0b3325812a32a54f59;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h196ed10e993e706ce88278d06ed3d48c6cca094b6a8f2c1b4edd37bca720f84b8de3c1ba502c1ffbeac5987ec6c5f336c234deafca7a70d1b0dc8f44c399cc894d31372b0a5d33f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb00dbfc5b48d79dbc9daaeadabf4c49f9b7a6ef8c7ee1d1e9b4bdb330d77efeca92c00c48da7c4d4e195f6bb3cef31106329f2f78ccad078a418bbef8320232416cc05a0f798680f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h241b1853c4c623469054836b1021c9048dec60a2f8dc615a5f9960192578fe0e28f64b65f42f51eb3d45207c798ad02556fd8c19db62429ca2e72959ef028e8a67f9e9532546dc35;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h384ba287076a67f2dd5883419e50154a9a0f7e3af71f03343855cce2c8273adb4e7cccf36472c21899fef30bf41bc61909bc89089f21f3d073b64928bb18db6768f499867d1b4453;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb9ea8bade3cca8dc7fe1416d26a970849351bff2f02fd798bb5852e7b4d70605964bf27144f850832783832c7f979da286fa169c9bf29c3b3e32a4009d38fc20e08f9f926d048b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86288a9bf68aebe6c6890e415f19fd89d7921c8ea503c4815073658dfd72b1a1cbe4a1bcb910f27b378b3c126ad6cb99f871daefc39b917f56f5d02e63af51a675c7cc517acc3d6f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4562c826b36df8fb46da73ca9c15b71f090fc885a7e989b2b71e84f654b9237c616726db20833f03a02de3ef9c34e4981210386ca1b29521d6a9bb6e0bfaefc6079a40c3cd4d9e3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d598cba59b2c6341bb8c02391c5be11bab36cf3137e8ed453bed81f6490911c37fc1b577d67dfb33c443efe2aaf55e4f74d2ccdc676f2c5c92e68f8b2c0375274a08c29f9215edf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h835f0de9985dc80b66bcdb61b83cbff90cb521b44bd444c6755b69e77faea35b4a26d15ac9727d99dbac763fef60b5cc8e9a974930dd02d3d99b368d0ec1a7536cd2dd2d07cae2a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7624358ec98de7df65c8eeeecbbb9e90873e7a2e13c109ae2a0f3b2e7319e92340fe3c7bd1eec2f684b28accd738dc955b2af7a57ce6b40379de2c171bd133fe255ef9293dbea84;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12f09b1d068d3e8186ddd4dc28ca7fb5301db75b6ee17bae7aff87c318bd6e8d15d466e1754e133ff14be0e4bc8b90b77424e05aeffcf968e7174f4a382824c05c1b0225f3f908e6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bf1d3af1f6fe7b2fc6be1ef23122ff8b022b0d867db4768605bcb2d30d0d65295a443b349a939b59662f242dfaa975e2815782126c7a3dad3c1f85e298e5f726a3dc2e4469ce97a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb360f2249e0874afe7c6e8c937905801f452517f4f2c5040b3f2cf08e6f16a92c7c28a8ce9288238da41ed49d6247043c7846708309c38062fd0f394ac281a7647f3e83b9d4e35b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6de1002bf286d9f63a587a446fbfdc7e102edb21790c3a5067232040a02ca0285de0fc5554d49709425549629b9ccf454efe3f2789f0b72a6a114a3378a09aaacf8b7c7ecbc42b40;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8e104809207f29bc971ba09f072bee2cc402cf33959af20da9e0c4960caf418d1174139c88fb1ec3cae452d86d3cb501773ead88571a36b249bdb5fe51af434d1ccf16e2101459c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28e226cc3c400af131fe172d3d66be27c05d0c88f26a3a0f4919b9bf9770bb4be9c163e5ce5d44c32b2a7982d4c5acd6945bdf8c6777ae76fc9827706b344fbc0124417315441d44;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf93e542745d4ba1638d8f77b831e7bfbcf5f0ddc5fe18235058830984c3bd74156075cc14e3103e3d995ccee6bf7ea7ef62e2208dccadc3ad2815590c67184478ad714b72526856f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a4e145ec0828bde4300c919e731170459f1307648e43a40cd2a2d68cf6a4121c32963dfb37ad8bc126ebf0235fb495b1ff38395c651989b0be8c39946ad4ec14a6a32cca7c5ed51;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb194dfbd2b2d2690ed6eec440f1db4d862e8d6d6b2c66d2caf54076ab7dbf07b47525f9ca1b7e99b8b89c1baa7a6740ffe5a9fa7d7ebbf65b63bf35a3d8f5379208b74b4b5d2999;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1bf5796d7a4119d4598727eed25b05b9e6a265662d2f00f17dc7e082da57c02dd92fcaf03868940a4687229a96285157f7385ce3920aa35af64d4c0b7853989310e3b5cd42518b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd082258f8fd6af350e5ccdea0df802ba5d6759556ad59786627ca0921f7c7440888a04f2a7689a407edb36e17b7d2638be013a4452842c9c5d2dfc31fba14a8ee69e7dac10ba826;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9749a45fd6367b414e1d9b24ac3296f24cd712e402612f67c0f6f346b00115fb672b5fc49129d60d5a0a5e5cc45dfb6e5043f5ac60c93b5d63770203a826ba84273bd5e60606653;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58477261d0c8739654e870ca9bb89c3b7ecd8eab6436bc2d793b07f9328edabf4df6dad8d04ce2d1a525aee18e37cbe0bcbefa9a20877dd62f3a8f502024e1715176bc41fb0d2dbe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3729e8e4481d7a10442e41094bb41e4b8bbce9e2d24a225b4f2c8a2018c35a297867bbde2e22e12a9cd7130e073721a8a37c445b2d5e2114f7f573269958c8dd5c380f9bed74228;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98cff8409d9600bd1a934d1c9a7567655ad2a393e9f5f7537a2f001867ccab8c6ba76b3fb96c6fe9eb81aaa9e17e54ab6f0938cc9f775811b4ed023d894cbd172f6e848967f8c70e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e6538b82f9858efb6665b1442884701064a260dd6aed60fc3b9b0414bf02bd3e012c0d1c72c9ccc6c11e07afa5515f727dde833cf0db1d826e374310db1bfa4a1b15258e288aa99;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4848e1737ba215cf385a67a68cd895b27072b14d89d0d2d67371f2db1737eba6a70a8816303f6784c85f4b342b5904ffb76e1cabace17c2f2c475c28dc93e2f5ee52efd9dd5fdc4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68c845632c0b8de1fdad800e0f66328f37ae1b5a3c6ea52312814c1a4b5a0ea5d64b326c324c088c95bda4cdaaaea52bad498015fc7aa0a0f20f476bc4beff98a394a7a9556076e2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80468861fcf3af87f37981dc1f5e5eeef52c8280504d2ecd0bcc96f4ece6f5dc08852bd1e8a898bf1171191b617ec29d24a98c5411a51c84fb7a28b676c4a784a738ba0e0e8acaac;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2481505727f26472289cc4ef11ea518ee5b93e3fc4c0f482a990a9ace0eacf96fc18f77456a3f3d8dba11ad83814097286970069d3f46044853e250f327c79d57fbb7c101c406e88;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha12f33db69e5ecb76caadab582ddec9648d6c8dbad2fb79285771f4ce7062cd55426db64505ce7b7f5bc5067baac3ca55d9f32b2840058e37396df1241c37c55178603a3762f8615;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95b18704ce8a7eb4a2030449ecb8b3c69b0c1e93c3211ed4a24f74524c6d2c58cffc0ef03968ced2842276c106351562cdc4e900a6ff4fbc6af8e9ef2839c4b3b791da985be4c334;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5f1dc075c29765affe342adf07b3a43a0505f058cf6c0ccac789101613cd8890fd947cdad42de3b14fd4bec9ae9690b21fa6c4e4548a325a096db25dbfaa550abe5c16323f5075c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6b1af6dbc4e4dd3288273b12527405a40ec40a790ffa9327e7c5a9aaba55dfc305ff3c14556863af09101872937b9b39709e0ec4b6f734abb128f2a2a6ad3c076c0348a2dc4d3a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3cb476c43689efb5c97b2b19356768786b25a23aecc1817515d9a76208f9031666c277d590e0c028597fd211e1e119b63044df012c5592d333f34abed1ec02cdcd5bff3b859d9859;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45512e299c5d3a8f8959b7bf9fd93fa31b7a16d63d54d405572fdc1e556d1e3664232f5ac4dad4c6d8dce1f075cc001aaaf6d1357d4de6f760c4761a1f1a5014133ddc5f866fcdfc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64dbb170100231bfaa90e57812cf4e0206576bc0500f2a79db88bc4b2a8d93acdc47300dd729e566605209f9e7480c7d542350f87453a681e6b79e24e883f19f03df4d83a6b6a2f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9ca626ae0ccbe3740fa89102d1eb333d99d86e52deaf030342f007a8b30d6287949ed9da8a771e08d2ca3889dd4970c01cabf4fb8d0215e81908045772e8a47b97da2d2798a7385;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfde961d561cdac386e7518925b57f60190c011ced5f7178ad147dacf9b6b2ccfaa03b59005c68e3afc0cd46c5f1056e2ce6e9c33da6ffa3b88926e547cb601d851223bf9298b65f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5132d34886ee1de33826239f42fb164facfbdab39a1593fce986320017fba9b70b4f8fc70cc295bd85ff7dc26e3d78dfa757a6eea05b3080b131e15ac9ab575827c9f2651040c9da;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b79c90ba962e826fc7ff70e785c0e40b158a8d1faf634203e825da3f40b882dd939c86df3a3956b9a7b3443c0787114b4d6fb52943c6efb98757d716a1b1bb0afa58cc6f9a1de74;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb896716a792df96e5d528c002f951966b27eba2ae00fd2c0993045d40e4bb880f63ef548708aad136ff5e6bdcf1d0453a2582ee63dc0bb43f9b73ece105a3bb63cd9d16d9d625f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74bc17753fc15049280c24484f4ca342fd11226f55869cd653c150f26e1b35f94671b93b02c2e444c9520e55d6b731053dd0d7cbcc6c2e901e66cd65faeddde2c2d507db9b9a234f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbcc2c78e1514fd544cb14988dad2dd443fa3a618e5496964cc437275bf33456894f0c8bfe854f020940b10a195daae0f30c35c446012558de8dea1b12652164cdb8c19970c910d3e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb28fa7df3f3c1d93c1ea538b3acda8e9032dd3637a5e42a265cb3fa2ac06d1604a4c0c5a95df1024f6f6d2c2569f9364e96bb3956b75de996c91fde288c80d8bef17a2a930937c83;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26a380c8a270a2fc74eeb2f68d2fcf283691159a7cd79ad2f99e993b9ed7b5ff4250a8f5986aaab62f9ce1a68c3b3a50d40f2b2b2a8ceeb3eb81724c00ac2a71d0e69e18093184a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f1f675b472c7064ee474697d65b32c72038aca9652a020da542926d70e730094b8a7c056f2046943e90c697b669bb9219966900b452c234aba9f26e0ff304a24693219e7e9a91e2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d8cc1a1a2100b0061f6523a9bbd5abeca322c0e7e8076b9fbb01f6df20254c83a7ca58e34a0639b9c9881c2187f538b1b3a0f0382f702faabbf526b6270d2c10d97231103c59521;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5442b9c8775a3d20e857d8be554a2be6fb4a83837b1388b67cef3282827844cb15b5501ccfb25d6589fc559d353c779e045f59090444a50d0cfe3dfed006a09db43002b0bd730b05;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66f4128b0109329cfa2dae458e21976d7922377358f8bb97baf0e0c8fe40ced948552aecf18e89f12851983a09510105b0c29893380b6a4e02da9c26e756087bbba4b1c3428ffeeb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67af65162f90ca405a394d967bfaafcc7e8f4a8fe37cb9cdcad81fa6ad7875b47918004fd937dcc553bdae07f6062bc058c28372ddc4987f1f6173d272b7b6f025839e5ff237841b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d7cde5d2eeed85f8fa40a9ba9be7d335a9ab4982bc7691d30598459665feac707074c5d0b40ec1846a2c59f9ab7307fcf73c904ffab5f94948a43c56b5269e3e896fd7629ece55;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa4f8ea19dc93f61c27bb49d1902c61b1988af13375211173f144b90fc8352e6ca003c51ec4a5fa5e78a5309a50122d2d9a220d6148b40565aa3ee8d3a2f4847796984a170a36cb3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7490d24ea63ab0cbc3d68694332e606ecddcf9a473b6c5d539f25ff45f88d1d820b239ae86db6d86f83d051930b54cca2500f60befe689f3ae2e821e57b2d98173240cde33f2ffbe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce00a84b984285e8fd8c84054cc13db27805b4835ef8cbf695fbd855f69e1e961acb3eab7eeae3a0ad8c9c9ef4759792ff7d2e0a9d32fe8536462f0ce95e9b1c1d8f61aae2a4a914;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6799ff665c07d58a2ecef6b0c816a85b525df8a8387348376f283b38b2bf1aefb45d05827e32fb0db1d196f0701e2b1d48009c691bb0eafbe766fbc1d2aa405d5304bb3c733e4c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb86e9bf20813698793f5afcd4a703dc8a3194a0efbba0c7b8c2cb2ca92233c4552941f7311868d7722f598205bc9b58213a310a6fe388b8579166da1d03dcff9a1d67ddbe935d413;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd239816a3169eec5c02aba2cafb767e2f1d83694bcdc181b8ebfdd0f9dee3ebb288029989ece9c035a5608fa6982aa4944458346db6f5177dbd03f9ca2698bcf3099a3788810a1ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6b8f529933aa0e5ed8f3d639ca065fc0aa7c5360ecc05621d04dc73f5bfcc5c98771fe3774e05a6e4af2c9642e0f8f084cddc6513c4ff9937ff845e3201bbf97b76b7f2ac45e57a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdde58f5d4a6f1e1d3c82f4cff723547fc5a98070f2b82ce209c4f4b93dd83ecd56fb523eb4b0763bdd476171e9c6a09296e63ff569ff60199a90c5a151a2344ca41df883f7df6a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1b946799a2f24fa84966ab3c099f167c7c4c1207a3da324ec3669af9fb1bc16731ff802c74aabb6638b6f76a4f96c32fde96f0fb00a47bdeff642ea3b8978f7dadf7899d3cc85db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6647615045c6559d63ca8226839970d9d49dc2688752b199dfd40de8f3db35a982cd5603d7f16c5b3b9f0fe24f93997aa1a0786749b6dd2f10567a36905b568b6d1b3c72e05c5ba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba224d1adc1fc59a9c59057fa8f961c73b74169e7b4e6a8859fea79b2f78fa94d28f3330b077e1ec859eee5b21308fe4f5c31980d0c900013c335af61d0b391ef2461a900b6fa083;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7d59c480f133b85923a36c7c1842c519b9d2c2863c1a6c9d51c1f38ca152a8565f090125c093068a7014b8f38a7137061e4700d394118066c1af5b04d4b6f1b9c3717acf4ea3733;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4323883c01f2dfff0f74203caac1b188d7bcde0ddc318e73177b26975a45079c010e78dc69c2278094aa1135d25404dfbd260011e4727c69a661282a924ae0aac3d37548f66e2aeb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he44498d5d4d74e21db6deafe820a95b0322418c09c398e3b0020fb24a03fcb2c3893cf3606bd6c3aae64f1f91e7bdb8124c5fe35f4d68ac9bb47c1053329aa81a2de4ceafda4f2d0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9bd3ba0d0a6300340d9aee712b0a73cee59a351eaecf0b479a42cba9305921785c20917e5bdef0a871e8aa91976db689b7a629f5d21e0843b0eb197a8c14b4474c36c6cacffb0ba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53d891870bd81410db400b925ed172d28eaf9ecafcf0965b32767ce2f4101bc0b0835129b6768c470bfb5a54ba1cd5f5c624e0697eb66cc98c3c614902f47545e5922248dfc6ecaf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heaab3171c261cadd2f2b20d37dc1c49f65f4b562e067e4733b3d96362d68ffccddef6be2b1d7a34147076aff206e269f2a433b6e73d57619ee4d754b8c2c000ba819f918fa2533a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfed50eebe60d5469c93f305b4b67e67ce67b3005a305684f768e348d766fdb17f8d8f31f1e8f6ac5b4e49871cf0268085d928d9673c1e1ce2252635f0036ae75ebc9859cc83fb3d4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72936bd6f839eb2f025be1cac0c2ad1da214fa5e2be92841adce39566e4ea1483de03c6c6f9b407065521b3fafa2110845fee056344f93e425bc1c416a15d88df9dbc2584560c909;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h504437dd58ce21ce3119bb9f9047d124bbd42810bc552de8c9b7180a4c9ca27bd79eb52c445eae7f7015498f325f152d6b47d5959b8b1331b8449aeb697e3c3d66e5c76a0d423dc8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd293b9bfa5a0f61fe7ff77933fea0e6cb3a9936952f333502c372f71b9da7376e5ec8ae0e1df88f31f82c31eb7104d76cf33d1723d2a603fd3c4ee886120c92a94c0165f1105cea5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b4e1748055311b7d498c43f2843c706aa1d757f675cb1214792747f122fd4821a531f9ae7663eac477fc604b72b4db100b8da9431966f4545ec1bfeef6b93c99abaa3c61216e4d0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef3f516c76bb63ccd98c44e2e83ba5f44cf8d5a2a7714e787da07fe574b76b54c3db6ca2c6a415ad5bdca28485a43286fab3b472fb761859c64acfba655438993f7e52b1596c8488;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca3d9f4c7d081d6ddbae72bd126f5ebf35ee12c3e849e845cc24eef47cd0ed24aeab53049ea0f75780fac94f985552ce2f2e5aac1a6d39b7833865fc122bc312d7b8b9147164e07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heedfeb05433ea0b439417048942e9ec29031d8c84fae0322ad0ba7a66934860f3d63ff99f9f239088b144e1895ac90c7bb5070e224c456eebe6f4ce2938cd8396374cd16fe923e39;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf373fc3599c63920a4c1689fcc794ce95263ea85bb392e91027be869433c34cde3d8c61dcbc58410c110708dd3b80e195d7f4f259419efdf0ec654cb12e302bdb6c28f2f0da26cf0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e29ef220a5450d1044ff3f301e1937b3f08b1da0a043c97b2735923d0494286dd2aae1e26f0ec328418e4dd48bcea446b19ad20ef4597cc247e5aab3507edefe69077a3a3885372;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a01d4ba72fdfcc0387a72a3853e29abdc4d6e315b3044abec1624672f37ad61d62fe209e6effab9732e3cbd5ba80d8dd2fed5feb398a344a51ca92f19c7b82df9a64ffaaf71d363;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85903941e2df771ca5482878099bd07f3de64e2971461986cb02b088ed48f67cd55f1eee1548c614196141ee0c338f81ed22c8057fc52d3c29cf77dd423601c180a79965d7d81ea2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36f2467529ce928473d10f30d6e8c54b055f8d1ded3a7a6da03571b78f2ebec458824f9eaaea48095c1b34f8a00e429fe22b5db76ebc8bc2865d47cef956823b85857da5d56ebb80;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22f7d61f0870a16981edccd5e1e355b04f83a1cf18e956a43e75988256c7dde5814c2b1f61fdb7caa1fd9b8cace8d76e16a5140a6d6f5173d9e7c64c7d2a5b7f629b3f2fd800b74;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf22fe58db8b8bd1ba0e2c6ace43660679ca395b98fb1a3583fe1d208b2ddbc8d4720d7e34e3eb25df4882b8c861a7ca0cad3f03f8f5bad7dd151a833a96e55e0cbff5ea6eb573ee7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h333364a4140a69e479491ade98b0b2f6c469587afc0e8d6194ff441080ae1b0cffba426584adaa953bafaef94bf31e1284ca8f9c6d98b2c94a0369f0f8afc8de66896478e4e3296c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d50dccf0840ce6400cc7c42edade1b929a06e24930efd9aefc5991494a8f808dbcb3c462272ecb40935248b766e85a16ce51d92230a1261130dc40af2d24f5505f02f65362aeb07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he48eb6d588170fa8e7fc54a1d4db19b130861ca38a21b5df3e2ad9e72ea3329178e47898795b9d5a8ef468e15e90f5947d71dfa617f5dec6e15d6818ec37e681e8d8f5932a31c800;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66b1d6e5b665692177173fea5f35744e0b0eb2b7d02771029bdd7b0684602f817668e2a8bd442798f16128c6c78f4e58dc45328c97f18a11be85434688fc1c101cad61de311d60ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h641053db08032537685295dc343a8d669f22f25d700691e27f45518dc359bbfd0f75ff5d44428a1c94328f659f34ead38784f13f63b4c969394e6e26251ba14371c812c533ec253e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he045f7fca2d24fead0be923b02b1aa0fefbffab7486e3f191accab0bc9962368fd420825d3e0d196142f30159b85bfe22612efaa82e90d9e0e7a495f06eef57d012a5926a05e4098;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1464ef9c64b9fa361dd03a28924991671eadc54ec7dcc762046412088375cf6cefd70798c465988c60be65d17a00e4b39f09e5dc0fd8c4ea8a7cee62797cc36ed74053b2cac1ee2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5fc3ad9099876a0126d320dfc8089b6c811c537b606eaeac310b7858c094ce3ed840a743a743afe43b6f516beffa951309ee0682a7ba5fdab971e2f0d65dc08ddac56886c63a434;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34343c960a989f47f93d78c9c82086fa7a5be7464976048f9292c2ff3377dae422ff0133dfc6360c248cc802a9ff2c178eccab6ae9df9aec5430e3413899cec574c5934887f4bcaf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbda5f9619c69eeb661092f6b2780fc67c24518eabbce6a1ea567de9568816a81e8b7ae29fcac0ff024e6fc424d6940bf4f5b02c8946650ff469dc2fb20e03204f12ea94130d02665;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h810bc5ce35c3728087feaad0601a9659bbc435e537006183d787a4bffe3110a9e49cdbf010a3421c4ff998b0750bafd8115a717cf24ba3b35ec8d4ac6773a8e2e059253115f375d9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b2703e372ca19dfb38734b3e5bfae5d9196f96159d0d79484efc91c4e2870863f1127a5083e9d4d54812b1d87b1e67c16a011f794f5ea07ec76c775490e4ca7da43a0357de07d8d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4f80e1dc1eb9cb5eb99798a94764e21ac84863411c87f466f88aa5f2c06a7665c509338e123a46ed2a0461ffee48751bc8a858919f9c0d94a0cf323bf629a5f86723924c94d1881;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3d44026bd1a2ab201326937294bdb7a4aefb0bd7e0d00221e26e628d9eb6cb96ab481e13a57248416224fcad29c4cd25fd1c724363abef563e8713a27ce88457fd8565798ba548;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3a14336034d70b83ca1f8d1b6915d80596e4a99e99dec735b9d0edc22e2c500161afc4b04de66cdedbffa31fd08bb5eff545383d6d0c5edef5fa5e72505028987feaf32ad15962f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ab317a89a648129b3d0f7c2c4943fbb1bd202c1e9e62b1003d6da1dab7008ff370951d5800592aa8e70a693054525a356422b54cfb0976fc5c9baf36236932e8dfa7f0309232255;
        #1
        $finish();
    end
endmodule
