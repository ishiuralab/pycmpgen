module testbench();
    reg [18:0] src0;
    reg [18:0] src1;
    reg [18:0] src2;
    reg [18:0] src3;
    reg [18:0] src4;
    reg [18:0] src5;
    reg [18:0] src6;
    reg [18:0] src7;
    reg [18:0] src8;
    reg [18:0] src9;
    reg [18:0] src10;
    reg [18:0] src11;
    reg [18:0] src12;
    reg [18:0] src13;
    reg [18:0] src14;
    reg [18:0] src15;
    reg [18:0] src16;
    reg [18:0] src17;
    reg [18:0] src18;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a79467fbee7bc66dbc2d463dcbde2af764e34371faf53241f1457caf7952dd37703f10ec0eaf230ab8cc3d3c9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c47d0f1eaef751a57e64de8e1f96f450459dc55ce6f5dde4af43775673df0fe7aaace9fcf565345e2719ac8ad2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e385fa4efd821ce13cc4c9850d0155e3264e762f8c952434c7723d1362e26eda94fafcf1e49645ff9a6c1f947;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb100369d04003e54699eaa629a61a546b01e6af2bde3cd4ed674ab8f602d0229625274b8e26bed755faf746837;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93cff74c56b1c053b1b1556a6c88f4a5ad08c212960b620b14d50dda1ab707aba80b916e1a0d961951d33ca8be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42b1713eb36a5f0072f6a86749a33f1fc083a6b28ee980c013cf0160a407cb0671045a5574578637e558f0889a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a5114e6ebb52bbbc264236b999a1d99c995c3dcf6b9be1731df7c4b5e2856d11b1c8281061968d416fac64b13;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ae88f43b91d5c7f49e658ca3974a87332ed6cd45daceb8ddd44083ba41aff8ef6ff9715f71384793c00e7e369;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a1d18e46bbe62ab569c9bd078b2907eb355f696ba45c35624172ea3796382cdc46a14e6eb1c76e781efd9d1da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8e8118804e664474614588865f1022748f44fe9992ec4589d0a33c2d5c014696c1eb08c99df30d2c564f2dbae9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9143cfe32665b2405dcc1c0ca9e09e32269b440aa360947b507f760b63ba2a242139b9f4c65dc4ce105db59651;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1244e58420f90c1315da0ef0784daa2c9ec7b886de51a01a14212b9bba14de00240df2085c836a9777ee7d151e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h39b22ef5c292bf09367175142873cd5fbeb5f4b65b95f7f8c7ebee46729f72dbacaf9dedae9a8210caf48f75d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hae04c0f8d4978abf8c1ee25114d75a643da90ff1203c7cee8e5d00ae0f39b575879c2f7caed0be177e048de32e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118f2aa8e24331c7f1afa91ee47ff5dfcf9a565f4186b255f55ad35f123e60ca405321fdd68286494f96beaf098;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab2e1b8683dfa6146b96a480cd1e157fa98f7e25bd5641b1840794251760e3f8486d4547f0fb698ceb6d48ff41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf7432f47947bb463390d1e064cf5bdf54eac42c16edab33e7d6551f3f8cd0d5994715dbf81d723fffadef0c0b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa8d6db9023b0279f26210fcfcdd213789408ec9e0d42d2f6774d5878f6c36f02a06d92dc46f39ccb8fb3ba6a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf3caa772cd387de2720c5dc107e086815811fb8bc474a366706a31f20b022502e9ac303cc3da51c1fcab09bbf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4fa00cf867dd892de60b870ccdd29afa5cb511dd7cfde6f340742f43a6ec16c5429cce3ac7898f049a4189993f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h178eb374dae4bbb4784eb29e8a0c495b59debd19e6f94bbccb0c1f8a9e00f4683da5cd12eee52cbb0083ba3f693;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f2c6fdfc6945aba654eb2ad0614a120c00f9b928dbbf7df93996c1e393a8c100b04e4df5803fda91f12727d8d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1862b12dece7e2ca760aa55f644870accadbd13ae20d152caf0b0c645602020e369187cc192384f09c5985ce86f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h759123854fb5c3359de080e61a26bd27066e0f2420d06d54c9595954a5875eb14b0667200a81d5559981cba87a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aef755a013c490e61eea7274511162be46f27006327079165053a4ae76888421f7b743894f680f49230f03779f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4b7f53cbf9376b3adc1361d7560b46d84502c68a8b1d1902e045d8955ffa67ec6cf0bbf25515a20ebb98ca65d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6eaa601bdc7607bf7325827a4f86dc86ba09920c7a4fd87e1b8a49c5203fe36543415db0321f400e17f05b08c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h146dc65abc93ef6bb6a6b29f9b4b73811a7042606d582ffbf09ec200cfe02512622e8d34329c6f7425ebfcf6411;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hccc09a1634f2cab1a26d4a1c4ac884d8a8a59c9850d4a4d7fa3d2aba2ab90d8e529a02073a3e4bf6418c80f07b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147a0c66cd4f2ed8252702ecde6ad4542971273906ddcc044b5babe7c1175ac57712289f7aa9b756f3cb84913ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf3e77f2e06c7fba30cfe9a4803e8adbb549a8339cc4fdfdbfa1bda4862ea400aff0e71cb85a271adb010e4fb7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be8f23cf9286e2dfdab27e1ff6daf15418a89aea757db8d73f5047ece261f88bb46c674d753dcd2abbe8afc775;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c5f212623a7e1d73d7b2a650d662b654f607e434142e85b416c154f4300082e933ce67f2161218a31f0033f0e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd075dbb7d925f01a495a6b670d82c14de63b6ec4aeb275046b346fafc173d6948669ccc8ea843a7266976c957;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7feecd5081d599790d0547347831f9ed561df29e69ea4ba83f5b4a68a524d313a53be1ed3b3ee0477ef1a3ff2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd9505e923242658103765b880316a3ad7513e1c3ad13af8671d167150b1ee62e96bdb0137ea1e2400da2c5a112;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd7f55ba1bdc8f26c983226fe26ef7596e0747a22be908512730a710a2a855c749aaee7575d693f9e1b0ac37fb0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea7fd52e7f47d9793655b8dc9e1012bbd59bf5df1b60796587c742032a7d1d796d3d5c591e72a36919509cebfd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34f9654b71c5ffa8151585c1ae433bdb0f3d042493d1b539dc8692033800893472f2bd9a39c551f465f6a60bad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1287c0af355ff766b33690d023e7331d1f8e255251bbc805c1321cbe3c017e4648f889bc2b552cc38ae68bb857a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64fd8693f563e43f7d933c0da9347a6094a276e142bc1bb69917fc541b6daba90a4012d25fa2d21bacb6f71469;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9a4e77a49a1b8b1ca1da46ce2bc5601a23f803973e8ba4f1eb3e3a8431df255c7ac5bd090471c58fdb7cacf3ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ee00cef60ea41c960d7764fff5acfa0b77c2f169066231ee8d7293cc6c4e7354198ef3320d2d760c34c2f3d16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c524541e32cc62f8802da8821b6971d21a3fa776c16602193b2aedff21b075896ff7d51f917adb6d2cba282c80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b5ec58d2b2484b6706a85b100417fc45b933778e8e1210d39bf07c4e6de4fbfb0015a25947ef0efddfa651924;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h101835f3484d0a5f36d37dc806234d0e275f6c14f125e8a00d67d731ba53b180575a112da3d403159f268b734a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1415c44c6913cbd164c47351071caf6b52ac9ba908ace2c7227f2e599144fd377caf9cb31106e33e95b25d6ac12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h63287238fa07c2abd18bf488ac00b8adbee9b4a18c6913192b1dce062822d1b043ca3f50491cb08d3ed5de71f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e6fdc633a7ad245266b11df04ebc76ebe0b559629408da052f05560c7cc87896dbacf0b0a2f8b5399ad277c88e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h78c84b80a2e48bea1d6644eef263389e854e7647c9a209925ba81d613486957e119c990910a5f0d9326d613b29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1666bfdecfcd2e8f204f6d83d2fbeb630ed602c2d0e29a222291e640aa199f6fa5f6c0b0840aee9eb27654dcbdb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1931f1903285452af7b170bdd702dcc7c1c59024fafe4f073da03221967627e4781eca8cc87016c32ca6a524b69;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136d3816b19f8bfc66d0a606b8a959ff37a034190a07a1eb4bbbd1c5f3569d3a04a0dbab9cd3a9e173b3ecb6fbc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe8d8508408969440c03f420a6859ca658a4777e4f6e0b396d657bf8388d3a8269fc2d39fa54d5992d94264b68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd285babbc08dd029900a9c93ad0162fb1feb657a67a8b87984f0c76d156d8e29c1f5083a739bf851f1620de3b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h778a53161192339bb9c183042da93320be5b843afdaa5e1db8826bd29bf528d35b02557f72c09e3192b154c06a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd11dc8fe80397950f7bf218ea2f63f925398bcf877d30de82979fea8e6051081241e3cec9440c6db942009c0d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2631e53f106336d42e69c78d7c97ec4098704fa285eeb10c4193d05ad02c05bd8befc55975848853f9398629e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5891831f75b55071025e744499ce01c5b9566eabef2e68027adea386352bedc5382807ae23e48bf67da9f93193;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ee3186f326100f9448661219f1ab8eb74b4c99f1453152f6dc1584dfdf9ce89ab2501701b843b6c6422d1c997a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11e97b69b5786fe0823eac237d807db26731c7d80710a36672acf66e81eb269e506340377702fc214a181621448;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18c4c7f356ac910ff9012d7b35e8be0fbc98995e9e52f93e776a19389a2f90b8ce92dabfb5bb306223a3c815546;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h48791260a0443ca7979748c4dd761c841b66fcacded3682c3a2d42fc4df58cd97031f7683f7a590e55ccb14640;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6eef6b04679793663951e950b930af95c6db2076280577f86b46fa5ea10a46a8c737fd9dae7594b0c6690e0e0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a32800170fe3cddbf99764a73504150ca9d21432df49cb3a26758a15078bb90bd35284db4bf1a021a3da4d9f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h153cb06a7a9370d340427586704471bd76996a3cb431186c3e67a9245bdc0bff9b57316d36b0c6a8884b9cfbd44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163bd2c091a2e4826adbdc1cfb86a84bbdfc712b7a9d754b5c4007cf5ac91e20dedb98bf7535e0c10d2a3986562;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c2908d6d14dcc8fbc3fb6f7cc4d48047dac5a4d1eb4a8151da159a9e6c874f15bfde1d35397101dd0dd645e89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc637d2fd5bfb7d3399e78f0a5ef5f57c57670e17ede148c701a349414852c14861dcdaeae80121dd1805f4f004;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11958258b1d44c92f0174ebf7067b144817ab652ba34bcd5a3ee5924870470e18957b713335f62bbd89b4596948;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c90ce6a0f6a47ad4337274c533791578d04458e8642300a3f0f7f1efac2dabaa38eb8dbe5552ac5ec47ca2b285;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c12f05c5ef97b0219264faf631529faa0a251125a861368e6c8dd0ef6f73b859ef1853e148416f5839fbb5d02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199ab5414815552be0f91c07e2bfe7a08537c10783434e6668963b55838c77cc0429a0d2156884352100cae262;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a912c5a2f122fc81fd2d7dddf6554676f19814e3010925785e665d51f7fac79ed52bc25129b647a4a628d4552;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33373930ce9d75c39a345418bdca2587d9c79a58ab2be5be7f97fc6dad03b6e9d3912a9681beffa26d1a5da8c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17346f31122a2884b189bb494fdeed5cb227011363a5a74430076e08bf687ad23fa2400e4c606930534ee637f9e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba689bc3670b709d60869a923b26d8fe2f4035d559e8ee209eb60d5cf9a1b4bcd1192a28aea1e43fd45a47d311;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7e423388f5d503c4dc4618da06c56335aee6f1b6ade0ebe8bba772be4a6d6f4d9fd5e1e2d2a5fb5570f885d343;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6413f75ab9159e0235b3fdfeef3b6927be46068c474fcadb7121e3142fdf65fcf5807d85c863242dc36fe613aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14145686b20243472859802eb55ee81ce12efc2fcb8028f5627641ffab4278347fc9249b961ac7b2de70f590ac7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdce3478aa29109c52475da50a1a53360380668855bfb1536f1ebb238fb04b1089a6f9c32a2f84c36abbe05cd94;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5a9d25e1f1bf4979d99c63978dd8bf1fdd85e1317a8cb2eeacdeddc60b452629b66ac18a31289ef06adf63282c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fe689b166d3e20aaba03054f64b1e1ae65cf05373d2729196464ffd8ea600e58b867c04dba50b789603d5a19dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f677598cac693e497f81ee899d161512a0ff69a1c886c4490ca364b5bb7a9d105863c0d20291a662088a402ef4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff6e642bf176ad2f466b2c220aaf881de51cf610c4af98270ba5074a70f93ad4f94fd7ea31ae9e87275068400d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b20a6c268a091db741255ae4080e39b627e714e277e1d3e1069bcd10586ea6fbf987a5220e6304e61f186f51ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c25c0a5260a7bd6b23a11f842c51fd42624735016203d7d30067c480999cb768312fcc0e1668cab8754bfbbf5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h126adfab89cabdb107cf48c7f2e8028a17d056cc540fc15badd1b230f16625a58ff0a2ce47aa71aa233a151ff7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hadd695032258e6905d3ca4cf391d7f444ae385a8f06fc5920faae9f15a9f6d58d122892af0beaf56da80838cd5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h715ed48777431dec8a65339cc3fa041f36ac81f90f5d7c9d3b94b3178012b65ee1ea9bd0c8b5501f384f980698;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd0e046f35ac1f12fed066ae93861cbd9906938fbe2956f60b317b2c05b381d0ffd0d9088af6b6c2b05c8b536a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8da076260a9e9592765d8c5ab405f8149109aca73056f370ee3a0f7ad6895fe2c041cf8177ecc0a0a4e2e9a578;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6250a18a77ef404fc91a5450b19d01022648dcc1512779d22e3e3bd107a99a890a3f7aaa4f48ef4856cd795730;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e88523b5ec334acd7cc15675b4ba313def72e052078ea8e81595ff565836d23380d31569f41c945a11e8ac9c32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h38a71d31638545a0229ca6005c89addc81cb34155407d0ad6e27da8233078f0399646bee6aebe5b0fe470ea142;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc9c8532978c9c3be27e25c8d42101f607e2b32abda89da55ccc49016fe9c93ca0d2b3c967cf963ea66b9af8f96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he56f5585739ba05770106820d74b645cd2b159d0d69eb1a553ff0e23a05652e5585bc9e33b737b7336a5ff9732;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d31085f5304dd5f401d977d5f35f93bdc9430cd52f2d4ca8098a3375f4589bba4ba952fdebf976b63de092707;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce148f5cfdc0b71c0f847e4432b3f53aa0d1ddd757e2461ac72f16bfc62d9bae605186b1624421fc655f025076;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'had7bf63a2cb9e88aaf013f209e391dac22a0b4c467ec74ecf11c963b9fb62889cb26a725140650d578d22eac1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159550b0523786b003fc3f0edf2f08c049f167c72776e6ada0fd756bcec5ee1fa6eca2cb7581194b53c5f793af7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h104d7d0371472dc6de82246502ef2af8684c27edff5a36d28bc36fc87b7863ec585c58ad125d49916a4ec83bc3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h840a95747b7e24406ebcb1219f8eef9ae775d7bf66a110828ca13ddac7da7f66366b36a4c0743ad1ac33bac809;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he0b5f9841b4bcab09d43a029402008ae43102b4a27f9131c8f23528ab0b4089ea909058558243d89e937f8aae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5b9abdcaeaa7717046ac3634ab9d6c0c31f3a0777b325aade67011eeb601f001fef8465fd15a29012bce336c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f57c6834db12317f82234faf4a15e6719228c82fb2707f81e5f6685ca053cfeb2d12797a0308332ecdc75ef009;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182c28b08a5bf5bdcb3fe08ea3908ef020c6f18a6334af4b9c434212081ce0df832d4f8a2d44bc5fe57fe90a9bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19b4869fb37445201b168b7a0905c46c0105421ffd9fe7cdb6f537998a7033017bfda2837f5f669e88cb05d9f09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf5dc608523461aa9f428f4c1cd4db4e9fb1955e099c18e2a6fc5ded89bf00e6a4b661463e0de1a7eb1c8687781;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11954305e44e6b23beac290b6abeca0036b998b82acea7671b7ac65adf4545ced49aa02685bc2e7eb02b93fd678;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h185a06b7bd9a489892e5adc7cec27d126b37d354ed73305a6d071980c2a75e61ddc07deb168a713c06bcbb97afa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c928ebef6298d51d85a80b9730f32f00bdd203f5b3ff212589fef866f221592a6f50a24b0e6e9dad2207c1e81b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h103d85807b93b2f62593b7e2456d6b45fc081206e7db75e7085c727b626cc0e2897bb02d5acd19472896019f1ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h235834ff3619140329c0d8c927b2911f9f9e86c6d4c0723abb160d8d648145a1f20de1d07e42c5ae35a15eb6ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h124e19a936772b0aec69a8ebb8c47fa49bb7bc06312ab92b166e3486d703db2aaaa34c1d3c3733d99494521c815;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha396a84f35d40f07a0f1dc74edd23b80ce9437cae2077e6a4d62c331303df7d8f54851ea6628a1e56ed92b6741;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1911f6f9aa3740add394d5852a8e19f0d0f41224d5a34ffc51b5b62c88e5440877b2c8c7717ed116aa5f7d24eb0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9bad99b0ee7a8fbd2e97718d5bf911ab884f0f69cbcb94f022ff81ea7d002bb41f771275a77c26c7138bc95cff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc9986fb71bc5fc82cf2f7453dcf470bcdcad52f27973e8d7caad7894570ed912ac78a949c4bdb5fdc1fc66645a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e723a53801390749de60016a20d8ebf43a8596694135b1ebcd866da0cd118c42bcc2045a99bf7a338a6349c89c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5a9229d07a3f2469fe8eb9cbcdb7236a737aa1dfb5a6e254dd96ac379ea38d5e4fd3d575ffda26f505a97d67b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd929ce59ae99e7d7e9ba01a0ad0d2ad710e4049c2ee9be30a617421dca0c187ee89ac011891d80dfe3a67d30ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1495f8c0c28c8d9af8f6c78efc86b5324e1f3405dbdabbdfe420dbc451c178f39b00d06c8174b8b743a1fab6410;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e0d1d244e6d030a2c069e173ad1f92da8d7329c7d881770896bb37c1ee266c156ff34ad6b1cec366ebe38a3200;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10fda967ec83c1b1cd227b812ceb67423d7da58ce9eaf062fce905f6a017715af6fb429a41f444701d6d7a6ca52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd1df177cec971dea0aafd1a52ea485da0855af66decb818a83f457f103daad0b8934fc470aa04fa290b7bff323;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19b5f71b5cc46181651e974511fc0085e4c95f1423b561193c440079a64d9778c071cfe8a17011ae582ad57137d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d44d0aa5e75b2088779fb34cbc429e5c1ab94d7771adef523ce0d15de22e6ac264291d012fdea2e8d4992f06b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1598ecae4cc07f6b209fb0be97383386aad38b5259c8c1636a1f42b245b3a2652f87a0015ae2c4959e92aa0dfd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h967ab2640bb9d1e5282d51bd76d18bde9bdda650e2c6fc20765bf14a6f8b511afcfd87a66cd1412a5dfd3db146;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h662303e99e989c07ac3cfed8c1dc4b8ff3f877cce0bfad0d7a103e881a6fbde6bedcc878b5e0d04f190f5c672b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h127052966d2cdc459a3f46ce65c084a2c814fec40fdb8195c72d39fa3688bce39fb63fc141c539e008bf7408ce6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he1a091ffd6709f7214d632e20575aa0c53cbb68940c17628d1d9932a46885dc75037b88102e21a8d22a49fc88b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1729c5f0a14056f0ab916ebb147863b1859e912a1edbfa2af51f0dcddd2991d35aafdf5dc9d9185c75db93468c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h184b635ba154a049d6840155d4949b2e372a72b936eedd787dab782ba023ea31344f76dc248bfef2411d7d4868e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h377351b22d2a35dd40de6ca5bc7f9fb8146a952c208d5a86778dca7c7dedfc69a5fde8be047ff796a7d9d09aeb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h48761ff93cac4530968a2227c0675584eeb123d462ca1ff9bb0c3f9d8e2ca1220acbb7ffdd586ce300ef478b3b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b7fff344bb1321166c1de6c95f1f8ccd8bcd9c2109df98dbb42c052c7ff066d137ecb59802cd35c499ca84358c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f11f0f7ab1adffee1c5c2372cf48b51869d9d3484c2d5e9ecbf7b4d9708fa523da0419f4e041c854e70cc18e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11103916d06fc7ceb8164ac7915564ae53bc8a242e20a62635d99b629bd53f2dab83b2205b35df6ab4394882405;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c43a7ffff38099d420db47c79a3e3ab32ac07866719e4bba24777efef4a26dd2439c70381229d5837cdee27dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71fe2f04921f23f6652e5dbe4a290b1289e53ef8bfa107524e523b89671bd16c3556e67047012cc06f9ff1e2f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a5f1ca0ec7fbc2564666a84cfbfeb980217dd7d29604f54298231dd803b1d7a9c6855ac7c62f7a910c56aa3a5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b382bc7ee16f039113218747afa51cdff9f6c305884de9742ffbb1eb2ddf45617fa7c95454521df0f977d445;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9194737c75a3942ffbdf4a7cd7055f7d2662fec1e18879fa85dcb05260d2a5632bc99327c98b9cd445ccf203ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142603ede61d7e89c0996edf9131ce16ddc38a10a94bfc74efe2a53fb249ab81f5902973ddab419492c5e4353e5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93300e98cded53fe3c08c40321566b96bfb5349436168c3226d79c7693391df5b63f578cc78a6c0bf895674e44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h63cfe2b930ce2ea7013533cbb4b02737d8e7ec7a5cfda325e9166fd4d61374c56e01212f963b2cef7905b06157;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eb3ac7fd132d48775f929e61c710b4048652ad63daf7ab6c09e658e87e1e6c14b006e7cd89e324f2ad838b13e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h26168eb3f20c4570c8003e26ee1e6d5c80b10cb259fea2f4fc46a789bf4fd046a75d98d5a3a87f2e2248cc2046;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he32998cb19388e58fd3b9ff14e0167a47feb0a164ca3a4a7d21b13607a46761487e6ae93ee9971803b4848f0a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb3d59436ce27cdd0301bac4aa7ffb9cd27666fbbe5a73ce8fd09d8f748b29e048b364a9a59608e67ed9abddc89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d5d8b7cbfa6f237cabd4446c25b749cda24441ad2a624516ed122741cc7bf22e6c215d2fba89280a6b98504e79;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a8f7cdbc3ed6a9a4f0f28a6195274429a916eb190478efd8be9cace744c4a8c3d75a69fe06374aa5cfee1c6d1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fe2aec34174f36c587cda5df5175245d5799f63063c6d4371d4d30a85bdcc74a2080a9f3e60b6374aff38bf074;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h97aed519cae2b7762102839201b4ef3b87310df06c63537668026b2175c237b0e4a391db505fafffdb49374005;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dfa9cafa668bf532027e8bc3a8814c7f5557392d406b603a5b7a87e58041a4d4f34bdf76cbb42abd454c92c5fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13568be495eebc5bd821fec9bca5ba7167db398cbd4520ad292a34855b39eabf7b6e7734be9bdf6ea0b82c8eaab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3b715d6114bc6b4a25cfddc234b5f0f3070465bd08ada811df9104d4bce182f3deb1f41c08ee345f2c38168c58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb9c910998cc50dd67b7c650e0e0e33721e432d19152fbafc045beb1e55f92803dfc77ca32a0bd8b90bfaeaa865;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h169e1bf0a2b2877a7b34ee5ac3c71492e9266f0bb1f6f03c384b7d0a95e16149d234a406c629e1214ac62bf08;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a87c4755d9bbb964ce9cb98a8d13b548c85363ec80e8285aa79d9c9da6728d50260b427f817de3f8670a3f09c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6cd24da3ecfa12da79cc15217d5c4420b6db2a7ec7ecce97bee668800620688360e832358b43e15a0b70286f88;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1edb0d8a122e00bec0071c048c8bb42a40e8693b3fb27d9fbee1e81309ccf477bee95d0f36fb5c11e08b92ec02e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd844fd4f9379d8b19ce19d9dcebf4b18d5ac70ca4114143ec1654597f6d67ef0d932fb247e2f744d57d273257e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haeca3f7ed296c9a86af4b2a536e814a0db5516d4f07cebceefb1e731a8cb9e205f08c81b1cce338fed6ac44d11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h292c88f439a3eca73edfed4a00d948239de3528ba22a79c038ecd176c5162ed9fa046ca012e2a517bc21d4644d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h824e524a1a1ccd862d7c32b181d1f090765d09998892cd9dae55e4548b85022da292185780335be023ac2954b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13724e0114fbf8a93f2e2f29111381a7464c878a72b045c0337e6743ef33314f013623a8860efdd5cca4cc8db33;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb3efd2147fb9b2da8eedfe4a340bc813fb6ac8a225c603c7a7d60a188293e2fe36f1084daba325a6794dd76f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h60839a78575c5b9bedcaf0c4981ff788b80cf313008eeef364905fed4dffea5ddaab337bcb222a7a09287a88a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c96bc158eee8ee454b287783af54c2c21a8f868f31a196c8ca97f8011ca190e8fa61e488c09ed47eaa4733b1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1709c2e887eac0c12d25d9c9c6705e482c083c0bf85e6ce51c35ea1e1a7b6bbe888a267d7123ee2507f0812f1cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c47477f458612c3572a95b41d8d84a689fa560af673a8b21a7743db75ebd17819f89369322a3371cb9b98cd40b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h153b3f0e1d9b3aa415a6b65575834462c2d854183fec6be3f8dbd7ddad6a9cbb5bd21572cafc9672598367cd2f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10878cfcdef772f29bb6348553750817bd851a5ab1c9be4479960069880b1d3bc0ef6c1a9c788313c00c7c5779a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4d53154b51723469d27ba4c63f3416d816cf8da69e0e3fc236d607c989b313d3e1a43c33ec8c0250b3599b2b80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h194d51af43bc53d9681e40b2ade105ab6bbefba9643469526b42922492ecc43a2284326ddda81d430b0c991019;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h44cd1bdc86636ce011f908a5a0614b9066926dfd5594f521a13d8f7ce65cedc4bff734086b19615855d4a487e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e92e2d6f409036fcecec20cd68bc3492b350296038a161bb899bfdf4a0d22ceb14b05aebac162b38d1a0b92d0c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fcfbe2ec9a10ba0732d99813cf19334ec31f50632c26f3cc53c44bf6902ef0fc077ef8dbf017f03d9d01069417;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a7bbc04105defe72ceb7b2da38708d226588a284f219a230cbfc3bc9105aa737ac81cef5894eabccbbc4df6c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h61f405650cb6cf44698352cb227ea49338aa84adc382ac55d2152f447ee736d03a78f7accfe0055d6842912a34;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd239fdd3a3bbd2c923c73c04666a84f9bb50ebaf2afc6a17a00d70072dd7ee5c23eb1a566775d16dc06579c643;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d2376a145798ba713199d3180b897acb842bfbdb19a866ee1b98fa197cddd26b87136edf63ff119c8b0aeec66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e30635853735afbb11fccb67956976caec5fed88588a7132b11c50845d5d74dc8a5436dcff9efae3c7123a994;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156c57ec2a410d6b360b6fe999f81c18f25201a91feba9a1fbdb0ded6bfe98c2af5968979a254881567c61ad2d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75c3747914ba2bbf1bf2d7d3dc3ae749e69394f2557a07cf56cf3863ff363c09c38c9b1b3004eb695cfc174c64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he81bcdac9810d204f9747a22baa853b25edb3e0f1bd8ad9b0cb3060ed353f14927dd37960b231e826959862f39;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94a9523b628a3998933d8a045999ecd47193770dc1f7fa6a4bbcd4b771532c1bfc1177c365706d221f05115da3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hea017f5d623c9e146af827725dc6002c817877923c6756eed7ed251581750759678a84bc6b77f8a5be68a8be39;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d72c3708219ead1a6cd579bfaa9c3414ca7baba0934ac8c0b69ecd42d6b5cb0e53d0cdad530ecc48e30a64f93;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hded48e5e565de5d28dec0e82463ca7578a0ba786f7f8fd3b3acc4bf79f20b9f30560f9a3e822daa855ca479f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab0d8b92587bc715e394e6b6df4b9c638519d870a41f9185683a9d173c25c686d71d6708c4dca7f4f2a3d74e59;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18468cd1a7dced7515744ddf6121508b8f6fde78f115264354ecbf5106d26f486c1667c98d1db265e118e6d5174;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70a15a74145655feb263789ffc71c99aa87d9ba031ff59177421550dc7d25c1905c0a8ecf193d2ff9d772a318;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbd8b9300e389e7112275241ac2ffbdfb0932deef3be51931dced2bbfe2fbb13b03a1779e3fccd14e1546eddfdc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h188facf477c10c6491b537722ed82670ae8cdd7411016be8f6b333f98d6ce6b331054184b2265654c5ce21af06c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b1c9bdf21de9cd945fb29fc0ea1341af481b441becc2c9fd3d39a650a9f9412c6f2d1041c4c716c45c4928f81f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f46031a8a798b12aa8991a6fc9ba79f0df0109a7278c34774b89049764b9867c13130b529a32d741617d64365;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heab086d2814d5552c811b9c4afad5b2163257ad55294b262ef8124813e82fc59931a71ea468b8a11e4667ba0a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a3d2b29bee891bf8fefd5f5e5fa44ebd57fc447a44c7dfa328f96a6bfbbba71ba2196af9f65733933ce1f2600;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1410374a763952898a69532fd4c4e0c362ef6896671d353f820b0ace29c470d6ba80d91944e0bf023ddc732779d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e494610184fb23c17811f7d17befd063431e0ddd3e7198303f956bc4669e6ad632812d13b1d08d60f394f62364;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf59a9e906b34bd884cc68351de4b55d3884352d3acb4d52a84a1f3c98d317dc2f9255aec143ad57516fc69044;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d2c87df4bcb55b9932266755c9222932493fe0d8751707844165095af29995da47c1ba596ef3a456248bf1b56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bdcf1042ad7df212f340410797a3e5f36708fbb4f01ade0453b90a4e57fca0b7e9de2e7b1f090a473abab1d476;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75995cc6f325122604b1228b7fbe04d946d5cd5a3e9b5cf0727ce0820ac1e70acbc93309a2505e7a8d948febbf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd426dad3f309067a0408e347e4f52dedb5379e2249b92160127885969777b572f51a2fe982f50c9cc515a48bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc451bedc2e6eee407db55fa32606bfc779cdfef0e39e8f0317cc762dc967e6694b88264d8cc76a3abee1ef4d8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fc44c9ba16c1eba2802aaeb45e5a154ea9381bba0f8837db3950f62522669c5e6ed722c11a3eb30238bb85469f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1137a436cc4b53ac50f3771103cf6bdd237dd14b99e0cca823d180d62d0f66c00bfe5939a96e88227cf268f13;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc12a8e7176647f1623f487a9ac757029be4160beb57670f78b3b6ec8629667bc99b8f1ba180c654c443395f44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b381a0552bd961888d8fd17f37c8ed42156adcd59da5f8445d66c5efe0989c819886477fea4b0a2a4d6428a76e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0a1feaa562596d65acaba4ec52476f2c33aca40b1613b239dc27427195155cbb3ce35116cf3b589cad7bae638;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h281513fe60c7517992e550d2a5229c901c4d557656034fbdd66ce56ed40821400d3d86225f83ca646536b9ca50;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5782eb3b0fecdd3fccc16a0037c6025f782d256f2b4ae7101537bcabec58c72c5365acee23b96df99a720a6c5d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34d11a173792a24b94b0acc530003cc61c6b17aaed6a59258e0b602f9ec90c29992126fb09f77d4f4f2d5e7125;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e4c738eef81c3924b5f2aa485666980f5958fdae3acd11132de7d607e645b7ab7ac8820600e48f2cfc51a961e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e21d7cb0de697cc1d2c59b061fa9673a39c74104fc12c8e634f392477438c4c2f8e36a56d81c2f52ba5ed94e0c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5e86130a14661a5754847ca257d849a093cf241613618506e35ce64f3ecc60368430b14c47a6e347d6dca3784;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8e76e1525e86f23fbb4e0b32b9b16bd14e5d6edadc5f1a914cb682d9c9a5660ec375f4c4f199a1dcd2c54166a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haca2c7abb022fe7bd91d8905421195be5e775471d3cdc775236443ca1416ba9009316e2ea61a5798da631cd42f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdc88bd66ecf563b583229e7a039135ed7ff55ce7ef4b18dc1ee4ad08d30035c72f666097682a83f7b43ee7513a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba99a0b00b57435755aaa7269ccaa48b162df992c7c5d43dd6ba8b574e31ae843ec9fa11dfa35b492b0653be69;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4abf0a7eebb6148bdaab3460bd3f517dd4cd916cd70e2cf5becec1b1b4155dd5c640e55c3630f1bef7d2ea7a23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he069fb587d305b83a2eb545d0416f70f37ad36094fe3e0f68bc95c38c57ee423a9c3031165bbf7f6ce64718fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28ffefe048445475f07ab6e22ac33c38e02d7da48151ed2f732d07dd783a579c620856b1d14912ae5311e607a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2de00422cc20bc88847c898fefd6eb59912dbae890cbf5425df74e6cb020f465ae5c7f57dfee8aa55ba33ae67d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfdd4e69f360472bf28da6b28e591934407d9236d0537fd886971b360f38cbfe4636ae7446d7d3728e9d229aa1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hac135ff577d74f2aa43db3133974b18f0df15c7e75fea2d4ea8a78625c8f062513d2cb1319fef2e87af0f823ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4742934817fd40e981dc54b7cd3e923d478f99132654e97274a9a662332e0077c8b01d19461a868cc07c62dc78;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ffa1de4e47b085211744f964b8bdda7e359f7657563fd057d3007771278c38756a66723d8f13be1f9c14203f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2eb45e01f6b240805d1bc61fdc3fefca04f13e68addb39a78f16ed50f6601bdb73e86e5d896ef561b9bd668d98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfd1d5fed3fb040e6d8b67b76d46d33ddf87729f15c9a01767177997e61edaa498e681bf2da82025293c9b84974;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33c390846c1c6088e6103d86c3b9f37414d84edc815b98d51ab5cbd3f80e4665709c9e946f44ca4654f6f28940;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h564aa40a5d6ff6c069e27717bfc00e7c338d252d736886e7b35c7a01040471ec66ce48ac44715f0bc5b29fda49;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98df64ec751b599b7a0b743bb545620fc96e70730f42393c15983f874acc83ab2d310e65b8406535de6408aec6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h77de490b825a5799092b6f10ae56de41a1f98b50d80f11dbbc8ff0206c87bc9f670bb35fb1b8a20fa794b7b6e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128fd611a1e38c6e382cbf9826a8de20e1fc764d1e528078e4825f581a65216a33c0c19cc9995ac1ebe11ae0e68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3b01d05249b303d2b3b29c77377db805ff825d92121d2edc21069a52ee5e392eae7a6053a249c5c1382e535d40;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h111edfcaf331148fba865954e5653889111454e1e1ba60535b90e7e7aef6218bc3cfdd317e2a9c479d3e41a80a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f5345701306fb5b534087f6b8f50e2c8bbf32784ee28d4205b57657976cbe173ce532ca89de0deccc5d9650e47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h327d06d4bc23d3e9a65e7d26dd443d6351de394ab0ab4de146dcc3d14d07e7f543d5e530d01f75378e849482eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h456ead1f2ff544783d83d4849c454c197ebf6145a689b8928da0eb2dbe9cf8f05641831d71fda41ad1ae275314;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cccd87f53593b9359b7c591a985e128cb605f41916d95fbbe26f2857713c82eb15a93f887aa8dc71fa6c7edd02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb97cb78f24e7c1d55a4d2319c1e1c5d5345b047eff061bab662a731d495b70c87ea9900ba8f2228a8357d4da0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h194ebf3f1aaf1327f88fe6a9d7102c1ccbaf02593a983ad1afb7429987e03a1f72a9c7518e6c11db0fbd29ce044;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb1dd7810975ce0ecd34c0956fdfc68cc96288a7bd5a5b4ee9a368c67fa532667799b287ce7badcf46a3588a9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f32b6c0df4aa30ed15e44f780251ded72322dd681d46b62623324de6a305513ee007ce4a08ffdd370fd886d334;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b62744c956353c2686311511595b49dd6eba13a4d7cd9624467455075774255059443e13d2ae3f491f454138a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h495b003bd3c61fde180f25d0385c94c187c3e0896c0c1e65779c8efe563a7789e1e42458d206e5f974e3450abc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h347929f770962ecbd51a9adefff46f30db1801d08397bec47b9a43b514e8f1ff08d74d6ad844222106aecbec7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e0ea59aaa12bcc3f082926f40b9c9572be5fc460564fc371c1f59a6b9a526d3df535774e5c8ddcd1ce2a895555;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h688bbec7b2be01e9f8edaf38fb6fd233d6a938874279c392c08481395c4bfc6c2e146c49ecd0a2da725c5bbad2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1289c5043e703528898a8ed7ea3762f354b047bd050eb60427f65682c8c401f2544510512c9d469c3f102c46d1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e064a6e619e39ec2f446d3a93ccb27fb96025d63c6586be7ae57d881c0d954aa3ab4026051c7d6c960bd7a25e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116964864252db237508b7dfcfe8d23666aca302c4cb2e0232fd2ec65911eb3c94e626308e84f9ae9efa9575d8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f1e2b076d39dd517ba85ea0819f99cbbe5c4bb22a7d4a646386091ba174eab9f47c5c33e4c9fc114e8108a838f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d32fc8c14963175dfcfe25e7eab25c083978e156f5793332e8346ebcc24b41d9e09acab3aee48e95cfa8428d1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c07132c6dae7e8193f3bb4edcab561844e4fdab91a24fc9ed1ee1a61eee2ab050fc84f07eeefbee62d026f7b04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ca324ed06aeb842621fbe2db8478711157e1fb0ffcf7be69353b6f5de0db1dec9da205514ee97774bf2c1e4c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a47ee7a25d3485f8b30c0fe3aaf0623e2cf9bde2daf9095cccd63806907e10cfab247bdf6ca5ec611f103a0efd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7db473193c2f2abcd1323c94973c9ab9e4ceb11fccb5c30f396f3f58ca7942a2ed24bbf116dd728d69635db11d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf8c0622ff067d7c85b602545ca21ceb656fc91e726ab944438b5caced27e40e5c3f61e086658a037fd7c126ff1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h846ef90cf8f077baf233058cd39eef91f88844f6d97cb5b3b55abecb8c5df71caa370e53aa418d57d9d9f239f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1da5d1697802db49f04e1abce68924e93194ff89a24ad7c51b3043983438b4f0d8b68e4328e6819331ac7165a98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e3df006bb577f24161e0233e2902b7726bf694b48ccdceaf21ec894d615e8d5c8f7d32b3cbb74ba2521b597d28;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h325571a6ddd37e93c03552ceac8b766e0afd714475b381215acb2661541204a5909fdb2ce0a138b616c799b2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d965a0516fd97f240cfd3e8fe75ec541e07c839f7a9f23dffc1c5f8ff8651794950de614ef6dec1fcdb2034f59;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd708df47fa8edc5c436ec146c32f0eb2a676a7774d1b741092c728d29c3b239286256640e69152fb9ccce48060;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h323440786a4810f89805275f31d3f4727521af3e92195680bf05fb2e8c42c145ded4d0abe39a8444abf1e38bc2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h489ad4d6ec168980897dd5f30300ddbd3eb0848bfff33daa4d9f42dad3a71902676666bda4e16cebe8e27586f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc2dc3d812d3fc3a3b0e0307550eb9cf9ae3d60e6d5a7e4116f97518ac97920811c838c38dc542e1aa6d57463bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1978d6ebb6fbc48176673f982ce92386799f4b640b09b5c9de1c632022c9255656455787f4e829ccd53e3b8a063;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35b983e0e6cabb822437be092dd865ddf1ac9ba3c526d51a123581b95f2adc64e12eba68be1fc8aff8b6ae5f4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e058973989cca683fa93b94489d240996486513c00588af030531890ddfcfdf4257a333fa2f120c118c81fa1a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h119df5c8e8d75c796c377aeeddd99237cec8203869690cb97a7b60913d88896de7ae9185e436472dcb373de947d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf14ffb6e055befe89d8aad61b33637847c1b15bf1d7a76bce990c649ebb1402abcdb7abf4b4a34bb585248303;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd4187e27caad3004d6fcd8674eb96ab7e194cb7db4fba1ccd9f849875310301e42ec2b80d7597726dfdf1d853a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h197f30f18076edf16d7c863366e71fad7cf79b0af11402afbe177826bf44906b06dc4b2fdf91c5bce2c75263730;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b04ffe98e66b05d3f85a234aefec7cd00a5e9c9e4e67b6fa90eb12336bb224e6ad98a3a2258d4a626054092e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d189c2ded01059cab5dbb0177f5d73458e9436742123baf7c000dfac1f4bdbf59801e83a86d90e1fa83bbd9ace;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca6a1d613bb82fccbbf9ec1cd158986dc8d907a0156ae927f20a144e6729a25e85b1819fa4e82082d1f6e49085;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf29b46602129eed81e924ba01c35b034270ec1076275e344ecd92b982ffada5acaf1336b8c3977d8e74ff1f40;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11b7335cd4e3a896082e9030a615042dbe50520492cdb8a51757364bc944d01b87364f4d0665bde73607c7c60ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e97010d384a57382621aa601261bec317c20a4e40bd081243335cc936b4dd08bd902239b91eaf9c70b29bc8e8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19b3d3ee76fcbbcfae1068a27765a8b38ee30f9fe0d9f5e98cfc2addc9db095820df576b83a838e2b6e6c5e35b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189155b099ab1691770db2c45bfb168cd1ac8635cab033e91cd92e15e083ee29e699179346f3a4d7fd015043d06;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae69752efe36b540f4514f02a62b13da43e4adc94d9df32327e7006d7971aeb39ac99039d044e5072bbf8f89af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6481277f2f494894e9f133d0c039cec6ebcacecf2c9d7da665b9ddbbed3df78a2fbb2db597bfd36f4421b270c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf66db461bcd7d67d6e8d58840076ec1ffa1c7114c1bf31e76d20fdae91a4bcacddf4fe1b094d23210b9088030c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f48f79fca65de72e3ffac8ad019a90291b11368671ca254f2f2a68c79218b61b607da80c345df77a5812049e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1639c35760bf0ec864fb9ab78a15a535c1d6f3a141c173523c4d592f06009c72b65b54fdb8885a1219cf1459e7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d281469c77a72ac3457b9af0e6fd8ca499786a051ba7da8efb5288f2cb7a25145a99b58c60583d845df0b9d5c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h779ba738c6074b4c047e4a2582f7f68d9136a67deba118e83276f79ca477dfc3de346bb53ab2db0d8fd9044cf8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a285ccceae18b6770c1a8ebc6fa32ec66183bb99143a4272416382997ad5d20bd863bab24266456dd4f80afdbd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcbd2c3ae26ad51bf9e0df3994b2f6c3467760da74522453d945bbdbefffa46bb4334c6ffd360d97ee8f2532d95;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7bf3d037ec1c53fbd789e43ddd0ae21670f5c0836030f80acb3a8ccd27a250b77dad8ef62f79628a04d86b2fee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hde2fde9c3daa3473eb49dab7c917f35dea843cb076e95cb7deceadb22f7277931a49bef24f833ff1e3f82a0fcb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h30a8f6f24d1a4ba2c324a148a97091981cda624f5dc3b447930e679394d579c427702dd16651f30fc32ec286f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h183fd5d95ee905b3bc3417e2edf37e2cf54a9137543ff4a29bfa6a6d0dc52aeba731778276b05fc4f634130edd5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1894fa10c6800e2e5f8f54c0ef335793aa53c3dcb4b8ed4177e932c2dda7524502254cdadb44ffb0f9e6f662204;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h86ebbf51183fa4f49165338747e895b2cb57df626a9f73f053e41403179b613ca50e259fb5f4f32f8ded199433;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc45ad02d0080930951398fa754f75ecf3bed22ab2511146f923754bd3363ec4f9b5b011e797451217ca5cf60b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11b136ae73e1bf95f9fac9e17ef067186014ede668e135ad2597ecfeec9a1415cd97f03b2753d7e97a35a5f2fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5e4f1defeed37b52f9259d938bc5aac47d6207383e81ff689ea2c38d20d54f1e818948c048c0218c678be6c7b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hced6b729c8221137eaca7ba65d989254141709efd95c7682d4c4e5deb9fad9d3c51690948111f0ed8f9bd84241;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19172b4ea516c93cb368a68a9105647f35d84a390bd651b698cbc711478be11881c86b170dad841beea8e9ea84b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d27fdb0d8d0beacc4e63b78f43c1daf7301a0745b1bc8385ee3c31507900debf1c316f6efcac9d405cbcd05f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h139ad241b4cc726014290fe8c56544596f5c7a9500b9f514d7fefd8281bb6464608c959daad063c1ca059c739e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h145105c625f270bf90ecb734c27880e5f1c3b25189ae70111c5c6516e3f324c8fa0ae03f017bf759e3b87f0b4a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d643eac34032a7f8fdcb6826571b55821729d689ac1ff53ff3b4815461c58c6ac042ff95170ad446d67af33994;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13896db9e2dfc03cf2ff21dd0cdb321c3672c4a54b3e5c2eee2833b45cdcd264bbe62cbde1f85785383eb371c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122737fac61923497f72557d770f6339548d46131f0d59ee7fa24544126f0554abd106340c8f0deeaf1a93c06e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he70f48de82c36325970a98d80ee32943dee376294257a51c0f4203e593248c3175389d050ef5948ca673a7efc3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc94a670100145ecd97016cf6d7718576781361f7da1a5ec9f87c606846052cb4d5e3150e769ad5cb3ad19ad46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1188cff1deb0c2ce7d27ad9c48cad76c99c4088ddf5d01eae7bc5a0c558e3c06684d9470c4c49a0ad7b38a89ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107d6eea8cca361c842871c6eaa6ad32735caf3c304bd5a6e84bd647dd7b8bdb8dc4f3dd76af52532b5ab64cab8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b32328eb1f980284345137fb21b4f1c873ff4c45d11668372f951504e6dabb9a7749eac85fb324fcc459f06c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b1e8324d91ebe2d8cc6b3906aa541ef5df468a78a585702228b28971e6f0c3d376d0a2c538e9f4b84c78b88597;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb156e331e2013a19e0eed67c677ea9c0a6f3c67fadda08146ab7d79ef854dc99cde8c112ff0f531622c2b921c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13bfab4a6b9c057abed196bd272b190f3191a3c135163e7d276090128fc4e31649a26c5acaa0e2183b5280d0426;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42c0a2f4f3467d4a55baf3249524ea42538c10f98c5470efac0d3ad089dd366da7a4bb9c7465a0830e9e741094;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11eee33da34e6079f5d3154f44f4cea0cffdce813d0c07a966dd70f3d317091ed40ed9fab5884d4de5c362560ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h188fe56a4882db6bd766741f274db5deb01ab75aa43410cb9c411ebbfb0c5dc97eb34270d3c0900624832caa6b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134aef350bdf2ad89564287c3ee21863e401e1b96dba6432599942828e2a0b36a4d0de7ef9b20330532235e7883;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he9ab1fe238e84e04f4122ce79e2018a7e669926e045ea142b322f9cc055f0add6501f21caefefffd66b4eac6e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e2b80894313487ef1b42c6aa8badaf7e814e913ed6bffdcc8b78d120a69c77adf5327504bec5661d7cde9741f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a4d4eee50726d064498979369d108d1b051e000fa03ed33736eefb637914d90be4ec73c7a4d2bb588f434df7e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10ed62cfb65c5857b8ebd9939a75f5ae477ff0722eeed477991078f7dd932529d1059fb9c0fee00dcc7afb6f98d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10def9ba6b6f8bf61a67352dbeea5b2576da9b3c05cd62afc18dcf69bf491b3c213e13e4f2cdf74a3f0fd33bd96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3407c4d1c775d0f6cd5874b71990596971e084b3c69077d3b2b29128e4839f7f8d4d27fcc0a61723d875332c29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hadcf3d638b01bffa01ab17d03f4e2ac58f363fe9d03adca090f003624c9b9067012f2df1a96a1cdab9fb140625;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb834f9491ad61034429c1ce04646f6b554aa23d7f659275a8bbbcd705d8246c6188649970a9e96593389735259;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h139ba49dd91a7108648fdb23bd15af859bd095bf46ca24a6c9ca38a56396b87402850b0fc25f58caa447c0b61e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h194dd47a19eec998b96c0f3b7fb3505383ffae7f6476a36b220e5eced82556ab95f27b4902b420de7730f538ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc69f65568d65798c097d90ad88f5a04ef0321fcebf7fd313d3e06bfb82fd5b0d5d47d435ebea8638c4050fadd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a7f23107815be3f6e2b9b133e2d925cd5c8a738aebef5cb8eb7cc22cc4b1bc9be0529f6adc3886c6dabbbb6f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h962813423593572b5e6696290ad36e10f658e1ad101397ac166581bec881f9b4beb7fdb880c4307f1cafa67138;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dce855399e6d24cfd62c3413aa119fe7258920bab43685e5b4565fb32bf9938b9b33a6add4df79d837d1493515;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a24fc48ff96a400a04f5f5abd7eddd8cd8c1702b642a3d81d26205831a18b6fd76b3442efa2a22bb3172b76bdb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h38a4d2df53fae0bbdf1f0025e96192e07c88e69a2057b0464c63c22a909a807603cb90639872dfd6394907c5c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbffed96a2c76628229893ab34a7bab99cf16538f1a246b86b7904567cbc57e5e980d0250b804c8cf2ef34a1c19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h939eb8bb6ca6851122ad167d850edeb6cba09280ca515e63d8d3d4c37710d59f1adc008bdd55b2e25f94e3630c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h135018139337a34d7d74675f6965688af40658dbcd327e6b4dbc1a89abc621c73c967c28134cc2ce8ea1a80979d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ca9b35ae4ee2bd3fd8f546916a79f476c79dcaa94b8da97b70aa63de96b9f11e31c642290dd1b835916c0f309;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha541a6e019d8b58cfcad39e285e31a9e22584c4b7f6ea52219fc4dc538af59247693f1df9f6165e3ef93efa80a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1887926bb6c6655ec19ecbcb9c401904cae6243524492dd0b49a2a81f9377288c02896a2c2a1aff0efffeebd4c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he4cb830e9ce99f108dcf9fded4b74780eeebaabbc589b540290ab16c3496fbf4e69da2d77b998729b097dcfd20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee64806c8fd634dc0fdb4ad81e9516626bb759a4e7d252aacf1cb4b7777f17183dca013e41a7a6351c80258678;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ee101ba870a28f3ac9550dc47c1f08a280046bc164b86715029dc89d1d77f21faa4a57dcf8cfd53588331165c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h111d5cfee50e6f09c3f8c8ec313d38f41a3106287cfe10f21bd111babdb8290aa028527de5e3b93da3f5f8b2a17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f5ffd523b6b53dc720824e103c186a28c74ebe2e6ee090dd8e9ef7d423fd98f0c7f7a4b333edb1099c109e72ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71c5cbd9be44a8961ec7380551277b8584caf27ffbc464e3c7bc0d8a0b0ca49480cda925a9356185ddf6829c74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e486fbaa05646f24a2939560606aa4419f3899010df67bb8f9c5e13d11f047e375c852980fb6ff0c1af6f4d0ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab3e027722b0fcab4fffe1c134d367704f0f5244044f14159c7e2f6a0a817bda8386eb16d0fcc67aa06d353b4a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e2f6d4f1649db0aa630a9340573d680c028ee103112e335aa0dc804eeb1c1e406b05647c13fd7562c78083a43b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5be68852fb6161c4de6a79a6fc279d01af420499953c1570598e26013d40fad1c1fb98889c64690dd9bc11f4d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10ed4a27b000874b24d6ccf7e5ea60a3a82ba33fc178b2a9901ef00915c1018bd12ea6c2afd2e4758644840ce6d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heef3fd4391ad33536561b3bc60da7450816e17ad690db6101a18a8a107e6058ccfbab7eb96b9b0bf1a8b4ee17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ccc5c726f76b20dab62957f92246b16e781c744b81a0fd4e25ae73a3b309a2e2e08b42519228fdecb82644ee1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1511c0f77b62fcf6002a40eb51ca70a0d3908777d6720f44290ef72457c045b3cab8612895e70b181f6e7075d74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a75a7a97a73e3b3dabadf65e0f622949e70ca3d013225255f5f1e59d1e3aa63922c740270f57c6ce2f1a9cb68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa3c4522598502e176e78a2b15b7bdfe6739753ccc5de03ad23fb20311b066554972da7179852326892624ab7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18309dada0adfbea87503d236dee1612c272b9742a09156279d60565ba602fe21aa320b9a80ff5868f354b73bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h697105103e076b5597913569ec9c95bcfb6155c28582182c3e3149a0e871c28758c570f24051f6049753fa0477;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he1d0e154c6332dadac11ac38217e11d0497b1882bc77cf1cdd241516a54ad3a9518b2504c503fca27bee9fb70b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33a58a165f98548afad60e08f259c048c2f06b077436b4eee0ef738f9c0a7c4cc2d2002b1267d5ca9226016e19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae52518e2e22ee55e3a6453c9b4a7e7cd4ab69577ba0066c034f371d380232a1dd8d62abb43527061fb54ff8ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd7fcdb79aafa4c29d8588c8e18c56beb8861462c4ac504e2b3711a2638ec0f7c9d11a7734537b7361fc777cc20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19cd620e57a0a7ff9ce133ff5fe27f69d53afe04deb52bbb6a38db605042d73b79299e968eaae234bd60d7d2b15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13b817766cd95155dbbbbc964441f2acf580fe1e310d8767517743a5e034048f39cb67db6361b0ce95b8d9bb10;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d93be5e75698b69b9281b0810dbb6d9c243b9ed0b8e15db4ad7d970f9defee147b0c6da82eb686208aa60f94f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h100af21f88bc992330bdb3bc4118c13e449fb92f72f8cc84f5f547d41879621546141f3648f93253442bf7e7e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3545d23b5a7cae2b1a34e565e94c700dbe9140b26bfd94babbbd0a9b82e3039aea401deb3bf5c65335cf375cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha336335edb6a9be0e96e40ecf33964b40c72ba207eb363ae04e61e03109907a829a0614f4b3d580a98c8d814dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d56bfe4c15aed269b98104c49002974e3b44305edc7241b8f78cb3d26eb29aca3286710c10924ffc7356bc61a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29589b8d577fad0aac3578cfb9d0cd827689852f6fd3ff46480e9303598b033b51f50931db3fdc6fb85efed16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa86b3394c6068b3f3e487d17f5e2e330962ac8ae6810a59574c48ea450f379fa82c9ae7fc841046b82534473f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16531de4140aef46705c494985be8d099b07ba425ab39fb6798de8eb1b6a1ec6acb6626739fc14dcf95d6f85086;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed241c6f003f5e76c53baf73c0b6683bc05e2cec8a999afff1a4b7eee39085ca7a2b3999da26ded659b77adcfb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ce379e90b6c37bcb15d7ab36198b13697a0ea90391ad2fe2a27507951b83660e913fb6cdb7c4e146cd05bf5bf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d350f9b4730bf7ed03f1deacdd3fc6581109379045159a5bd59149cc5fcffcb59244178bea414680ffc3d25b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1528e2d4633110d40377fbcc67749e013fac4404b44d3aeff2b406d164b6847fb1c01a3459f7db8655b892a65a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c6b59e19f26e3736704a336dd7f8fd28fe224b516dab281695db275f7a051ca88a192c21f4a5c9f336691fe61d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c232432103222425312a3708d9d264cff8017c83373651d0edd1d2b5970457cd5728076e614d6d43cbd81ac273;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e1b2947357a945105bda7ede041d1026068d1f0680c5f2eca44ccb2293d1a39ac47885922c6f9ca0579aac48b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5cebc3250324e5752ad9785c9d90d22f2b5099d981167e845de0fda36f2b8ebbb43f125062cd354cd0e530041d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7822ac1f99a19a5ebf31813756b9ca31084677a61a94846b7aead4a2aeab1aa4bea5b57f06a8afdcc3904956f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7e16de5a00c83c2a9d3693fc1051c2b7d85e68cbab01bfb475d95c48d5b7969c63e83de901084220b110e24af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bc513821524960a7032dcbb41d629320e7cc15e4b746c0cd17a22883765fc16d65caac6ae7b303f0f3d6f513f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b3eef0e7d5a7796fdda55a144a3c505b205054cf27055a2c42b2814024aed99ed892e0f4cd5815435ed1eda22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba2c0ca4aa3417ade4417918ed3630f30bd28e7c66fff77885b077ae5aff2886611f32e31dbfc6455a5e0dbafb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2669af1ecc96b69b7ecfa0837895b375fcee26fdd65ba90a42ee6b1f0aafafe4527b2403685328a11ff051020;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffe0502d4eb9474adc8e93f44a7fad1773a3982c4975934832304e473a5fff676ec5d209ec240bf86f6fcbffce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1147fb90d709b7a736b0e52d10fecd9deba3acd93ad053c414e98bb18ca4fe51ded270e11fee5ca1ef92c6b15b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h645242ea173874b778e4ca995860f889a98f3f61c85c8fd90a9ed2c14e4edb027618f8fc7f870f38b81c50a36;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h111c2515c032ab93b2bdaa4c67a0713916703acaac0841bffad0d983bc49803cfa41e31dd06db2c826fb92c9a27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1303b2b6c3b335e38f00f892bfa54e112ab7cabc22fc797990debc847eaedfc544c468df6d500fa46d7a00b307a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8012212b6179f14afbfbd74061e0a2d5dacc759ecaeb525136021708c07343cdfd5345bdfa16804cac03553750;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8456249643df0f8cebda0cf2ec0fd0310421a71ff621433c8d1d3eb48e936258afb5789605d3dfb13054688034;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3825a028202cb33a97ccd44cc17cc3cbf5ae49e5d7b381fc4d6876455f241a3842b8fa9acd0869030951bc25ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h166ad0c4a302d3736bfea4b4ef7f57be86a3413b5014ccc31a45575ec9435e84379daa02702b8acde9b756a17a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13d351f381d5b947a9b85bffdb7866adacaf480329bb835f8d979a443b32380500b66d6130825019c42b0bc3a12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf84b7556f0c853eb98faed44bfb29fa61e16170ea06575fa36085b2c4707986ab34308556186ec7c9d23bb1f06;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf9f23fcb04b9b69344d295c851a84f1ab2d3004b6b429faeb6c85e1f21ab54ba867fbdfda7f690b257839a0d22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13472e1d82c0822d3ddc7e2fa7e0ffd7ced2ee5301956130e75b48ac4e1ea38334bf32b5f952107700f5452c7b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c1f60e9702870f008be1e6dd1da9862ef5f229729bbdb42211df5176fb80008702983df91b179946da3ac33f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h642c584d38c6f6de76b58d9209cb2ab304bea7dc6610fb867d83d07122ef84f74bf686c37336eaac5be4282df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a21d08a1f0ff530e62d793243bb5c7c968a4bedb2cf38deec7b76079307b1c8c195526ba2989f5c43f91b9bf1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14952b1668e36a6303a73e982274a37e0e09eadb6e79156a610a987f3b2b8e3d52ea02039721b9111e66dbfb972;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136d6f1edb6a4eb78f9f323fd3c049251617c5ffd5ea7a6f28beada49de618866dbd9bbbcb8f6e32cd3e245311e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf46e14164fcb0ba35399ca78ca88a190b1bcd1830bf735dec43019c0e0219479c2c9014c8dc744f74c9952f6b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d7dbfbfe2370bbf88499c6015d18565a531526c66c393f2bb2c2319fe5f2d77aa794da872a4c27ec90d96dc12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd9482bee02c225801baac7b8b4db8dcf45886c4187656529b89793881896ddb505cee82d9c4fb0b7185ad88f78;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h68fa5f6734be3a33744037b80aa156ed69087e59a51ff911157ded3c8aa85d78a4bc3cb0314ea7dfce73a9e90a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b936628478efee2430e074cf7044a7199e41bf770e4741ae6143ffb700545b3a60e1198e1d87cf834197238d58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12e395dd60c7d9ef9ce98375722028290b79944c428deeb3b69564b858e02973438c36fe63ed59b56c3f417825c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b91d2f9f3999393fd8f07c6a7c9efc6e398ca3df1d0da41a1415a2e0d55c472e039fdfb6a9a5893a78aa31851;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8219e9634c7607aea0b88ffc6d720fde0d0654e90858cd7c3b99bd9780a03f71dd720209715ea1e42f6e7bc6de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12d69fa9c15e10a6b2cde66001563349e07ae7adb97fcfad6e065ba3d27ede0d08dab5c3d2fcd7b548d69d05fa0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41cdf810f07c6a14510afa558737ce6e54542fd99a92cf3b0f8f2049a4ab877888b0410274760b99c3f2a6567;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf5bca56a45545feef89b83bce390c3e320ff75f2b5460cb03d39b521d6c31ecff9090b00da80ec9532e9d029c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a4a50c519e53cdfe368e53145b677ccf5ba8f2701af2b97c2753396cf025d7567c049240ca919d6e663b1d8ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4ce98cc7138525178f145487b149358bf302fa1bf28fcb4588af5614ce729a9a575c80a5fa88c8440711f8fcaf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda0ab9d425a254444e45d5d8f3343430832e8d9e19c4a4b090b2ef871a50abe1409af303385ecee5403dae694e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h533690088e61a1daa4f34c1ffe1863071be378ab31b76b63148d4222f81adf13e5157fd1494ec440370829c20c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd27af0aebd34ca0ee3a2ef352d0d4a5fb79e12a9484a866a7383e64f0eab00a1e22657e1a89ec2332897b4f99;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1ba49e97b80fcb30addfeabd46ca477b154cc8adcb310d664cbf9fca3bc2997fc0c30a303dad6ad342c37c79a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147c230f1435b16d8fffc629c78eeee1dba209dd36256e5340352de3c7cd2916d3eb1dd93a308f76ab425c9db68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c78a0568ffdf9f5b6f945df56fc7a0d9eed36f90ea01e2ab8604da4676ebdbea6eca8b3bbb29a7ff53518026b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121459ae59b18f3167d5d4d4e261ce790316147000c28161ccff0c468c767583c4a82427483e1a89efb38e8ed9f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc1fde74b7097647880713617eae6d511f450af29a617d0844d9aa5ef59f0774ffab1fe19f702810f74ed03233b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10bc5a9b0d030776fe17556ed00fa0c4f58bbf1b0d197368c13bda76cafe82b9df9e064dec9e93cf09092ec5e06;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12682dbf368e7cf56eae98ed10e4275f557617d801fa525dd390686c7f0ba002df65b1165efbcea89cb1bd5fdb8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c92ed9248796a797388a6e39e6c9dd15809bf9a20f5e96baef91ba13817eb41832df3ebf765d3135f2a664e3d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b7f099d55dfed44e72caebd0db247a0f6c0ad5507e29e65aed531be6fb2fbc434fd162405f0c050a60687ba67;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a1d0ea473f03368e75a8c2fcceb4f5b993d4b68d786949079bff7b33331b154f6b7c1bcad26d57d1785aa116b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ccbd15c35d39e3adea50459d3fbadce9336270d473f082a3bded6d5e0e9af7ba9a3dd24a38fbc4a4c68262640e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e365c568de39e1f2a5d682c4359dfc67217806258784fae45f89227c7ace6a0b6f914185e76cc2f7d189f2b255;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e6556a4b23eeca9362ca09ec5c0fe70611b64e2104455f0445b31aec82f982922605a8633f3c59b284a83fbcec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he79520a515fc99eae7871f599929e9ed07235b1943d70f460331b1f027391c217acdf899a0315898d230782bff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h67e8e8c77d8a320928adcd3ec89dc6d50daf6813a56170177c4f884a8dd116843c7859e8ee2a3cb36f685afbb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b28365a7be17098246d09f745f8d8ee43726b913a6833f8332645382b4ae48b1e4b61090f066c771149726d5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17ff489c543028ba7f48f9939ee91fb3d5fc4450b1d4777b2bad6ad7a082908498ed56a33b11466dcee6306c14;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128346fdc4005e7b3caccc82dd51a72accf19f9712fc45b21bf69248c3108a3d85b7d6356c701e9b69f4c4e960f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12cbad78bcfec184e9923eda71ee69b6f742c6644da9079ce305e05cf6b7b3423e090928b32641f792d6775081f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha09a4f7c12ba359895a8fb4a99e9bb032fe1d8498fc6bb8ebb7b64a4d2fc93c1eb032ff878b1dc955503f5bf6c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8fba18ca78f1fc5c8af3c2d7eca760f4ae6de7c52b87582e1477a969a1155cf5fa86943682832aee745ec7e02a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb437095353ef10309cf4038385f909509053e44206e41266b06a70b550ffda1239c712c359ec4bce0522e0ee66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h76708575735c4ddd213d5320899de65224a13789111d00802f3c4034fa83198984b9b182b13b266fdaf813ba64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb04dba1981de98d91cf2731eb15a4b8a0210810f823af3cbc4195fa6fce08611cf192f55a24be0195e82a4d46a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4cb7d81231555e72c1079f5073aacf3ae8998bbef8ba17d6df5d44f47297e56f8f831eddbaa0523b5f6e8c70cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e3b2feb5fba28ad76857387a75cef788ede76688f8e4964505f46dfeded218e0c9c194ac19bfe5fb330c9bdc55;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11fe9d89e50dbbd3bed7017bcd6153d4ec7fde6b63c50e4c37bb08027235ba097399467b73950e891965ec2da7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1573cb9054b1331327fdc2a7d13fc9ffd226f4c0f647a87490e06f8df4a65fad5190ca53c7855bcc81864cc795a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af02e276ef702a8b10c51e9ba89be01f16b79a9565017ad380e40085754b35dd73ba7af67cd27ad6778ea8369a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1074464d41d5b9348a48785c551534430b6869e23cdf0e2b79df91e25a6d168d0a9f09e3d1a172d9b877b9c5c76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c907636053b1defe3d6627c32831e60547331cc778a5347aad732f2e79a5919e747fcc4226cdc5f003e24cb60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd4fe5073188cb213d5343964eb256a558b797286fe39f21bc41c24b83d8f09a90aa7d182862270b5db890a8bb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1acceb3e86108227bdc193db85e6f4a2840176669c9f88717699243a4e33dcb67541ccd18668af576cf7d415fd5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h152bcf1d652e53860e50ac7ca0f611e770ce9291d39aab7cde1373f4714b3e4286ff5f9c586e97e69abddf43e2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h141c5095425ecf97b8a01aefb86376a3ae43b5c8cee40bcf6db6ca3e1c884aae7e12cc1b8599ee1facedca5265;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a8f99b4c2a99aaeca805869a94fba3a4dd60d6c6f67a438add3399a476041b20aee91b9646829bb7ca3279385e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7d5a7bd429f49fc81624290cb1bdc5abce58d3a8095fa756fdefbeb5b9b05bf2746f09f5a8256ad214e602220a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h61c14e0ead6cdf4fc994f9b5b7e4fb597a64cbba340524adcde3a41f41bd1e26fa504dde2febae6a52b36d107a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h262fe54fdc92e220b949e9a5d85ad8ca8366e4dccfb471bc9ae054f3fe3e3aca686c39e001cc5314920c5dedf9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h124891df3c0968a837a1a4be2f53da79a3c872ad765fd4f7643439b217a2a02e4b63294d33418852f2baef58fce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd9587a32bf1fc505b13e30dae012d41da0c4f8f13ee29b37080384e5f7cf2fbeaa475a5461897b2cdf9a5a25d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c35ce42be88c439122c3ee59402d29c7b26f45981c19f16ce8adcd5918d7f1765c76f09ed15ae5e481f43c2776;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1397bdaae7c59011c5b5684eecc99c424720cc1119b86181c617f954ecea179bddc5297c47fc1c8b275d20e7712;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e0c657b70b15539c3d652a8e0818904e259866968fd00c86c41a57debe84f81120dbf579abb82fc02be3f04da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1471454b9dadace529578df46ba9e8a43492651c22e531d4c09f4efc754001e3660bcb5cc4c8779a76828250ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16fa2aaa33cdbb7a2ce67e92c5a63dced3050d7b62a9c464582e5b2f6f58554488e94b391e0f76c59123b00b0ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha2343b5d8b52e17e5d4096c4e9f16ae8c70ce41eb634b8856e53deb54fdc96d472168b69b34057f256f66119ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17fac33faf32e5a94046b1824cc31d50ed1f72e82493b672995cf5272e40d594b3e1cf0edc56ec93fc4b2923ccd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb338bd37db5b295f0c72d784221faa9203d7e4ed816673254c0932ea01fe3a386dcf506a5c78790c826e04af0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc878c40445b55931aae0a8ac7dc0bd09f7b9e25cd236427a393c6825c8143334f152da543fbcf9147f5fc5e9c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h91d87c5bcfbac16c20af5a1d01d8fb54ce94cb6a23225d68ac8c5f0b59c679b05a8eff2738d8ecc958862d4cf8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fbdfa9650c1941e29a88bcea99b2aebd8ed1d898dc6dfa201abf7e304e099d8205e34136db9dd211527d1b947f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8f9c901bb9c5ce3663f201da3c960abe04147d98d13bc0fd3bc8983fa7441bde5c39a9da6411ee8364814136;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h85ccea2a4502859ce6d2f17e91e64abe5614ace42623755ddf253cf12f9c58166920b27b1f63314bfc4c25ae2d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199de3f93006f6c134d9fedaf3823251cd2664f80e028296cc71d60fa10920dbfbd4c28c239d3f6a7ef45b16435;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c9a33762190996e48182bc72dacf864e2ba35296b98662e7235770388a0fe96724af36f749ab1feedcdc541ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h158b522c7d8a72f35f88504acc6bd4c892bf4982b530ebec54a996d85344381e7fd1f7b5552a3c17ffdd6b06b86;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be5500f121a987f57571a38cf7e2cb9f46a6c99b280fb635a7001f3b24fa6d1cd1cd84f156a4904265ecfba335;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c646ad86190ec9d0e9842eed7443f05b25eef14a4e370fd359ee856dd062e418956a4167a969eff1308273610;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h106fd1ab5342e05734963686f197330fb647815920c123200da2610c237a7596f792377a8644c66fd5972b98c5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1952829b2b77ac59625212729e6f1f0df2a4a601561c867cf53a4a4d4a69b42826e33c7b400cefd4ec758af5f5a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e61e4a0925f6e8ef4d8d50864b70fc65b94e740770dac2c3697097ee9da6f4220cc7354e8a4bc767cdd1c750e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h256a0241a2b6e500d412fbeced92ba777bdeffd794d7ff685d375a7ca5e5fca4600e83c7a8f109af6afdeee542;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4f7a54a6caaeed369d49ad99a730ef9cf1333fdedc4283439f503fa5a86c1816f4d0365fc7b06a9688d2a247b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90174d596b6a34a97c97b051f4a09168737622f29f81a70b73e54bb79d904f09d34347601ead0edf2b4ed83132;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3a7b21b414a79bb5046bc65cb7a9f231279368a848459785c4aef4da995e44cb612280868593d983e7f7d3052c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h383eff2cb94efe31a2361e29ebc9841cf9d1df1d207a70e3bf2b919cca097ecc06132af87b7fba2abea482a762;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1afa092ddfc2ea269f30cfe29431e7e63bdff678a288c3cb46bd6fc5f33a35704400f3b074333f51697c7a3752c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16b944b2d8cbddf15c0d4996f9021366fc50f1ecb0720fc94c21419b4f83f45e27fdc1bef698821f7009ced32e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d0416aad370aeee0bcca6b27646a677d58305c953ffe690d53816d2ce302941a506cd4d8e9840705050ca46fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a86272bd92fe3afc8dd970043e7aaa81f90c4ce875461cf01d8df37423ed1e2b0b7f7ea7019f70666d2d1ba4c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d3f1cb2deec7144186ebc6c424f816d9919d9014d2acee1f783bb96b6fcda22abee5c3909a0691a01d7fc0b7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16dfa0be2c2da099b8df3b74eff538a25e9cc3e3555878820b2a1eef5f88b31236cddbc22687e448534f157723e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d76217aa095d931093ac7173187649094010e6501ce23f53f296d0244333e6a1aaf138eb8eb2b927d712a147e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fd3e18ac3faed97a1b8edff3b9201695eba9c4152804c779cbfc349e4866b758b2c670ad4571f88a05cf993fc6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha2723bc2d00de24b86b47b0ebac619e0f57563e90480fd795f1301f93bbad1099dc6849be958b716a047c29d04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfcb255055116bf0bc6507e7383f29654d6ef09bc2a5ce065dd9be5de5e721b3be50fdf3137be4f4edf131885f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19e2c7e5f03683a4ec040221badca9d44c1cabad12be39ba22da542578802e8f81cdc04a0bb267f16bfa187ee6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd6c62e33f0504d00f264734bc8e337736cdadd28c117c52f5cda5163dde254565f4e695a1bfd23052232af9d70;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c6f89ccb4fd5a014dcc825a31372cb941411aba43d47ac51f6a425f7e6832714f230f8401a619b390ed7b3b5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h712ba302baf9e0c1bf66820af7f4356124ad30b85b7f15dee695ecea39c3f62938c02dbac128bbd9d1f2649be8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c5359e25110f50ab2ae667ad5bc3475fdbd444298beb075090a9e6349cb0cf08cec6b3bc6b3568044ca0d57a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfad6a382541f56991252df234eaad215507af00d31bc8fd220d309470b18682bebf1b08ba7b091e95bab869788;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hac1d1193fcf039f5f89f302302b7d79f19496d607f8512f5b26e3f4c2a13a7f2fb9aae1fdec0cd832800dcb866;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d3938ccf10e0487833d075daf56465ab25842806237b97edca16cbe13e626c6b11db06a7b4597b63c8cc288781;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7514d2043f69e324048db3a8ff532af2a6da46ecdee9d68814a5eb55ac9e19da214bacc0665690cb31d0385857;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d22061f24178de158065075836fda08e85c91b77c2c42a3fabbe81a6ee085bb96a39b4cb5a0b7cc453ccacd6ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b670b90a15f8b4825b180145e49cc15af04d9afd2b613ca04545acebd129d3788afd601ede1a436d3291c3fad1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1245678b55354ecabe6b570feaebbb6c8df3390bfa06e311d7a7bde254c898fe6392f261f7a87982d02d05fa2fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec6eccf70ff2ba50d647d088433fb46133c86c900c792c160af0b7481d9121c99d142512647b1a18f57f44ed14;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ded2a16cd0794e349063a7b22bcddb4c4f2efbe98420641ee16bb6135b765fa6b07fd64734c2f3a68d80a31d77;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b9f4e8edb8b76a8f7290e6b89b8b103823c4273f3822dd6ef35863ca477f6537d3720b362610f795ac83a26159;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h668a94446832bcec469948bd2d041308f1de4848d43a0e0f45ad0dd2046f67beb7886a3c42b875e538b4a68a62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1406a4b9bec0d05ec28da488f2357979340f2a82711f679cde3d5d6292f13618ff8b695e7c677fca2b7b99f2a24;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h103eb2a405bd96852b651090c4f1480be273900cf8dc824b68cda38f4936b442c1e2bc5f18b45656231f19dfc6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d4761ac17f47f5b4b532e92f5c773a6dd61cb7db94f5ae19d2487856921536c8e963575f8edfac3e5886a0ab38;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fe91aa6a9c446527491b53cbb2aa30894eeb0f693de65647912164aec5a8ea7b6cab236268c7964e7462e49d72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195da09ef566f4009de46bcb347553cb9c92f95cef27f8edd6d9c5da46e26d0ffc07483a6fbe32a644693f8c8ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf72cc6849523679bcd68ed797805362a83c3163a4fb49e9be8219dd14b742c55f7d2829799f58b439738a4e00d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h597ad2b4e05b2ca120a67691c346d0e4bd1b671ae28747d8c18112a2e16ad73dad31daba835991952b3f9f51e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1deae67ef9887faaa2d4ad19a5e5708a139d801c61f6c07562913ac88e8bc747ad2aa89942ec2f06421ee80ea17;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1620010e91195cf941cbb9a9c188de96ffe84ec043b44dc29a7b6b2fe43e83f50a9c4321f1c808162e34a6c464a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f52224bb013479449390ef6a34e93be0c9a366b853b25e18593a3fd08c45e0d4df3cafa208ba5a8907787a0c1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h331b3f2067d0b47989b5c37adefd4719a7be918b5df49b55cdd5c6601fcd28e40c225890617d7abf0cc75cbee0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h304fb152d93b46a2a09f2916984f63076b22cf30ff3b52163d34e135bb0c4c973b02f37cbc989e22ed84be679b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e301305a73d8d09acc8e240842d01e9823a4289f255aff41917d326a648260b2c286bf345c283454ce2c0ae15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6e0736d5e6c72de2a59bdf9e9be599b6b05659e0749c1b5e10a87712f57dc4417e1e1010a932dd66bf208f1603;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h66ee85478c82eb546acc36883846934d58fbb8b6b218d5bda83c37141b12b28046160085f92fc8d91032194db5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'habf98b06e5728783bf4ec073ebf319f722377563fd143a462c228b4106d79b330e3a94b2bcdd7030dfe7a634eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15e6664cbfa3522065e0fc61b827a587ad2452834dca37582219423061485e8b0c767ba151ad46f885ebe1ee429;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h92cb183eba2c57be9d503f800a40b80aee221228dca6075af4fdec4bb19f81cab90100fa57fdab13a381a18423;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e28b39bbb1a76241cd8e1f1ef6e2154a7f6b05e2624fb6123d83ae16a05267829cc5ef6ed70542f57ca580c52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7fb831d581e587a48a70df592f23553a78368e8ef0847bdf8c6c7b4e3fea95f6c14d45dfba51f7640b001443c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1088141485dc6e339dd9933e4f604594660ff047f374c55ff533b54cadfae6b7ed0a6eb499c8c466412c07f7ad1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he2b49c9a31114c9ca18e2a61656c4f2e8d14f59ec5aec42a94420c4b6f7377f5852fb571578d98856832c4e64f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1edfdbf635945d6ec679c192135086094d449e94a73e13392b1386f57b93f3650d86c2d62b05c985147fe7c81e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e755f2f0a61c7c5a1c016b21e1dc369dec8424943be23559735f419fc0a6e38d12a5d747e7db3b42fb86a1e612;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7eab5f407e6f61750296da49fa770949b41c736fbf38ae31b0219ca14470596347b75b4e19872a919bc05bb672;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb2dd008a75ec63933cff1ee28aec82199ecd39c55b81c018674934af636dceb4f6013dd3a411e1bc6891bc6d11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc6a6bf1312054aa05a08fedb3ea6841c1eb19bd971629c0409b45beb5b0b920e1f50dc1131b7402c75b4fa4ee1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h185932d61c2ab7d9c4f23d3689f0e6762d92facc2e0ca3e286462be6fed4144efed068b71a9e200a326d8becb3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94c3676de8a0df13d530de564f2ccd43af0ca83ad77559a83aeb6d71d803d66288f3f9855ae2fa95a74166f11b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10f552afee286c148b9961295ad753e6cabb44c3146c404398d78015a0978c803a3a4c2a5732459cf210a66c908;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a828888e2a0cd35b434e06bd4f626a7a5ce597d77802954a26db98abebd507b2e9d192625b05b350b91d4a12f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a4f21b5a4513c2d109acb83e084e9e634cfc024a83705fc2df2d117762ac3c4fbc2b68912ae3041f24580bdbd3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118b5c5344d799780d2c9d48c19827ee72122dca93889a3dbba5d95566665902d01a2a5012394a4f1b8b6e1cd74;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b203c750b357660b90fed90ebc9ed40e4eabe96affa0bb7debc5085c9149b6d0ab8ecf2338ea90899e41eb7a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hde957bfffef8249b3209c8d436d727d4c1d3aa210c9e31e46eb4169b0016486c1ebbc27f2dbf93a309c209a456;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64fb1abad95d6b5a13b3bef60aa7af0cc623b27e92f8a2c8aa631cdd82871342dbbaf22aaa5fb1d94f332e409e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd95e6139b8cf29a91f0900fe9e25ddf3d8d8b677d2c1b1a525db8fbb6505df87e307d8c0a12cf35d9cbd3be7e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha566a971c4ad5cd814f5178e51db03e6b103c4234402433a313f37a5d8558e01bc5f93dbc6874b1e79b61c9290;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51291515cfb64733c36bc44117de5ba37fd7ca54536e87a08bd9af86415a632a06a58184ed8076e661fcc9238e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h62b2b85c04ae0dd1e1badfe6c9e49d38b89a760572f7ada67712c3e13d8a81569e403c914d33c246f268616d8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd27e48aec791d76c2a0d495c47f2de28badbb7062b6f4ab655b4377b4126d56573f31763ee737d1a34a8d81b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f8242efa201c87068e4a153303640c6b46ddbca301e6381527dca0dace0887dfa30b01a1f868468d9b7c8c2c1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hccdb98704a3917c1041ab349d7d10834a44a63956b9151167f70a166c81e6bd552ea81f2179dd19f8a00876451;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h608855c9064575237b0fd51b774d57a550580d82bbbbc97809c2765c5b6675f02c70e5aa984405ac644016b9bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb6be9a25d969c145192cd8dfa08f08b5730461129169ca6ba23f1dc608c37f74431a6c0251d4307365045e09b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a727481c34ad2ab67568dc5864e81e4073cae8ae4758a56cb2439949a9030457a507019cce0d0a777d539cbfc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fab34232164abd5fffb582cd9539acaeeb3209517721ad5e802679f0ad7fa3d698bf12fdeea8e44f96ffe4314;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10c77cdacd828fd9219a0d0272dfea6550ef354fb66c8984424cc470a1fd1d6000f1e5cac6f6e2f9f59bb90fe38;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b7fe2897820c9a80ef07fee242f028e19b5f14c1c663e1419a403a8b42d6331c59e43ec240635d5d3d2d193659;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10584f71ac811d8c76c3f600f66d71e90a2adc3fd4265c38ace94ad4450f80ee8ab161778255a0203a880d48b1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fac6b5ff898e57183b2487443644d21655d00cb04fb8a8044693bbfd7fe70df9e06431dfde3333c84dbc91b32d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c973fcb3af7220494256b31f5b8ea4307d2f4f0015eb6a724337f6a5d61ef985d6425707a8d62d2054433bfb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c7b433f0cd3c25be41513ca8b9ab51ee7ea0983c5735c05000fcf4991e23da25755da6be572a46f86f7ff1d3e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h110da78d3b9cab9585ecc12776336b909d4cbaddf9da2b0392c3cd266b9f6b0c0c4850c54a5d32c39db8ffbb631;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e57d467571461bc98f49406e4e08cf0b9fa7a689516019d7cb93b74893f1bd739db3808262f5c8a6e827ce0a6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hccd4cc99d62a3d14ee7e012c1da971b0a68faec80a5794a87fb278250cc6e8c50832c8c3b26be35a56ead560bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88d7bc868fa446eae9ec3974e79d1119efd77478b46c9b8315cfda86f402e0b8ce7f754aabb4c91bea58ee0b93;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a7630b90a4952e28a92240af0429c9e6e8458708c55ccb1400a6782b410bcd7eec4ae3f8c0d96c03c092357ebf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9def53e217ff8658a58bf670adf0731b547f08ae76db3eedd6a6a402906740ad262c34d01facdea516f4c08162;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h97910441624bfd32a90625dc5245e5eb4a67a2bfaf362e4958f2cd3879b9d9d9d8eb3e66828fbb55f834d6397c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4aa1e62b9148d646167355eeeeef883759ed36719528de6dd28696bdae4a6645fe16d55eb0bcc175c3e8ead805;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h920c06425a4831cabb590623f76da3344975574f87a32cb5f5b8fc9ec512f4350c24b87e39faca9783f1cff015;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35d5c275ecf115986d30a59dd97ee5089135fd9ed6f095aa0a8b8706660810bcd0bda8b0e0f3bd7c9a57e36b6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe69cba7ce69a3bf570febbbd3021a20fa62ebdd2132c09112394bc63269d04c1dd3f806d21b0a942487090429;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h108a297e3fc4c70889ef1e3dc5fbb219ed5d83de02ac5773e4ee414356d46d96d63c401f6d033286bd85d44da7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb88a6943a4b3fbf5b363a781125cadaf9270a7c068857c4889e542cd0a639a30667867d5a2b0ee1ffdf9bff605;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ce34ad0224373c4e6fadd0aebcc91780e2f74ba05526644fa1f7a2c02e144fdc1459b98c5aa694a46a5df2fca5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a3be7f966cc41c7562ec147e0c89fa559c346412c827f35103e43b774d6335507173c0091ec1d0500537008bd5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94afab8109ef833b4c2b6faa5abeed9faa2faf734be365b8a04b05cbd18fe5fd81c3ae30eef2d17ec65eed33f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6f135f16b4c77e8be36bdcad41b7ba2b484f87056854c8f90563deedf1cbbfb355af6c051161b678f2b99b6cc6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7af802ed74aa501164e17f21b05bf0003288eade3042fa8ab451d4162d63ede48eac2c322ac6b7d46c198757dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8bc303b560df51e1af8872c60d779e9e716f1dfe40c69b39e2b132aa2e066b52dfa84a72586d2ae220563e0386;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f362f04c3d1db327b6d38ae2d6c40314d575044a7d6ff58dddece06e7e1bd73af1e5ac6b91fc06c084db335237;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he44aab497b818fd5c40fd65a1070c37efe323319db8ea7e2188b25f04db8a0046fb620a434603d42ff6627f83d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b0c448da913152527b52757b83486556e4439878fdd02410664a6bc6190b251e9ae92742af39e76a9930b52f87;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c892ec3276670962ce8e6d7d8aad0a7de0b01675c22e5c27e279632acafdf4ee12c6699ebb96ae1ece67745d6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1263df53c66bed846241b881ce965487e2d7185e22c3f15f5a6d18647cafd0c4481580d7d8f36da4a8fc986769c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5fc42a019bbd5c99f1726bfed07305d35d3ef8e1a5fb8ee0f2d613c95bb2afd422a0cac7da5306815a8b0f480;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f756b1189be05da9afbbc40f43cfe35032a214e364498039e681a5796f9bd18225939ce707816d22fe2fd0ab86;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d96fa38494cac8c1258db3063c4a07f3f09fa504aeddac40d991d395e409cc91a4ad909c7e9fe093a4b0bfdd54;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfb4b10f2a1e0bbf1719e61f2d3afaacd57f9751012ccf564bf65a1adc7edc1bf1e0ddd479437f3c61aef7785df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5545a109d14bab9c89d9724ee408b95946c9c8d5f15dbb910d743cebe7884fe2fdc05eb576a752bcc13776a78d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bbfd99ac0117479f56547f53493febbe0a07d65b5b248aefc3c75aab9caf1d7546b89af9c9cc4cb5770df9ddcf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19054464d5baf488d96f854acefe28745a89de628f42b29073ce0692007f5ec8df7165640a120ff3e42248fa252;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f9aa030f1f38f990bad35618899270a466c653e0fd9fa74a18cada1a1f7d9aac2409c9274566b3c4fd94ea15c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h31a9ea73c40609e77fda7ed324e4e856c3d805b52c2adaa13b04f14726e9d0637cf3d8bd0dfdf28009e02ec8eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4198567b36ceae76af88ed6242b8f9fa2a726e3ad707a8dfc8ce0819b2cafd8da59ebf684766c6fb38728869da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h62f59e510a9f512496b5e7d9b9aed14c90ebc048a41605c3ba82f17934514b38af77133c1d2100df72dc22e2ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h194fd74206afcf157087c0b250d317e7821555e31db672b01c6a9a994908f1188d52014a84357e7d83e94bd39a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ec8785ab6cd255e1818fdc6c53857924e5f5674b9dd843c45473b81c2dfc885468482c9a91fe3009e9ba069e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d58085da182bbfd29c2ad862c984c12447949a1b5e2bfa5edbe62785c0cdbebc938559188482c716f240132a01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35a9df4969e06b8ad2ded51774036db0f4737c7de69d1e489e27c2d1f84dabaa9ba4f21d76ad9d679369d1cae6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha36e64161127dd882213ad50dad84e1650ae35de151197bf115d1eadededb6cae0ba4719434704b42afd525b16;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h178ac16e690935fa3f270b8b4fe77845bb808c37df7ba654d1b34e1f6a2e10f0df289b001d10df1b68abd9955f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha6451008affde804bbe4ef1785b40dc794e6205a3afa081f413f5ca7f979bfeda1ca460d3964cb9548c1a2ebc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a2320adfb9cd8159365893eb425bd7120f47709c111943eab5b5c3237a7e61252a535fb120cfd25a20852028c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10306c9c1ede9c47cea9a44860b4ff93b94019877952eecd0be37ce0358870c2f69e13014ae9885277c1b01a5f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ce46a6830b1da565dcdf83efa545a6af12eca91cb630ba635ea4b43cd22cdf0843f74ae1f0c49cac1ba5d1734d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f22deeaa4635b81c94a067648b56126b9ec54d9ed1c87382bfea3038413d164438e438f582081815a3c04b853;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he621537eaba6232efc772240bbe3467d6b95206e40bb7bdec0e412a8d02614c4d99352e649467cfc8b3e2e7614;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df948e263c5fd38e67656ed5efe3729946b0547b4f5c01b309ef47a5f1acccecd48f2946b6d93eb9b33e9ec2f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15078456d46d730871dc533020c6770776ea8d383b9fe2dee7ff55be191caa63c30f7b85276da1d7550ad60da87;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14fd5899dcfc57c5ecaf1d5ecfec43ec2f372a8d230a9f7891bb17330c576b553df21cbd8e28f658c02063b6a5a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5be9d75828abfbcf87387030faafcaa908ae3e4dc19bb5d5082b81576701346b4b6a1c70b57949b32127c69018;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a4f9a40af31510dcd98b80996a8d2babcde899e39d9d1d9bdb2b6907ece167765b2b96b4d88d0b4cacfdafc7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h936e820cd4ee30774753f154b1f6c6264f9b91ccb02a41fae377129960557c4de0cf7d3114013b5d44f1588f5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee88109e05b13fa55380dbd372adebc71bedf089d8892103ffb51c05175548282d14a7b1f885a27144fae9a08d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18e1c7de72bfeca567b06696ae64f9014529930f17bbaf0e4799c1150d097cd1b817e70f912a50aade9676a6244;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1818d0c0563a330d43692def547ec32ee6bc530c7e2eec80ac7840f017d6b7a687231eb7b9631199a77186fa138;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d68c5ee02dfed198ec6674f58609bc68da75d80ef2722080b4a31339bb8f33f1de36fd06277c01982dbe253699;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce20f9364a1b88915bc2705759b09ee179b77fcb3896d1fab594757daff3b371e27febe48959cbb2c08f6f34a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8961fb1117d3bb8b4dc3690a938452c7791cf58803d582913a6b2a9fdf3a6228a8c3f27b6647d9e9b0f19d2e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13b90f850117acdb968cc0358fdb8ae34c0c3d8ecd1b9c219890806bbf3bcbe2a3bdcb7f2616de60f456d9993a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1050cb336693e2ad6005b59d41eacdb69e1b7b2e36245fdd218d02f4bccb5167180efbecd624c2293bdea3260cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf0c1721bf446ffdc9ae4095647072668424573e0846548dcf7ef95d91953b7625b99226160a92cd70714a77d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae124a61a79b0ad30ffe5d108c5da48ad909f6f53efae0dc8b6c0e645d86c4d6053be81a12347e77b7e74f2487;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8e0147e947abf203a203013b1dc1df14d829df17fb07b8437a1d5d4d8f63063a5c94155b671ff7d8a72d26cc6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10bc23dc4cb737dc88dc94ef939bd7d296a2828eaa830e3a7efeeb520d1bca687cb82358bde300d35fe42ac7bdb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cfbcfb60046acee230d38d81fbb15f59b07518e22103d460ef5b574cd3b66e097761b0fc5c15ba19cac1ed715d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4d016b8abe9260d3e4aa0906813f6a029cd2071e9d75643d82bdb41d4a34a6c333b23264deaaa66065e3a20538;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb09bf97f7f4191509a0e2c11907f4f168584a2f0a2848dcd840f523c74fdc548b40b77248d006ead753c2bc0bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19b13563bb4f6eccd0c6a16d340119e145bb07180d3c2e1f9e6b2d13176eafafa8537fbff89b26eec31b8c779ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b60eac22f63eee3a7ab5d31db72469b00c6ce4a81f02500256878b48780bcd85acd0f67f2488210d2600fdebdf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f70831911ba3bab31484eab4517a63cff4dde96d5259fa023ea54b0911fb98fc336e0b5324926fce1ed6eb2406;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9d45d1ed60596fe51536cb901ad3751297c3c689f8440388b21cbe6699e651b65114d7beb1554964309f1f012;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d3979df1f65e067521a993039eb0df1a7dae44fa1535f5bdd3feead5b16a1b741eb9756866b6782c06ac3c5c84;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h651b94e3dfc94914e89540b75a5c3270ae3265fcc4132bdb8eef82e1f029260acd14c0123e5aacbbcf6952b2f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h398c2fcf22f8387627d62a75c648fe0e77031c7738733de7351ea2b516ab2181b2f95b4e958c167c7dee83703f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3a9088b4018f6cea713eb526245666984fb7efda849ad9bec59de597c452677cc6ef2a3db4cdfa32aafa56b206;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2527cbdafa0a294256f49a556e7d2c09439c5842de99d6e550e1b72d4bc28a7ce16fd3bae53a6ac358c9f3dd56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae790436e3d8191d62d7ca1ed2a816d8f2412d1a400b4bbaeea238c6b37e34cf58b799d11d465fad0029aae033;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he77b36b7258e39d0840d78bec1ae0f2be6c1dfeedb889b1b6f2e65827411afe60ae2982ed82001a9bbb21d1806;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5cd1b7c029cb5ded443611cad7d0f3cd7daa11810c33aeeca5a7823356c3ee1761e13b68acdfc4aa99fb47d00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1138eaf5d0c734f446fdb1d45a21bf154da272657c787d9b536e9072d4b89e85791782fbfaa8c599e1cb94d5934;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bc5b0f769553faff00b37ada95880061c4adbe2df05a360e6400952c818c7710b8b7270193a5da0dea1891c961;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132810f4b59d5eb8fe979c5b5b4b2dbfd9c66f5a0c3e37c7a43e071071fc9253eec14e88fdfae1a1fa906c66585;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h420a97085a42d4cadcd0ecc022c547e4024494921811b05f218d57b96fd7f7ccc3c59cf07e18df690a02dd0975;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h171e7a08ab7534349be9e8b3c8a6ae489f5a187ce0b63006b0ca5e3863d1f901c4f4312880846d36b64b5e0d802;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b05b5e2222d1b1df308cf36ef34cfeb3a18597adb3ac37ce21b949e52f00226310c2df1005e7728aa5698b14ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a0bc16da3791c8dd6f0ae7a0aaf11a1d9adc503550929a8c7683f21805d452b710bb136e58ba2ae644de1da51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156f2624300aec73d82bb2961d6b1bde83945f18f5fcd9093a4f99df00ad33aab13c222415f57b779bce2979745;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2963580dc7ca720a53beecea34b9dc2a850c4752d8ea52e57af226ef83bda9d3470183979a1eb36549ad0c235;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca8428717f17daf6bd117bd830e4716950073ec44a4fadb49e9ddc3ee078b2feae75174a0e276c9baa3f0e65a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e924401d8a921dfb733d5c032fd6382e47464a02849c41ca6e8479ba720314eb07e4deb3787ad3be381f6e8009;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6f31a1c3264d297c4abaab68f2306103c1f353c3ce55af8652991f3f04d01f5f7a61d97a4179435e2759c59e40;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d6abce38b2f9431854aec6a93ccf6accc0fcc20279725a022df1918e3705fa43a50dd6fece419522ddb18aab2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcedcbf4233672d3316a7ff223fd77374dfb856108bec03d0e5d8d494cecfc77b22e7296422ffdc26f42ae47b72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h65588ae263bb613ee86e5436a81aeefb1ef4b39624139aae7a2349cb7e96d4a29378bdd121a6953a2f2f693cb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h148ce722bbbbb5492932d52d379e17d9fe7945070be6110573d733e2f2451437ac9c3c3183060745612e6bbb873;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c419f18d40f221922d7f23fb78e0f1831fa8906bd41f5e29b18cd187936520b8fb9d59fefa7e39edd6c18ce89c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haefe0dce5f08ea2e82a57c9a33473b3ccd1eef5cf3fa3ab9ef24e7a69e4ccec9b7863dd7ec7842fd933f0c5e9a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf31b8dc1a632120fe43a6c09aeddad309898eb132606d1c25b895bba650f12e6c6345d75a97b38b53921d7460c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c3b8883dd745e57efbeec090550c4ba1023e63b5545fe7039a350f955df742a7dab3c4c9e4ae72764fcad24a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19e9882c1ce9e0469a5e69c06ee25fe59fe8ff5e2e24d47a5ce7d3bb8db9b09ef775224e8e58aba1bd470836474;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37adeb6fefc7058b64adc696046ae78058495c99170f104e17b2e64c61c51f3b1400144f616c95d910a2197b40;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc06da5bbff641af8666d2590bc25afd676cb879b26504a3b14dcf16fbe02228d71bd0c0583322abbd262b7da80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98e5137e424434917e5a1def07f0980b505a08562f4e88b6ad7fb51c9623d743656839223a0ef92bea0fa8fbd6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df9ec7df5496e679364e31f4da96b11661de402dcac9f617265d0353d6c560a12fe15285a2761731ba3b4152b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fd98c0ee9aac4a0a25a97211fd26a2e06e95c71a6da5a6ccce98b489af69594b1836199455a11e57c0d0c70b5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb377d16458be8c174975f2b79c01ad55e79c34f86784b6e6241ed8b0b5499971000fcbfa3e0b548eb8a6a33f3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1080f1e2b240af597c1a1acf7558dcc44b2e048f0d1a7ab8ed47ca34123aa58e6c035e1fb0371b18eee6761e511;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf700a7c8f2afb58166bfe458e55859800a37bbe1d92552c831fab61893be6c9e1beb9719b4bea80bb55f80943;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17bb4e36119210847a053b6a5f6be48d245161cbfaf283d0263f41752f5e28a96a4ea788161066a0da4d82a613e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h197dc713c299644ebd09039eeeb0d1c060662d5d9b0637cf22642f0439023e56fbd2e1f25e3a65ad8720725a303;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10b0681d1b7e94c511959fb40e576b76618e836c2ac0d7f85d824863ea3a26bca154416e68b56f2a6accf68e192;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc27b5d1071a7b9b2f13fdc48872dacf3cc01734e33eb0f947d65f679741033dcc32ddc80c71b6b0f865fa54572;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d90ba5d83ef34275ab5eb66f434c7fd1f2806a7071efd5b5e13592a4c16e68e9464c6644a645d14d0118ea3db8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h205610be8ee22cc52560f5a379713e39d46392e51e74e658d24296f770cab9e9ca30dcc1ff87bc52d66c47c955;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h670e3de66d51fcbaddda8eb2bc23908c06a4a1942f376976d1d236bff00e34f8630326ec3b98f97f615186219a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10ce6acbdab8a456f4e33a1de4fa4150e0f2195e9dd5a9dc764eb0df2b256a2d859e9cd4cce420bbdce1fdd12d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h136a1f06f9ee41ceb49833d0ce63294bb11104a76b04e40aa1e81cd7683c83a43a377e4fae118a60f8790ffcfb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6563fe830b2b90e23424f8952723ea2073ca723932c44eda52dddfebfa902a330ae45670cb8b3dda98bb3bc934;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8eba118c111dd3762dfe98efcbd4ab09b536678ab4ba53fbf82ed3032a10311c4387aaeccf3d58c01ceb2c2dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h180ee9eb19193b86c34a78321d51c5ba068e259d42d2229b3fc2a33b1b3f7e53272dc9fc68c1be8e07c6f960670;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce7d72d7e5e8091a6906b8084bba7c73d3040d71492e04dcac855824d799e9d2c5b1f3f1d2bedf05a9af9bd3fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcf1a7355f7f8d25fb3c93f31e4012cc569e9d7022558895ae91603805911824148a389e622ccc26cd5e9bb30d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e3566bb1a8c2ceb6fc53dee28a4342565c720c7ffb6cd6b444412247ae2c32304913137d6ce7d628cf7d8d334;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19cd56a3c54ffc73ac83cab71f134eabd316b6d8d81c27ae97302bbe19050a16187933fff3e1c3e02d096bfa1a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f749f92a2be2ffb744db9ec326052e82f82ee4ed4d524a5b34b33a34a71f3b3fadb213ec88811ce39e549ee8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b5e4c309f28062e34bdbc431343af0475aabadf423ec97cd2faf7c2e27656f5bc51859881d4abf4dc9b55b3149;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h744523e524e3d15d762654633075cacaae6cf85bce1e016135cd037368ad210e511e720c1945a4f52d03996d60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8ea323c44120af63dc0104d91ce6006388bee6be3c679500e00f9825151149632283d739ecd83ef0b10c47656;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hde00655e2fb6af5b8accfd2a4016e031f82d2c2b57293d77e8b5e2b5526b0ce06c27d57c7ae0f2ecf9ce6d6db9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a468398262e6ae3a16ab4127676b259ba1b0cd1416f923bc4b9e2af5642dd4cbe9ae91df0b947d69f046624ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d21e5008299df834a22e6a03e5da581ee11a92d327bfa58b5c281791fb3c2c6e5d915bfee176f1de56d3c3e153;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbe731ca786dd827ad3fa5261ef5197b4e42a1be607e69b3c9182b2f81fc284a3d8ed2983fc66463c6690752e6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc2cf3e10379a26dafedadfacb045c5234e3d0d6487fbb0fa605507cacfd2dcb5810e2122aa3839b5d56d31803;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he4611916548d1a4592235d76569e115e2924e8b2d0a61d18974e08ef326c3a9403dab9eb2eb765f3310ac52a44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h146d1de4f7ca80f8f9fe7f9366f306ad5336dcbf668448c8629476a476a48a7542ee7011265ca2d4e4a8f52c5a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19e3d0032d94a6b690a7e48e075ea2372de312b866a1e15ceaaf1b1c80acddc2cc3de45ddac3cd7d27c8b5aba02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4eb633a292d4a20c4d09479915f74a6378dbc36df337464e7fc0201a93adccf87905396391bb56375afd0269fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c72644e4ffa970570e67a9431a0e7dd4fbec72ae66bf0b2d64ac21b047fe82ad8be94190c9e652bc947cb912eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c45c07b7297699e80bad3f4d7f0e156ea18d370672303b574e25c0fe9f15b699d4f80362c2e50a08f8c8ccb0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h165834f176c4d0a3a6ced8a58299147b4107be64ac4fa2fca4be21fd808d975975b08365d371d6f29581d2294a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1490bb1929fd80f7f48bc7e5a18da24205eec1713467870d28a647e092f6d7a8fd7761438978168e795894f223d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12377fc3a11a0211f9b637a3dd6baf761757bd28bb08f359cb0270197f2ca5ac6b55c9bd0e362c9687ce21aa000;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd27134861e18da5272bb1aade567d53376485bc9bfb92906e7c9f7ac9d2781cbd197c66b9870c7888cf2cf12a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h487edbd2157aa88b43535124954e21aef648dd3b8c939d0f9ad62856d1254c79662b7afc7268d48a1fec2278ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16f40a93f4165467b5e7ee985a475c2fef2a8364c04cd8da2309b1f01b535c1ac8d4700630f4250a9fdc99209f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcac4f0d5a95d1066a26e44b1b7f0e88a5fcf264ed7347e076ed953cb6ae65873af4a7a6e5523f017a75a0b6e1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c5ea6fa5599708e4b868e44780c7cfa3b0153d472f4f54adb6ecca3b6c7240ddb8ac47dc4bfc74213b490a753;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h83d80a30140f4544fc7d652524a2af701a5ea30defbec682ba4e7b6cd22e0f15851cfb6d2769a16571ebb0bbf3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1da423394ef31af23f5263accd9603a535b592305ca507997d13d74981d66d0872e90d07466236c7fd46855a43f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbaa57b6ac3d5989c054fc0fa66c42eb1c6536709b6261fc32b8f4752d9578d39eefbe236eddd9039ca28c4d57f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1338db716ea6779243b1748f8f2e17a2223756f92e6acda7c086e0e2a6f4a424acba41e4312b883a112d85f8487;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1810c5fb5c9d2ea2c0b7831dbd1e584764f6f58403e10c59d3917f1178447be62748c178b97924467fc4b12c08f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ca228df6cf8d213cba5d93393d53081084bf4e46243d788b6b63681aa3c23b115dc76212cb571a04302a2b1e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h916df612bbf389f0bf28ceba7d73f8baf2f4a2c044c4664b680ab82de72e0684e776da9fceed920d2935b3d727;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h990163d8728fae641c88c83c343efcf9ec88a01c7fc76888c087504611f8e48588f20e15de7de0ea37cb67dcb8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16f0f7f06dc9147653e0c7fe54dae6f64d04bf99b2a37e70bd7de23656f5ee2cf708e1dc6608440d7ef4aade6e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12cbdcf1cb0cac6c8e007ca4bcbba51635ed907143683954355fc547a83c9618d08a61d16873698b67bd040e8b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1eeb80ea9242e3dbb6f2f132d3218c98c8ac5d7312c097dc883650516733015ab2cc15cbba88a57fa4a13f2ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a32c0365873055049aa8c11600a10d44f2243ac93f5320d0a7c196d1761afd758854c5a7e41819ae2ad99cd0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d00eb4b4fb7cfe34ca5c3c31858d4803cffb03cf3ae057d07a7b965cacb720921821512fd0f886af715a53463;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h49c87f9188c94e44c95e5ccb78a6b683c919449ecf84aba9f1e5f228d71d2eacb49d8a4e2c8bf0b08e282177e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h171ed45fd1c29b6327c3d595a90fa099e3bc01c6b2b6217182f9a87e9bb641fbf5e55274692423ca05a12c71f1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h63764f215900e5c3e3676f673662f56fcd2d92b43d850ad8bb3e0a70fbfa58d4a751668937823069c4fec1f891;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163ef78d7402e812f4380a3d3149bb8cae2636e7cbab91e9c711af6e2376f88d98bb9b7f9571440ccbed724c534;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffc3c438188bf4f85469fe589c3c44a6e588c77a0d1ea121428a28bb50064d8639770da4feba8dc8eae7391e1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c23d96aeca48c68e1be18e3bc987bd18323e8d99df3c00ffe237129a68f90d54752530ac73ac05699bdd5de39f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b02736f018b132db517e40324e363a82f02c6c9ab37feae2d9f28bf8223f3bd46c38ca011f8ca0db7900fe22b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15744dc4f80e4dc02be0a878845d9c34c0c8371d5c190a37932596a2b37de7709202be3076b328c2c6493a80143;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199b53c367251de295052f6dd2e4d0f453f1e6759dacfc440935cdeaa26b64f8582a553aa845cb3924a4f3b3164;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h301d06b3dff9685e658312aa257a01f2187417a24a2fa258f67b196b625ebad76a90df0ca3a005abed1e3a38b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12d69e1ba2d59f132cd7fddf55b0bec0cc47b0926cd80a347c50d15d756d99edb6b087635ffedfab060488b1265;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f54be92e0df6c16d95bbb0758d16159fd06929500466fdc6f0ea0f7d009c0588460b7710146c991682b8dea11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h371d23f15af7e03e8a7969668d899aa7461d0366ad507acf54d936047840a9ec59a9cb49c47255d062ff0cc597;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1469f163a94be0be316b51a4d9671a8b85ee70bfd57f9dd518decc4e9dc263965050fa96dfc497827dc007b2d99;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h24bcabbda0540110247a93626d9b8898b119583f823a65864919bed0b7e9df5aede8f4ebbf2c5895f88abc4ebd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9fa282c4358612b58f990f7894d811e69c2a829c0b07cb45c4d0aa2298b04f1b39dbcb311d5a228b1331c978bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec5f5d9840b241ff2f7e87ccbc4a7ca4fda0dc4e069f965eb1762f8d5294499552bb229c0e7597a8ace9b58298;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1849086c5634dfccc650819062450ab3a0a73dcaf22f8276e0bf45311f03b5776caa7948ec6a1d0ed964c01baa6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h27468298232b77f232352ea7c4bf38bd3dec0250e79b78a55ec75ee93779182891b1f154dd954f8818765151e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe9911f9b2558fdde638bc37db940c68248d97874e165eae066a0e0b7e5628e46c1148433c571de60b840c33cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c3a9fe9d37a807c29c566cb0d3bafb39e491581fe9f6480d15b5af3e75a574dc74c84897a994c95f22ea5832d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha8d306086072ee1236eacab592ac2b735f60da17875ce7bfcf4db836d82e37c7f3dbcd45814c097ac694dd2c22;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcecf3addc94870893a1c48956212754c5e7793a19610e9877d164013e0641ca24ad3134a842e74cae91df2ded7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d5329e683f47eac8d56471d51d9ed18d5377252c5d1fe2e4e562fbe30dab1cf723d4b55185887d5c0d5419099;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef0aeaefdf540e9cc1ac4cf83fa33dc1415ba9550c267b9dd1d367f49528a84f6fbbad9482f10856aab9985c7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c0c6e3c7b7cccbe4903931f518cf63613c5a6f12785994c73d30423be6491d04c9d10934d99d4bb49422a29ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha6eee5b2b0ab48117d5e94c89104c0cbd5b0a0b79229b23701c2455d0fc142593122e9c5dee66c192ccc7ad883;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19f6b597692bbca014f53a21439c0967fd6563e24a290a1b0e685bc8c0a1169f36757366ef7257433ee3a584470;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb763ced40df03373fa005163958d0bed6770a27dfcc287048ca873df3b41052d5a6ab0cad473f5338433ddc824;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7f8214c595a362b5c7ccf913e1252f20a4c52428c4dff96484fa61641307ca3e6da4bdab198edf992b846a9105;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a9f74e02d4176adc890212c25f7d0e011b4e870421a8eedea8247b3aa55cbe37cab9c143765b5bba863537207;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h240a007e23071a942db02d48c5cad2442e24e598e67bcb0ca78909a953ca11ad2fe88e875c306a7e7206937108;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed281d0c4059380caf341803fb9c10269a400b7367dc9ceb5c437e6e73764468ba9f2ccdad0a5ac0bbd6fe3540;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a532c671e6faf38362708d9c7bc04207a9204bf4fac2170d4a58c3fae4e0c8affbf1d46b2afcf72067e6c1a01c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8f327e81f90e2f2c8d3abb104a4402e274d0e674e839dd02a0537310846381a97a8e736ededfef5c8ae085d20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b2524035f2c9f621b70de3665c98ed7685db50894b6621aff486b183617d33723d9220d6c7ecf4a4f4d073b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf382b9128c0ea095616a300623cc4846084fc4c88e2dde637d7aff7f0578ec9d8b2035c1596efdb6e1f695f6a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c80793985251ed439cd8f9a472e4df8ec3431c7df182ab14a47f70aa17fa813baba326d6b423a52e8a37ea469b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h63ddc54079c1897c707523cc292cbedd426578da4e05c835d08496209d81b1ce9e07ba6a2f42a3ba72076eb312;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf15041fd410b5b77858e434ab82902b68d0af851aa8155c746747e1c69113b5eb4092f98a4d24ca5bfcf8559d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bd8a79b915029b209e586c134f048228e555250359e4f93173cf31f6dbeeaa0f6b4a2795464b96ebaee38fb6cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc57c08be352dff713ca8baa2cf89780b1e0b4aeb4b1d98a4ec51e3fcf9b862ca4cfbf30a56da7de7a4bb66cd1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cba2d4c24f00d4acf4eec93c8c908ca2a7ef16e81799fbeb7c3e90bfd06a4462a62d0ffa43216b863f1adea925;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b96484aa6235671490425cfecbc439eeb2ac878ce44762bfdaeeaa77857c0d939f27b100ed239513a022f9194;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4e10410476e093f70280abe585d69c35a291a97c0bb3eabc525eff97f227799dd14b89ff01c76a302f6fb3f1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4d4d4129c4e0ea8208a47ea3ac0f388254910fcc3f3db54d2e9dcaf98377be8f4763a333c417a0c3a4f55cde00;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e11216ba9834070fdbec82eb3f2618950562a843390d7e96922d51ee208420497c9768dbd3ea0285b650c7fa2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195faaea6344996d4a37fef417aaa8c180de4458c2de617545b66201f65022437c40ede2887b7642ffb0d54294e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a18849848cc6e9ef949c33706ea4efd3096f75c33c144197de2aa733afc3e90a94a572f903323cb3bd1dc1b7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f4328dff7b85d160ecb3ba22a3580e586aed2c2c0a19dc2096ef9dd6df7c4bdbe7fda4ba748e53cc65586f761;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159e08e6cc2a4831c11f6e32c847e6872e439e2844747eb82f729fcc4ff0838d9c1eb57f73d2513f76692a7193b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156f17ff0e27b45ec6cbedc3f246282592527bc48a8d230a430b1f252917a7acaf5f6bd2a448a5c5d3d24d0a05f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf39b6b3cc7dfc625b527f77d96c878641471d0603ab2db31046768014a08255e7c15bcb035c8c93022865cfcb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h27c49d516afe4724aa4110a713816bec188f66c1007fb67cc3a243ce07d6e21829c9257184386728328ce13af0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42a9ae044ff778826321b8b39b7b325af65c1fd7831af31bb56ae22f72244ac5136933acb2718f75a4f4905f67;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he9e92ddc646a3a9b1f045ab77ec7c0b9d02cb5fb3c249d0215ffa91322d175da90a1b5a80549af0406d0f033ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h187511f9c316c2e8e2f0253e9c44d358bb1a08cd4ce33501ba4027d2162fd44cd4b105f9f7e6b0457bdadd01cc8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6810f249cb5c5019440183a2a2fd3cdbe8d0dd468ee7a9a8c42e546bd4f4374cb1819d415ea6a4db46dd7c1f7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29e61dfe0f6bf0d1d716a9aafa9574d5c1fc6cb9532dbeee8ace569aef3c4d1d0c837f1014fd1dca59c985d144;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cfca064432ac84a653962d31a156a43645e15d1be39154a496118ab8414f699232b3b0db817dbd7d0efb81e732;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hec13429a49322e7399f3be723a72e26ea2e1883c4b3c915273df461da89bbb62b296f064eb638c9dcef673bf5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he45d6dd93b8611d01a767199c37a7dba7a7762b66b7daa531ea7b36affae3c26be8f85d4ceb7727ab3fddaca6b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be4bd6f4f7f3c021b575fc82f85e7ae22627b2873185eb2ec66dc46422cd7887395c66b1f92650204660707613;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d5bd47972dcdb8d76e2069c3062de5eb30e0696bf870e22b3ff4210c8ec1acb1afafa29fb350619dadd1ce5d98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca3dc989f3c0ad87cbe76f3db60bf171315151a09d46dabc58fd80ae1332c9518a852bd9f51950c4f7a3db7643;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193483ce35e09263dd5be80859f53a902c995aa4cb230955ebed05ee423c65d536cce8359469b360c7bd33dda9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13fd00ae531085b693c60f305b1ebf60e764eb50b6687235ed1366d6686d4c34bfa7688f94ffc672d561b861ce9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10631c1d5a88e9039e86941511ada06e590473e50fd45580ea758d55e03c91f159e868a227527c49ba5da588d39;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h148c46529fa4fac6e99f1c169a0d8cbcf601ebd28ef4b215001297376f531e8e70a418f3b0a6895f1350eb9657e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d791cc570a36afcbb84be8b24e817b719a8e757721b706a9e4538106eef39a8bf55f14762f3fe8e1cd484f7d8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d8b04ec984843b1b0751c0f8c7c40444636ca2879a4c2066b5db6766c49026b7341ac1c4e063d418474a65772;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d10299b983605fdf6cdcb60618c3f77fdf1870f7f2014a89e3731e78aeb409b175f3839d02e1825b0c8f4447f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he2da5d10c8e4141ae541f33d04ed7e71803513f0d48ffa9507d4832fcbb3137ac9ef17777766a13b377b176a32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hca9cbdb9376e8875f061d34380aee2b4ef96ac204e777412c7cec783b92123e7fea16de4bde4259efe3abea75c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f0a4c9a41a37760224682a418dbf1407543de1c41b9056d32f8d871b8e3d928c12ce76a68f253f077e69875bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19144bfaad8fd5c9869ad56efb290899f9087e7fa4ae2886cbe0c59074a7653f645c851f5cbe33922f8850e534d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0a5bb67f4db87cd6ef4896fbbbf13a1c08a2a795a677c59bd0fbf688a05e9f3aee1c62b6d3fe27b76ba2b8e83;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe33a3e9d3bf175b94da57b4abcfcd7635b9d934154091cbeb4694994b2ee98bfa65232e97a5ac57c6a2827b82;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1677fcfd8dbfd5c736396fb6d6d3e924d4a9e15f854398957e24154f83d24b7ac84a51b8c7b9e15aa2dca4d2dc2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a26928882be3dec98f45504c24cc616d1abc4c6197193b63a65a473dd76f5a4aeae055a341d58cac19ba1bd24;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h699b4c6f877f4f20118b8cf3064874ec42b8b5b79a91c657d26c19a3f95b83c86b2832850506153d1ad40455fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ef09f781eb0ee3c39bc23bc53b9d008688a8e5faf523389378a377405c0bd3219da225e58dcd2ab80f784e8a63;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1976e43991181dcba01ba29b93e8f76ca343707a036dd72a2f261c84f3eecd579f68dd508cecd0fcfc040deebe9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db3ff82e6f64b4afc0d79bff2be9eaa8f40e4a66751f1d40e64cbf2d554d2f528c73ffb4663e3b6e3cb604ed71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8aa127ff0a7446ef1f36f0695144d27661fd1bcb9688c124452e79916d4351bc259b8bee4b1e1247b7aad5a2e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12ba14d1c6c8b3f0272d45ea35ac6a37f44a7c69612cc57efc8fda070be00bfb253bc41ccb0a591986661ff7898;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28dca91a4c84165f132ee780a81418cb3e0e6e1800fdbbca9f6e465fbcba2e543f07fdd234eb390c652f28942a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h120b9407b4dd2d2904595b4d6215f65be77566510d8407b4d8ac7b1f7911e1cfdddbca145941638aa17c11456eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12da311d31dc7e73a272eb08d1809f39c7a472202373976115154d05081e92de6f7019bbc1247c55ca4b221310;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfce322d7a4444ea907339490166ce08efa9d5dc9d1e10589eacd842606b11244e7be6c020dddc56559a2d92413;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec630461d25d8b20ba0d6dc30fbcb55e9661bcb70e1b7d7c55e63c8490e694e6ef705dbf4cc72abd85da54ebff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14981ed8141e0e803ea8c63affeecde2f4f5364113c696a87e0b2119c4ed1c34b58050fb86da0e7fb84e90d7a21;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4032a52c8b8663915ada36089e0b74fd068b849dcdddff666277912a3b3f48bcb6e52d7d670987c40d09cbdd44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b546d2d775b183c725d65113883a8aae2f358338a06517f17888f5450623de54934edbe8138d8c8bf6e2ed014;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a8d6eae4f2e4eb468435053e11676d58c347bc434adf2951ba9b06257f56cabda80b0cecc46c5eb534f500460;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0420a9fc8642a5747fb44e53140b39561356e6c81e4e7b8455671e0d9c81073b929f49d1e61fcd7392fbcc822;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h921fc2ebdee58b14c3f86d433e4469c5e50307c92d8484200883c1056a8b7a0a06e5213d64998a89718039506a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13feb36da5e7e43f881c631a39b75ac73f8c1af283507f86329a5bcd26ae75686985538b57dc6c72f53df9f56b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d5546af9459a1f19ff276fcb4f1870a8c16d95902be71a08da0e9732442233c6b0fb541c569b7a8c03c6741e06;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf7e0ea2c62742848263d3e0f0669cc770efd712bad37da7280f71ec591d7947f9aa0dac47c77c1cc14849da48;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdb8f27fd7190cdd51adcc379c48645b8d1bcf155dc2b2abffeadf1d9da0ed81b9c4844e0e90c0e242fde92ebb7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f073f15ae5cb031ea1a3dfd4793e88610c89afe28910910a5cb92c7bcf038aff9aaa2b546895bfe5520d66dac4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h95702ceaf95b91e89391a002597fd17637a3a4127fb41a82dc5e3e445f4a722fdfd05075638daa78ff222805b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0727ccf2dc29919d43bb06c8d32afd64bdce2d0679f627005d64ba3aba348d2b4f0ba261d57538efa78fceb5d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33ab764c652a8c1f85e9e8e3fccae18367932f5a03007af2e57474b544b3dc60fbd0005e973747362148b93584;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8c548af26314e2a77af0f24e17d17d1865e278bbef072ee3340a9fa3fc23f66cfbf5dca35865190043da2b682;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c932f4982acd7d78b4b8c97306d8f69e489bc6dd824f99446e67e23a0b5647194e4e89577b41be4226237aca9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1abe9193e763c915ca7ab93aa90e38ff22d04fa89998af787f70351285422a6230bbf4c61a6a7c7bb6f1e73d5eb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h123d54fe32d212c234a25bb8ff2b6c441cbc5b4418dbb1d967bc424902e1f704699fe6997d37642f8382cdaf092;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h799face5ae19256bd7bc4c525d7caefcd0295ccc4de4d60c0123032745979942f32b5d35c88f2dd1445014b7c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12152810f181f05112216b677bfdc1ca702cc0e504895c6425c69717ffc3b7b7b357fed2b8f8dfac8fe942e891e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a0010cdcad5b059b2423abbc604f9c0acdbf9497d55e512b56b128bce6c9cf60af7c3a4e5bb3dbae19e7cfe52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ef5d35826ca0822db8f6d1995360f075560a393cb4cc03bc6945c5896d6a2d190a6bc2f5701e79e168fa96d21e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4db6d77e308d92663843330b001556fa95f5bed627cf85ace0fa8a737ce557833d989874b6b705f52118471f80;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6dc8e2afb148a1a5bfdb122067183381d4bc2dc2423002d88400a4cbb7a9648debea0a436f9f3cc8ae3b61909d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7bf78b49facdbb1ac5ee7480a75999632214ed558ee90ea1450fce2af2551ead39c2c5a2cf9f755beffaf9172f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9bd627f018bb9fae9aa746ef2289d5b73426d640d8227ec4b969b298c528ec45965cdc28e843eaa2f2f3ee1ed8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9075bd0c05aa820827ffa55826b76780ac93f13e659b9e9bb049f49186a614388dd38bd4cb729f28b47d961084;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b3b4b0c61228fa27bf5dac6560d8a837466eec4da02fc6789bb7d7055c71201b55729cb43ab7b723a6a62fb87e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41c72a9e9504fd7000ae096dadbaace19e11ef8144a8d6b2ca6574d92713e50bb6fa2c826461575685abe46284;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd35760f680d930ea394d5faa6ec1a4be34b48c833c723dac4e22f770c0350aa8f22a5efe82bc3180d2c608a6a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1295d0461179a7256bc2064ec0105434eb9724cfeeb3a9eb3abb6dd230540780e3ddeee898131e056cbc1644fea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c1f129abb3c59dd1d7713c40fb604dc86d678e13bf88d803902485daf1b57687b85cf2336f95553e106c6aab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13008aebc4b6f03b978360b1fbda10ccf664b0b0baba9159bf52dfebfa2bcf9e8eb7fe5a6fef5606dcaeb313426;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0c0dd088d178fad05c858f24c3c2bc781c7af892f5660409a9726a887fee6f5d9dff7d3d9a266e89996dad3e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15baed84e240f0287f4d663bf738d30b7e37729fc2599a5561b7383c94666ca23c79cb0660c4bc756a6a34b4519;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41b7a338eba3fb6599806c3de47a914af2fc58ff57b1651f42e5106445c5c0fe1a8803eff2f247fc3060c87756;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h62867c3dca9a2ca01d57be1ebfc6cfbed3b516e12b7d3f4b0e2f03fc09d3fd5e28ff0a0283d3f88ee6696f4f73;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c59645e72c71f9275b1816d14663da138f3402d91680e41f01246ba00d0b18701872c22e0a28c4d7ee30eec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d6c27c3459de31042c411ba1aaa020c0d5629701e7e89a38bd3fd8340996b1ec2b20ec693bb79a5800fdeaaa0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a99a0af8949397c18ee318c2be2248b5ac9d7f4c228eb06bd0fc994c2c8e0659570e039f544018bb1dbbd2ac0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1726be1c30991775f1cdcbd569fd4e1240c6e16e87d19f1962b849d8110d9cec6ab06271c51ec0b430a42c53028;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c81039a95f2b344281c38a3206a891eb4da3a6928d33d92f4434733dd31894d29b970d6afa13d236720412059;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f93db836d365dbb352fbf4a08153c182fc62f2de78419d451596c1435a123c40fd14f8362b0c107277150309b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha60fce5255cb6683ce99db544b2ed6aea982450c6663c73e26cc1ccf59e1c350bb871a796ffe402c8e75f70b07;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11b656164e32654fd9bdc3cdab98781a844b02d10e3bdd9043aae51e0c0d5941caff2062db9180d0bb00077c63a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda2956a53ecaa3576b812dde0ca5baaf74f99e24a1b6443bbed2c29d90ca7beba23c8e82ef90616a2d9366cd3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc512e76301d02fac9ccc6261645392797d36f07b09f4e7f91dd5d39c0a19b057f872f7c60ef6e54e9d4104f95;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d3a5fc75eb1855ba605c123c89b394415d22c5b1c031266e84d9eac2be049f6dd2320beb2e94cf5a38db4d18a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114d31491e193ca20ec8ca75144491a25abc16a0f4af743f8ce5f1f9392607cbfcfb053f07ed9af64abc87d3767;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he37f645dc1011804b65d6a6b5e44f5a318cf65eee7a5fd9b72de75d84553d4c9f94b3ad7f612e4cb6e64cac551;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8b8659e1d5def49bff45d5c5b57b7d7fd5d26e1e3134c957aac59f01e46ceb602e2d462832f14fe0256acca9c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12f13822f63b42e568ba6844d4a57b885bdd612d7a53ab2e61e5c3c15f4084459ba10ddcdec6fed418f90bf4a9b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b6da8441679f929936d997c6c226dae21baf976cfac0b9de6c610e449882b14b31d1fc41cb578096501ed2853;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd42558836418943d88b2ea5da71115b062ab30bb9c1cd38a80ade91d74f27d8908b56f32f5fde9520d672296f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e2d69a5fea2e3486892490b9b8f9f79fa40ac38e704394a57cede87cea16930570c44dcb016844052340f31828;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8095f55d06122093a8adf31a36439c2dd8bbd427d0dbbccbb2217ea07ef508ea5bf9eac03433896e98ce8750a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he66a3c135c545d624c7d251a29d29252cca6680cd1aec16347621e6faafb1720a38fc45217ec945f2f51aa8f19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e80c45cd0ff6a03ca8a3b6783c80de909b5dd6bcdb5f4a26f1f5883241ce4793e45c068181b3e086ab531821e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5018ac9a9f3d336b66011e15bc30d1fa207a1ad147973ce3469d9c8822e6e91b17ce7f9be0828d78008cd5fec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19f0093a77f440f337ec9654488d41a25dcc0873daa563117d2c64dc1abc2b471c29a38e2dc5dc2254c05c0f87e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189397c3dc480056e162f3a9dbd7143d95f31e0ade721560716cd4564abc4d3f1a1798538fa8a00c50081f9cf43;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c277d38cbe6e1b8832994a30afd4ea68ab6b4209a45265baee70c76317af1c02af0eb3998bfcd596e8c616bd14;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d3fffdbf6e571e13304f375b26cf572cfc7b2bc40693c64a572b27422d8ae1fc7df472a97b03f0f9868edb752;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a79b8d50f40418e807f46798fa092a32cbea195c6f154366b1d59f1daa2fb2f6dc985f6957a8890af77bfb7cb0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16953965ce58b45eaf3d5f5d07517d8c98b80ae4c06e348fb9efaab960112b8987d211408b258f579fc80980731;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h124c77d752c03a79c86f9635035f93c329edad83fdc2a16688470e2014e7d1072fb0038f37a6b77ae275e5665c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19f389768a123c2792fd47388da911c4b072f404d26e7ebda1aefa06e89c325aacd45a9161c28969b6697a8e768;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1739efac67b33e065a4261b28eded121e3aef9e40cdb86e69c9b1f32c9261d4199c762dbc1f9b8c79a793c6f114;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a4f9f33ea46ab9849be7cd8f3e07c9afcb41736ce946bad4ef4465190b65c12e07f8055c0f9820c5a31eeccb1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed892471e1df4999719a9c246b27d5cf45b89a918bf576bac152364bcdbf5e859157e11a0482ad5cb731e057b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12413b8a935a9d0bc776bcfe4e239c86ab567348f6c9d6d3ec7fb62ddb202dfe37e2cd7e995ab0f65ab81c745bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17617b7c9bd6e632f8e95fa50c0823fd6e928cb48d24383be9d6fff1cc5ef11148af57cae566a7d7a81c49e9ac4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1599dd33922ea05dc8eb8da8a5f2ef7d4ee6ac6edde61ad09ef5e3c2f301ee54089046fc3b5952a8a04e60bda99;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c7e106d5cfcbdd939b09ac091bfd5847b34bf833754fa416c42ac4acafae4d390ba636e50240fe79833e3b347f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hebc807e1368fc2dcf30c08b809eb9d2265e8a589349d32c3776ff4920b23a3ceef6a14e4a9e50c76ea131a8129;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17055c4f8c8dc9c0286680434c895072d66dcee24f4ae1798b572d9aee2768f5c16fe77e81a8be13aaf10fc9fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4f753dbd7dea76881c324bf43c0877ea1314e40ea2a57db5d833171b58b1962a8e9b9391574708fc2d9cf8a8ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bc72eb42c7faa9f0baa43dcafce513a02364411375ecc3b0efb9087fe9a624b394d47ca5e850056182d730c52a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70f0a8bfbff5a27dcfa471cfa6d36486266fcaa7744ab6ccaff1731864fcb2a266db9b8eab0ee1dd4cdd55dd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb40fe755dc9b308e90381ee684d4e3499d527e177b162a6208ed07020040d95f16493859e575fe8ff578a85f5c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he62802b5472bf5d78468ed9f5a1c659db2ef5d9ea18030caaf42eae92f727e62976456f7fe6449db022dc2d5db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h63f70f9d0f92e94c5403bf6eee9c36f6cd038953332b94490b45b3adfadfdd1676659a4804d4bdb8d3aeec7082;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dc2a207a60dbfd9fe10937bbc118fe9bfd3db83e95ac0e81ee69f558531a0b75133bfa7265e073c55805c1a413;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0f76086dcde0bb31dc98dd187ff10feef31db41c47884c8cbf9155283a297b2477e848e4c7a87a4fa894ccfdd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf338076a7006149c572a16369627e6924c1ddd3805f1882eaa53c3fa53c9028dbc684ca240072c4f94f31cec7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16db3e3d5775eff02408787fb310359bc5d3d268e2e107da54eaa459db73af30f78f0d441f9f6c95ae5d46cc5b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9449958728ccc5a437c8aebb9c21a75205262c980ff289354e4a1a12764171e9aa3469ee5e056862a28a6dc66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1838317448a9a103a512764f786101dbe8ed72e996de5c8f74111a1ba44d4eb09c534f52656f91fc3c33151b481;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bd1e604cc4ae57ff2267d5337b6c40c54e02425d5a7a7be7dd72243223c55c9bf99e1ef7d9947fef4e93260024;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h64d7065c10d06c6540f51ba6b078e2b6eabe40f72ff1f84dbfe653ace89190e5212f2c7a84ad49a846af3e708b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca44608a5e8d55a722259cbf886cf654c5b1da15b8ea0d1329402c3216e1a38429afcf35e1499da9629c355c5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116170d9f76cf8c95b4ad0de92d1c6e51823aad31e4100bdd850de8fd4a1e02ed75929c405ceff44099e8b47416;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he7a6c3d78acd5208605808d9f94ca34b5ee5cae97822327de44c2663289c5e481c8c9a1fb9afe00cf1ff89823d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1991667a2a169ce77617819d4682e6f346441bf63bc257f4be78c5ba48983533d1bb3bf69888d8c711892172d95;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c73526a87b85c07b43457a8b5022e370b971f5177af59de25c17d30877648e731d390189be967cc45350c9c1b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h144f9de5dcc48eb9474d4e39d5bb90f3f35e600d6c914beb57ab66729dcf66b691bc853548a1789cfefcf8e0dc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fd7395a2ea4a87b3496e709f6fadd85787e542e95e9355ee4398311ba83c0c3de0d84c47abe02e98036f231eb7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed7888c11ac2063e5c56fb6e00f536d6d560cfbbb9c514ca2b13ff99f623d6690fbec46774d42c9a041e6aaaa3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dc6e83a9a24cde494b49633367ca78bd1e2a22aa9ba110c165c7514c056dfe20d136dd437642d45a0f3f2a0415;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9dfe1733513a9711857f4cda7043e54c7ab686d3463793aa87fe0add804a099cbd5da2f7819f1b48918b2d87b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19bb2a94e26e5113095de7c131c304cea68c4b62b6fec6c026d89507918286052b0ff9901d5b5ba14008ae26ddb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce8c2553374b7ecdbf9765abac61dcbbbc4a65d0b8b1da1f9844a3f112aa1f616fb475fc27ebb6c4bb1cccdccc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b1e5224dd8877f34199113e43b8b72a27a1acf47b459ec22bb39c8c7f9e323899e911755d97b123c0750ac4e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h102ff3f6f0a86d4aae445830ce6883402f36993a7f04fa1429d044876f18d391747d42b60301cf0ef775ef3c631;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ffaa2fed3861683d84da90dde962ab765caa689f8720fb901b80b9a1bd2cc8e90904819826e1b673e1584bdca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d6eb0c0021d3a6c7c1e16376255782c6b37e29a21cafaa68d6e4e487ad005747b5fbdd8845f4f5ce633ac0341;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h187a9af8eb9fafeb4f80ace7f0594ac17dcad999d8ddb964fa347ad85054ecb0a0abb1ce0aa3f4715858213bb60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16fd92a9a942ab77f977e89666fd740aab21a4c38953fd4720433961b3d9c52dd54fe0c3168cb81a185c2d2d3b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b82ce6830ea712f2f8180d6be93ac6dd78888da363de1e89c956faf7ad7ee6ba43b910f2b5202c47bef8bc560;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107976c61658ae22c50ee887e6c8887495cc8fdfc598ad32386556baa30e9c13c2e3592d30a421b7795bafdc857;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he283cac20836706f92822649889d9ea7dad547e7f119c68d784b691996dafb7e505e27ad7f6a8c01219c49dbd2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ddcfac236c6427aa255361bd44caf22cd9b724dcf19bf333bb3528a70c616c31ed4777afc85c2f1635b66445e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150532b6434f7e3fa7502ed94721e9975f6a0329f8cf16313af028668c738d2bcdae76697c39e94634793bad319;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba59dee66149622c6a87cbf2842570f56ea351aca95f66c3f93d70cfb9cd87154e6801fc0feaf208b6758983ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25ab2e0d80d8b8f7fb87b51018bc8dc18c94475e28dcf966fb35c8d4b8bcc18a770a663633cb76e6330e3982d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ebb64555661aaf160373ef3d54ad36133b522353ef58dd2331f3fda78ee81912420c2700e465a110f5f7e3b6c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1acecc56d4388b56c14431cf64dd08caaabb3d777554a9f3bc0fdd6c024c3af9bdc78ac2c7032277ba4f6b6aad8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12ec604db5bca4e32ccd0b29e959c139b4d93450d070c727b1c5e5d2936b29437438a3796740ac84a0d9d1da57;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14fde904631e44f4353dd358517e4f2e8955ac842a8b485506ba73995c0888249c1dec019c0a0304e26cc509b8a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h830b24f5acdb3a75897c88c1e8c4822e1fb202a35bb989db066bd23c714568d59d7b7fca9a323620b27245c1b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f7fd446ae82a524fb6cfa0469c683769efff05bd2e7e651f9c5423fe5f58761f37d8c4a3cc3d62dc8afe9aed4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ba8ae2634411f7e78c254287a2cce315d9cd5d98e2d43333255129ca01a89655bd1568a3338dd8470c96be48e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h789a424f3cda007a854f5556ac0e9c4c2988ca686a3fcd98f401e9f1ef8cc1f0dd4f16b97ae9c4be9171ec688d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cffec4623803395de968dd410a32e2b594f113113cd80d7a500ef03c1d9f5b38d8b3e9b0512bcf30291418f7d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf3ff6747073ccfe126c89357a55deb850abf84b1cfb31fcfdb529350f945f207f26c9a74ecc620240e965f1b0c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h79b95167ed5bbaa1c974a873da3b082740e06c2c52e4ab1fe8a994c042a6c149cb0cb23a48a8bc468c5a2d7f98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa90af9ecf31c8195408ed2609508838df9b7b7b8ccb36ca7a6f3caddd9d1cc84ca8ab70b4ee65e4a0f2033bc3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5bbd0f9ce1e83e6b191f27d6725f9c3fe78858a649038294ede2738bc4406a1c2a12449dfb71c94841fb3e81fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1502ab309d20462749cc9b7291afadd1096a1868c6b36a87753ecdff323ecf232d9f1dd659976970ecffab88507;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be8076dcaf90270079cf180daadba1ae7aa72cd153b5c3ac65ecbe265611988bb347ba6d420b63a7586bb9c3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1112370a980a1f6f892fd848a141f19bacb165f121efe1572439fa628e168643fa9f804c20b2409f3dc7c7d907e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc7b2e9148cb683b2a0fbef11bb794309a440f3df08f67dd3c3def7670ab1eb10b57f8fdc6a68053634dc1b18ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c5c921939b3acc75d8fedf047b7e7eb7beac0d106e20ad90e74c9370f56dba041a878d63e5a05d84a396baecee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h776fb3c65b6400e75ab376353369b1cb1866a16e4d1595cf5d23226b6c7a292cf486c5ee8d03cb68995e51aded;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1104bda5d838dd4c5909e1399c2708d584138bfc5aef27e8974837b4f2792370add1b8fe2dd83b8afe080237b46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0ee4288f11bf7336ecea381300831fdbaa68065f3d1f880916e02201547c7c8ae0cda0becc18c6fc73251d090;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8430c3ffcd0eb9b86d273b39f17f9c622237af7b92bbadc229e6da6852a4ea237f5bf2d686498d2e81301e8006;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11b8600ee891e663cc5017b24a31c81ee53da50f2ff2b90c3f720ead766a8381ebdcac7ed8a3214d641049a2096;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb813782954a4c05cfb5a756c53c2764b1d250153aaffd03190b1b332bd8140a441bee25bc9c24b13e0e9397b3a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fcad035a66d13cb25c331767d9292984701d0826c66a83b2b74c13791aa06e39a8b61560ab81bd4c5e15d5e85d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hecbccccdd14464bf2216a1598f9de83e3e2414d6cbd641b1b49ee16e23dfbcdb648511f1feb84389980cae5409;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12691549da80f44646486a687308507a4b746bb24336689c0124a213b81c2a4b0b6d5660c17f4b8ba967dc1869e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h850bf23cac266b6201e049f3e2c781edb4c43bcba439937d147d4ff980bf13854c543084110b06ff287eb92432;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bdaf0d359261a5ffe37f07d54f2cf8bc945e984f529cf72e49e3cf831d520ba536e1c2a5c3c803cc0386b66d6a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b91eddeaf3fd45bcb518e66b2c45bd352bb7de2c2c42f4b56f9bea2097eb0ad4c123c1c8f1dd5108135921845;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e2b1993ac4b84b748884fbfaef1409e481b03df7763e2c65760bf18d5e32e9d30ed62526fcd2bf6deb90f1f5d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdeed1bc6e906acde471228e133cdb17b23af514c052cbd10a68a0b9b18971b6586a0b9ffcb3cb0b46b82d1c8a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172cd79dfeb75960997c21df466b6cf23944739127fdf2b8abaaca42e7e1b441fc11206a49a945049740edd2132;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e786be0b86ea3378a11078a9eb3246874e0a1505e9d4661fac50f9e92d83e4f5bfd21d8afd30d35929daff5aec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1778915ea3af4a6692701307dd872edf9cb2d04bce310cb249ec9e4e8c245d9181ee4ac8f5cf2b69eeffa535867;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hefc3945f6b874f94e6e6153ad0d4ece5018820ca43556b2e01368ebe3c7aa00082612d347a7eefb80adefcf36e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195064742cedd04e038b99b8e80ad50985a20dd9857e42b1362d6c17ee9647b6787f9c270688ed8dc6d5c36ec11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b9d03efc6f5c9c751f59f4cb71aaa87f4e80c53deb8f38ce1c9249fef9b35c2aaa7ef8f0af77028a06288b034;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ea1b9383a21538bcb05069f4fcf6b439a367241ac857cec1632206c738010930760f2bbe0ded94661c3d51fca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha1b9103eefb32d617ce57389e6090563325753b60f2a060dfa15262f445dd537eafa64f8ae11125686173fc819;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h123ae09d035158724f1be34aba31c2c12c9125226c2f77a088a4948fdaeb8db76a68ac93f40ddabe0b16f3371be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2505171916aee7d4a1a5436095aa9971a49aa3dfc9807ec167b3d6842a936b854e40c01c8b63fabe641bf2b695;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb0f1d8f36f91b300c0611bf875fd722a66765dc3f4c29f6af14527a3b341c1e01331730fa3f50ffb103a380c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b52ac2009a2136545deb9b480f19a5cfa52dadaf17a70a5102eeb7e91555d7b7b7bb8a42f7cdb9e67b85db23d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3396b7687b0654c7186d1d34c70fba5115009caf099483e1d9cd927265fa3da8e7379d1aa70ff0ce86f42193db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e66aa8c7768464a70e1e1c92aee8d410bffb5cf9a25f8a1bb5fe0efa5839f7fbcc5bb79227ce6a79de224b7e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df58b25961f343947ed8f0df402158ad5375570e7e9b753e532741dc5b4ff1691c8e687dc3a84c17101491aadf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c6e24011deab22341aaef7e707c9c01eeeb580be68253067b163c642f7ad442ae4edb02a459b857f2542d4904;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33418a0ab260a505794d7072b71eed8507d282c4d2f6a5b77d376943b98968a030d6f4c0f6afa88bfe294fb3da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h48be546b2c13dd7129bdd178217b111e742889eafb461bab935f52cacf7adf0228d60e5592da590045045cd2c5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17196583a490fc488f144177856b8594c09c17e9e2bce3d2294d9ee759f724a7e5f63d28b17408b59d682179b1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128cac25d9ad2d036398a9c6828f4d4fdbe8a6df6cd1b46245e36ae03741e578595dcf68302de9f84c9e50c0345;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d3cae935b135c18f422b9582284ce342b49a1b0803eb66145f7d4a2a013a018c22a5142e00875ec15eaaf064c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad033c724474f2c82573654897443446310da691646fc935974482e43b006bdcb4e6aec828f256e45b3114a5c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1574376418206fb7c0e5688c86204ff4f2c736927f2250ef47d09264b25b27948659ec955ce889f3a21e2ffb0b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7bbdac8104eb623b378ecbf455d5abfba754af614bb19fdc1fb194d55c216b985866c28ce0f29106cd778d8078;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b083b0610cedc9eba97962a122c53bfb9d172fb37d1299f51c4c8dec651dee4c413c93c27a9a32f7d8720ed6ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h721505949eee730d2fcb6e439000832b2ff744f9c435af8a0d185d366535e401e7298d1a0376dcda86987a093e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c57677237dd9b636dd1752adfc062c19e00404549103ab876f203eb914d5a0c827a1c469a9cd5886a0e9d2b4b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdebc10fc12771a9020559de723c59365c30aeb10fcdf818f0a46b06418b414eb0db9cea317c170361170998c03;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h65c492955f393ec068e059bdb8a81587adc49876ee893d0cd3ba6007db4bbf9c3dbc07533cf2d1418adc0a1e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h111d344b85c8d2536f96f208c6597713d300f600bf3ad687d8cbd1bf462751dbab5246ffe8422df4a279bb42c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159ab094ee7040c9bb2f5e4fae91697893421dd0a1853a73927c98ffbd9eb38214a737b01f524bb542566c5173d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he04f2e303b6a96733f7f38d20c88907f65d34d23aa221a0eefa7d0a85e554c0b2246ec5edc75d0f918dad1b85a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8bba5adae3d59c83f66619b917de865755cd4fd29225f4f03e8c4494b5aad9d56014f0fdacde9d62fadb00ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9562dc7e7593521d1a75b8c4d1c5a77eb589aee2f9fd50bb01b6c64daa1f09eab31fb952820af23db24234128c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d797ad7843c0d86807f0468a62d93442bb96774946e28679d1becfe7ea6d474d7e9a31826153fa96a6f56c71f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132c604ff935c99f134d0706f78aebb773af159c2c02bb7fd9f828b1df5f0ac4e0ccb1655fac065be6cce270fe9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h43973551adfced3ec2ff30cd871c10f223056f7355076feda4c8a312da813fb84a40e00051ebc6d40032f85dcd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142f8f29e48a73a2ee19550fa5721520d72c7eaa77ee3f4ec38cdde29f4d3c770dd13f85cef92d26d1290d456ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6749e37806ee429da83776582228885d7b49bc17a34c2e4c46a18f046e50bda898a9417c765d9e843e51306fbf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb6e5ae49ed65e6e276de913f577930176c6c53948625cb66a0de1f1505420a6a77c15758ec3c815d7fab965c1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7d645709c6d7022be5017fd0573870b63db968f7cbef38ebb748b887d0a4631bc9c6ae538525061e059a1bb7a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h30c42ba8e1d68f067e5e0ca3972e58d722cdda8334342a276a05034de377f657a9c74df7e5a2c0b4168f8347fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h69706e38f68600e13322efc77583ace51b057447a920d3db59a2b7179406e33f002c8a43d4c19c831ed761a78;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15513a98d051ff7ef0c5c12a6ee2882b30554c1ba4868456010019b122d635283297071ee0451950b0e4712d0f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd30dc390db59b0008a5a2df7733a09c951290179ad0201ef6fe0b77da2fcbbee6c3328609b12c90a86eaf1e3fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h747f0b1fc603ddc0b3a46a215fb209c907c233d9d018e54ebd9be6902cd6ec124f8fe58eb0e4cccb3f89ebed82;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb0a4fd69f2274e590f531230609a3d88065f08a738357ec4bd6917c00ed0058710f9e453ff4892e8578b2be53;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a587a0c2dd5c41ba15498d3178aa06d2d2850fade35f5991e12930ea789ac6d10bc429e4abafae87125f87420;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1562ae33d219f0491e8531793dbe98eb0fe4f85a379de6e7fa749ed279293c7e2f6822d0b64168ee0b5a742e057;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h123583174b095a188c2cf14b911ea91e7015aad05bca1b7b2739a8c38bc5e98efd6daca8b19dd6f0f61bc804511;
        #1
        $finish();
    end
endmodule
