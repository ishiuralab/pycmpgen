// probclass: mul
// size:      9
// stage:     9
// cost:      10
// elapsed:   3.2576327323913574
module compressor (
      input wire [0:0] src0,
      input wire [1:0] src1,
      input wire [2:0] src2,
      input wire [3:0] src3,
      input wire [4:0] src4,
      input wire [5:0] src5,
      input wire [6:0] src6,
      input wire [7:0] src7,
      input wire [8:0] src8,
      input wire [7:0] src9,
      input wire [6:0] src10,
      input wire [5:0] src11,
      input wire [4:0] src12,
      input wire [3:0] src13,
      input wire [2:0] src14,
      input wire [1:0] src15,
      input wire [0:0] src16,
      output wire [0:0] dst0,
      output wire [0:0] dst1,
      output wire [0:0] dst2,
      output wire [0:0] dst3,
      output wire [0:0] dst4,
      output wire [0:0] dst5,
      output wire [0:0] dst6,
      output wire [0:0] dst7,
      output wire [0:0] dst8,
      output wire [0:0] dst9,
      output wire [0:0] dst10,
      output wire [0:0] dst11,
      output wire [0:0] dst12,
      output wire [0:0] dst13,
      output wire [0:0] dst14,
      output wire [0:0] dst15,
      output wire [0:0] dst16,
      output wire [0:0] dst17);

   wire [0:0] stage0_0;
   wire [1:0] stage0_1;
   wire [2:0] stage0_2;
   wire [3:0] stage0_3;
   wire [4:0] stage0_4;
   wire [5:0] stage0_5;
   wire [6:0] stage0_6;
   wire [7:0] stage0_7;
   wire [8:0] stage0_8;
   wire [7:0] stage0_9;
   wire [6:0] stage0_10;
   wire [5:0] stage0_11;
   wire [4:0] stage0_12;
   wire [3:0] stage0_13;
   wire [2:0] stage0_14;
   wire [1:0] stage0_15;
   wire [0:0] stage0_16;
   wire [0:0] stage1_0;
   wire [0:0] stage1_1;
   wire [0:0] stage1_2;
   wire [0:0] stage1_3;
   wire [5:0] stage1_4;
   wire [6:0] stage1_5;
   wire [0:0] stage1_6;
   wire [2:0] stage1_7;
   wire [4:0] stage1_8;
   wire [3:0] stage1_9;
   wire [8:0] stage1_10;
   wire [6:0] stage1_11;
   wire [4:0] stage1_12;
   wire [3:0] stage1_13;
   wire [2:0] stage1_14;
   wire [1:0] stage1_15;
   wire [0:0] stage1_16;
   wire [0:0] stage2_0;
   wire [0:0] stage2_1;
   wire [0:0] stage2_2;
   wire [0:0] stage2_3;
   wire [0:0] stage2_4;
   wire [5:0] stage2_5;
   wire [0:0] stage2_6;
   wire [1:0] stage2_7;
   wire [0:0] stage2_8;
   wire [2:0] stage2_9;
   wire [8:0] stage2_10;
   wire [1:0] stage2_11;
   wire [5:0] stage2_12;
   wire [0:0] stage2_13;
   wire [2:0] stage2_14;
   wire [2:0] stage2_15;
   wire [0:0] stage2_16;
   wire [0:0] stage3_0;
   wire [0:0] stage3_1;
   wire [0:0] stage3_2;
   wire [0:0] stage3_3;
   wire [0:0] stage3_4;
   wire [0:0] stage3_5;
   wire [0:0] stage3_6;
   wire [0:0] stage3_7;
   wire [0:0] stage3_8;
   wire [3:0] stage3_9;
   wire [2:0] stage3_10;
   wire [2:0] stage3_11;
   wire [0:0] stage3_12;
   wire [1:0] stage3_13;
   wire [3:0] stage3_14;
   wire [2:0] stage3_15;
   wire [0:0] stage3_16;
   wire [0:0] stage4_0;
   wire [0:0] stage4_1;
   wire [0:0] stage4_2;
   wire [0:0] stage4_3;
   wire [0:0] stage4_4;
   wire [0:0] stage4_5;
   wire [0:0] stage4_6;
   wire [0:0] stage4_7;
   wire [0:0] stage4_8;
   wire [0:0] stage4_9;
   wire [0:0] stage4_10;
   wire [0:0] stage4_11;
   wire [0:0] stage4_12;
   wire [2:0] stage4_13;
   wire [3:0] stage4_14;
   wire [2:0] stage4_15;
   wire [0:0] stage4_16;
   wire [0:0] stage5_0;
   wire [0:0] stage5_1;
   wire [0:0] stage5_2;
   wire [0:0] stage5_3;
   wire [0:0] stage5_4;
   wire [0:0] stage5_5;
   wire [0:0] stage5_6;
   wire [0:0] stage5_7;
   wire [0:0] stage5_8;
   wire [0:0] stage5_9;
   wire [0:0] stage5_10;
   wire [0:0] stage5_11;
   wire [0:0] stage5_12;
   wire [0:0] stage5_13;
   wire [0:0] stage5_14;
   wire [0:0] stage5_15;
   wire [0:0] stage5_16;
   wire [0:0] stage5_17;
   wire [0:0] stage6_0;
   wire [0:0] stage6_1;
   wire [0:0] stage6_2;
   wire [0:0] stage6_3;
   wire [0:0] stage6_4;
   wire [0:0] stage6_5;
   wire [0:0] stage6_6;
   wire [0:0] stage6_7;
   wire [0:0] stage6_8;
   wire [0:0] stage6_9;
   wire [0:0] stage6_10;
   wire [0:0] stage6_11;
   wire [0:0] stage6_12;
   wire [0:0] stage6_13;
   wire [0:0] stage6_14;
   wire [0:0] stage6_15;
   wire [0:0] stage6_16;
   wire [0:0] stage6_17;
   wire [0:0] stage7_0;
   wire [0:0] stage7_1;
   wire [0:0] stage7_2;
   wire [0:0] stage7_3;
   wire [0:0] stage7_4;
   wire [0:0] stage7_5;
   wire [0:0] stage7_6;
   wire [0:0] stage7_7;
   wire [0:0] stage7_8;
   wire [0:0] stage7_9;
   wire [0:0] stage7_10;
   wire [0:0] stage7_11;
   wire [0:0] stage7_12;
   wire [0:0] stage7_13;
   wire [0:0] stage7_14;
   wire [0:0] stage7_15;
   wire [0:0] stage7_16;
   wire [0:0] stage7_17;
   wire [0:0] stage8_0;
   wire [0:0] stage8_1;
   wire [0:0] stage8_2;
   wire [0:0] stage8_3;
   wire [0:0] stage8_4;
   wire [0:0] stage8_5;
   wire [0:0] stage8_6;
   wire [0:0] stage8_7;
   wire [0:0] stage8_8;
   wire [0:0] stage8_9;
   wire [0:0] stage8_10;
   wire [0:0] stage8_11;
   wire [0:0] stage8_12;
   wire [0:0] stage8_13;
   wire [0:0] stage8_14;
   wire [0:0] stage8_15;
   wire [0:0] stage8_16;
   wire [0:0] stage8_17;
   wire [0:0] stage9_0;
   wire [0:0] stage9_1;
   wire [0:0] stage9_2;
   wire [0:0] stage9_3;
   wire [0:0] stage9_4;
   wire [0:0] stage9_5;
   wire [0:0] stage9_6;
   wire [0:0] stage9_7;
   wire [0:0] stage9_8;
   wire [0:0] stage9_9;
   wire [0:0] stage9_10;
   wire [0:0] stage9_11;
   wire [0:0] stage9_12;
   wire [0:0] stage9_13;
   wire [0:0] stage9_14;
   wire [0:0] stage9_15;
   wire [0:0] stage9_16;
   wire [0:0] stage9_17;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign dst0 = stage9_0;
   assign dst1 = stage9_1;
   assign dst2 = stage9_2;
   assign dst3 = stage9_3;
   assign dst4 = stage9_4;
   assign dst5 = stage9_5;
   assign dst6 = stage9_6;
   assign dst7 = stage9_7;
   assign dst8 = stage9_8;
   assign dst9 = stage9_9;
   assign dst10 = stage9_10;
   assign dst11 = stage9_11;
   assign dst12 = stage9_12;
   assign dst13 = stage9_13;
   assign dst14 = stage9_14;
   assign dst15 = stage9_15;
   assign dst16 = stage9_16;
   assign dst17 = stage9_17;

   gpc433_5 gpc0 (
      {stage0_1[0], stage0_1[1], 1'b0},
      {stage0_2[0], stage0_2[1], stage0_2[2]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3]},
      {stage1_5[0],stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0]}
   );
   gpc607_5 gpc1 (
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[0],stage1_8[0],stage1_7[0],stage1_6[0]}
   );
   gpc607_5 gpc2 (
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[1],stage1_9[1],stage1_8[1],stage1_7[1]}
   );
   gpc1_1 gpc3 (
      {stage0_0[0]},
      {stage1_0[0]}
   );
   gpc1_1 gpc4 (
      {stage0_4[0]},
      {stage1_4[1]}
   );
   gpc1_1 gpc5 (
      {stage0_4[1]},
      {stage1_4[2]}
   );
   gpc1_1 gpc6 (
      {stage0_4[2]},
      {stage1_4[3]}
   );
   gpc1_1 gpc7 (
      {stage0_4[3]},
      {stage1_4[4]}
   );
   gpc1_1 gpc8 (
      {stage0_4[4]},
      {stage1_4[5]}
   );
   gpc1_1 gpc9 (
      {stage0_5[0]},
      {stage1_5[1]}
   );
   gpc1_1 gpc10 (
      {stage0_5[1]},
      {stage1_5[2]}
   );
   gpc1_1 gpc11 (
      {stage0_5[2]},
      {stage1_5[3]}
   );
   gpc1_1 gpc12 (
      {stage0_5[3]},
      {stage1_5[4]}
   );
   gpc1_1 gpc13 (
      {stage0_5[4]},
      {stage1_5[5]}
   );
   gpc1_1 gpc14 (
      {stage0_5[5]},
      {stage1_5[6]}
   );
   gpc1_1 gpc15 (
      {stage0_7[7]},
      {stage1_7[2]}
   );
   gpc1_1 gpc16 (
      {stage0_8[6]},
      {stage1_8[2]}
   );
   gpc1_1 gpc17 (
      {stage0_8[7]},
      {stage1_8[3]}
   );
   gpc1_1 gpc18 (
      {stage0_8[8]},
      {stage1_8[4]}
   );
   gpc1_1 gpc19 (
      {stage0_9[6]},
      {stage1_9[2]}
   );
   gpc1_1 gpc20 (
      {stage0_9[7]},
      {stage1_9[3]}
   );
   gpc1_1 gpc21 (
      {stage0_10[0]},
      {stage1_10[2]}
   );
   gpc1_1 gpc22 (
      {stage0_10[1]},
      {stage1_10[3]}
   );
   gpc1_1 gpc23 (
      {stage0_10[2]},
      {stage1_10[4]}
   );
   gpc1_1 gpc24 (
      {stage0_10[3]},
      {stage1_10[5]}
   );
   gpc1_1 gpc25 (
      {stage0_10[4]},
      {stage1_10[6]}
   );
   gpc1_1 gpc26 (
      {stage0_10[5]},
      {stage1_10[7]}
   );
   gpc1_1 gpc27 (
      {stage0_10[6]},
      {stage1_10[8]}
   );
   gpc1_1 gpc28 (
      {stage0_11[0]},
      {stage1_11[1]}
   );
   gpc1_1 gpc29 (
      {stage0_11[1]},
      {stage1_11[2]}
   );
   gpc1_1 gpc30 (
      {stage0_11[2]},
      {stage1_11[3]}
   );
   gpc1_1 gpc31 (
      {stage0_11[3]},
      {stage1_11[4]}
   );
   gpc1_1 gpc32 (
      {stage0_11[4]},
      {stage1_11[5]}
   );
   gpc1_1 gpc33 (
      {stage0_11[5]},
      {stage1_11[6]}
   );
   gpc1_1 gpc34 (
      {stage0_12[0]},
      {stage1_12[0]}
   );
   gpc1_1 gpc35 (
      {stage0_12[1]},
      {stage1_12[1]}
   );
   gpc1_1 gpc36 (
      {stage0_12[2]},
      {stage1_12[2]}
   );
   gpc1_1 gpc37 (
      {stage0_12[3]},
      {stage1_12[3]}
   );
   gpc1_1 gpc38 (
      {stage0_12[4]},
      {stage1_12[4]}
   );
   gpc1_1 gpc39 (
      {stage0_13[0]},
      {stage1_13[0]}
   );
   gpc1_1 gpc40 (
      {stage0_13[1]},
      {stage1_13[1]}
   );
   gpc1_1 gpc41 (
      {stage0_13[2]},
      {stage1_13[2]}
   );
   gpc1_1 gpc42 (
      {stage0_13[3]},
      {stage1_13[3]}
   );
   gpc1_1 gpc43 (
      {stage0_14[0]},
      {stage1_14[0]}
   );
   gpc1_1 gpc44 (
      {stage0_14[1]},
      {stage1_14[1]}
   );
   gpc1_1 gpc45 (
      {stage0_14[2]},
      {stage1_14[2]}
   );
   gpc1_1 gpc46 (
      {stage0_15[0]},
      {stage1_15[0]}
   );
   gpc1_1 gpc47 (
      {stage0_15[1]},
      {stage1_15[1]}
   );
   gpc1_1 gpc48 (
      {stage0_16[0]},
      {stage1_16[0]}
   );
   gpc126_4 gpc49 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_5[0], stage1_5[1]},
      {stage1_6[0]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[0]}
   );
   gpc1253_5 gpc50 (
      {stage1_7[0], stage1_7[1], stage1_7[2]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4]},
      {stage1_9[0], stage1_9[1]},
      {stage1_10[0]},
      {stage2_11[0],stage2_10[0],stage2_9[0],stage2_8[0],stage2_7[1]}
   );
   gpc1407_5 gpc51 (
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[0],stage2_13[0],stage2_12[0],stage2_11[1]}
   );
   gpc1_1 gpc52 (
      {stage1_0[0]},
      {stage2_0[0]}
   );
   gpc1_1 gpc53 (
      {stage1_1[0]},
      {stage2_1[0]}
   );
   gpc1_1 gpc54 (
      {stage1_2[0]},
      {stage2_2[0]}
   );
   gpc1_1 gpc55 (
      {stage1_3[0]},
      {stage2_3[0]}
   );
   gpc1_1 gpc56 (
      {stage1_5[2]},
      {stage2_5[1]}
   );
   gpc1_1 gpc57 (
      {stage1_5[3]},
      {stage2_5[2]}
   );
   gpc1_1 gpc58 (
      {stage1_5[4]},
      {stage2_5[3]}
   );
   gpc1_1 gpc59 (
      {stage1_5[5]},
      {stage2_5[4]}
   );
   gpc1_1 gpc60 (
      {stage1_5[6]},
      {stage2_5[5]}
   );
   gpc1_1 gpc61 (
      {stage1_9[2]},
      {stage2_9[1]}
   );
   gpc1_1 gpc62 (
      {stage1_9[3]},
      {stage2_9[2]}
   );
   gpc1_1 gpc63 (
      {stage1_10[1]},
      {stage2_10[1]}
   );
   gpc1_1 gpc64 (
      {stage1_10[2]},
      {stage2_10[2]}
   );
   gpc1_1 gpc65 (
      {stage1_10[3]},
      {stage2_10[3]}
   );
   gpc1_1 gpc66 (
      {stage1_10[4]},
      {stage2_10[4]}
   );
   gpc1_1 gpc67 (
      {stage1_10[5]},
      {stage2_10[5]}
   );
   gpc1_1 gpc68 (
      {stage1_10[6]},
      {stage2_10[6]}
   );
   gpc1_1 gpc69 (
      {stage1_10[7]},
      {stage2_10[7]}
   );
   gpc1_1 gpc70 (
      {stage1_10[8]},
      {stage2_10[8]}
   );
   gpc1_1 gpc71 (
      {stage1_12[0]},
      {stage2_12[1]}
   );
   gpc1_1 gpc72 (
      {stage1_12[1]},
      {stage2_12[2]}
   );
   gpc1_1 gpc73 (
      {stage1_12[2]},
      {stage2_12[3]}
   );
   gpc1_1 gpc74 (
      {stage1_12[3]},
      {stage2_12[4]}
   );
   gpc1_1 gpc75 (
      {stage1_12[4]},
      {stage2_12[5]}
   );
   gpc1_1 gpc76 (
      {stage1_14[1]},
      {stage2_14[1]}
   );
   gpc1_1 gpc77 (
      {stage1_14[2]},
      {stage2_14[2]}
   );
   gpc1_1 gpc78 (
      {stage1_15[0]},
      {stage2_15[1]}
   );
   gpc1_1 gpc79 (
      {stage1_15[1]},
      {stage2_15[2]}
   );
   gpc1_1 gpc80 (
      {stage1_16[0]},
      {stage2_16[0]}
   );
   gpc1316_5 gpc81 (
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage2_6[0]},
      {stage2_7[0], stage2_7[1], 1'b0},
      {stage2_8[0]},
      {stage3_9[0],stage3_8[0],stage3_7[0],stage3_6[0],stage3_5[0]}
   );
   gpc607_5 gpc82 (
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5], stage2_10[6]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[0],stage3_11[0],stage3_10[0]}
   );
   gpc1_1 gpc83 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc84 (
      {stage2_1[0]},
      {stage3_1[0]}
   );
   gpc1_1 gpc85 (
      {stage2_2[0]},
      {stage3_2[0]}
   );
   gpc1_1 gpc86 (
      {stage2_3[0]},
      {stage3_3[0]}
   );
   gpc1_1 gpc87 (
      {stage2_4[0]},
      {stage3_4[0]}
   );
   gpc1_1 gpc88 (
      {stage2_9[0]},
      {stage3_9[1]}
   );
   gpc1_1 gpc89 (
      {stage2_9[1]},
      {stage3_9[2]}
   );
   gpc1_1 gpc90 (
      {stage2_9[2]},
      {stage3_9[3]}
   );
   gpc1_1 gpc91 (
      {stage2_10[7]},
      {stage3_10[1]}
   );
   gpc1_1 gpc92 (
      {stage2_10[8]},
      {stage3_10[2]}
   );
   gpc1_1 gpc93 (
      {stage2_11[0]},
      {stage3_11[1]}
   );
   gpc1_1 gpc94 (
      {stage2_11[1]},
      {stage3_11[2]}
   );
   gpc1_1 gpc95 (
      {stage2_13[0]},
      {stage3_13[1]}
   );
   gpc1_1 gpc96 (
      {stage2_14[0]},
      {stage3_14[1]}
   );
   gpc1_1 gpc97 (
      {stage2_14[1]},
      {stage3_14[2]}
   );
   gpc1_1 gpc98 (
      {stage2_14[2]},
      {stage3_14[3]}
   );
   gpc1_1 gpc99 (
      {stage2_15[0]},
      {stage3_15[0]}
   );
   gpc1_1 gpc100 (
      {stage2_15[1]},
      {stage3_15[1]}
   );
   gpc1_1 gpc101 (
      {stage2_15[2]},
      {stage3_15[2]}
   );
   gpc1_1 gpc102 (
      {stage2_16[0]},
      {stage3_16[0]}
   );
   gpc1334_5 gpc103 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3]},
      {stage3_10[0], stage3_10[1], stage3_10[2]},
      {stage3_11[0], stage3_11[1], stage3_11[2]},
      {stage3_12[0]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[0]}
   );
   gpc1_1 gpc104 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc105 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc106 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc107 (
      {stage3_3[0]},
      {stage4_3[0]}
   );
   gpc1_1 gpc108 (
      {stage3_4[0]},
      {stage4_4[0]}
   );
   gpc1_1 gpc109 (
      {stage3_5[0]},
      {stage4_5[0]}
   );
   gpc1_1 gpc110 (
      {stage3_6[0]},
      {stage4_6[0]}
   );
   gpc1_1 gpc111 (
      {stage3_7[0]},
      {stage4_7[0]}
   );
   gpc1_1 gpc112 (
      {stage3_8[0]},
      {stage4_8[0]}
   );
   gpc1_1 gpc113 (
      {stage3_13[0]},
      {stage4_13[1]}
   );
   gpc1_1 gpc114 (
      {stage3_13[1]},
      {stage4_13[2]}
   );
   gpc1_1 gpc115 (
      {stage3_14[0]},
      {stage4_14[0]}
   );
   gpc1_1 gpc116 (
      {stage3_14[1]},
      {stage4_14[1]}
   );
   gpc1_1 gpc117 (
      {stage3_14[2]},
      {stage4_14[2]}
   );
   gpc1_1 gpc118 (
      {stage3_14[3]},
      {stage4_14[3]}
   );
   gpc1_1 gpc119 (
      {stage3_15[0]},
      {stage4_15[0]}
   );
   gpc1_1 gpc120 (
      {stage3_15[1]},
      {stage4_15[1]}
   );
   gpc1_1 gpc121 (
      {stage3_15[2]},
      {stage4_15[2]}
   );
   gpc1_1 gpc122 (
      {stage3_16[0]},
      {stage4_16[0]}
   );
   gpc1343_5 gpc123 (
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3]},
      {stage4_15[0], stage4_15[1], stage4_15[2]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[0]}
   );
   gpc1_1 gpc124 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc125 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc126 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc127 (
      {stage4_3[0]},
      {stage5_3[0]}
   );
   gpc1_1 gpc128 (
      {stage4_4[0]},
      {stage5_4[0]}
   );
   gpc1_1 gpc129 (
      {stage4_5[0]},
      {stage5_5[0]}
   );
   gpc1_1 gpc130 (
      {stage4_6[0]},
      {stage5_6[0]}
   );
   gpc1_1 gpc131 (
      {stage4_7[0]},
      {stage5_7[0]}
   );
   gpc1_1 gpc132 (
      {stage4_8[0]},
      {stage5_8[0]}
   );
   gpc1_1 gpc133 (
      {stage4_9[0]},
      {stage5_9[0]}
   );
   gpc1_1 gpc134 (
      {stage4_10[0]},
      {stage5_10[0]}
   );
   gpc1_1 gpc135 (
      {stage4_11[0]},
      {stage5_11[0]}
   );
   gpc1_1 gpc136 (
      {stage4_12[0]},
      {stage5_12[0]}
   );
   gpc1_1 gpc137 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc138 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc139 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc140 (
      {stage5_3[0]},
      {stage6_3[0]}
   );
   gpc1_1 gpc141 (
      {stage5_4[0]},
      {stage6_4[0]}
   );
   gpc1_1 gpc142 (
      {stage5_5[0]},
      {stage6_5[0]}
   );
   gpc1_1 gpc143 (
      {stage5_6[0]},
      {stage6_6[0]}
   );
   gpc1_1 gpc144 (
      {stage5_7[0]},
      {stage6_7[0]}
   );
   gpc1_1 gpc145 (
      {stage5_8[0]},
      {stage6_8[0]}
   );
   gpc1_1 gpc146 (
      {stage5_9[0]},
      {stage6_9[0]}
   );
   gpc1_1 gpc147 (
      {stage5_10[0]},
      {stage6_10[0]}
   );
   gpc1_1 gpc148 (
      {stage5_11[0]},
      {stage6_11[0]}
   );
   gpc1_1 gpc149 (
      {stage5_12[0]},
      {stage6_12[0]}
   );
   gpc1_1 gpc150 (
      {stage5_13[0]},
      {stage6_13[0]}
   );
   gpc1_1 gpc151 (
      {stage5_14[0]},
      {stage6_14[0]}
   );
   gpc1_1 gpc152 (
      {stage5_15[0]},
      {stage6_15[0]}
   );
   gpc1_1 gpc153 (
      {stage5_16[0]},
      {stage6_16[0]}
   );
   gpc1_1 gpc154 (
      {stage5_17[0]},
      {stage6_17[0]}
   );
   gpc1_1 gpc155 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc156 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc157 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc158 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc159 (
      {stage6_4[0]},
      {stage7_4[0]}
   );
   gpc1_1 gpc160 (
      {stage6_5[0]},
      {stage7_5[0]}
   );
   gpc1_1 gpc161 (
      {stage6_6[0]},
      {stage7_6[0]}
   );
   gpc1_1 gpc162 (
      {stage6_7[0]},
      {stage7_7[0]}
   );
   gpc1_1 gpc163 (
      {stage6_8[0]},
      {stage7_8[0]}
   );
   gpc1_1 gpc164 (
      {stage6_9[0]},
      {stage7_9[0]}
   );
   gpc1_1 gpc165 (
      {stage6_10[0]},
      {stage7_10[0]}
   );
   gpc1_1 gpc166 (
      {stage6_11[0]},
      {stage7_11[0]}
   );
   gpc1_1 gpc167 (
      {stage6_12[0]},
      {stage7_12[0]}
   );
   gpc1_1 gpc168 (
      {stage6_13[0]},
      {stage7_13[0]}
   );
   gpc1_1 gpc169 (
      {stage6_14[0]},
      {stage7_14[0]}
   );
   gpc1_1 gpc170 (
      {stage6_15[0]},
      {stage7_15[0]}
   );
   gpc1_1 gpc171 (
      {stage6_16[0]},
      {stage7_16[0]}
   );
   gpc1_1 gpc172 (
      {stage6_17[0]},
      {stage7_17[0]}
   );
   gpc1_1 gpc173 (
      {stage7_0[0]},
      {stage8_0[0]}
   );
   gpc1_1 gpc174 (
      {stage7_1[0]},
      {stage8_1[0]}
   );
   gpc1_1 gpc175 (
      {stage7_2[0]},
      {stage8_2[0]}
   );
   gpc1_1 gpc176 (
      {stage7_3[0]},
      {stage8_3[0]}
   );
   gpc1_1 gpc177 (
      {stage7_4[0]},
      {stage8_4[0]}
   );
   gpc1_1 gpc178 (
      {stage7_5[0]},
      {stage8_5[0]}
   );
   gpc1_1 gpc179 (
      {stage7_6[0]},
      {stage8_6[0]}
   );
   gpc1_1 gpc180 (
      {stage7_7[0]},
      {stage8_7[0]}
   );
   gpc1_1 gpc181 (
      {stage7_8[0]},
      {stage8_8[0]}
   );
   gpc1_1 gpc182 (
      {stage7_9[0]},
      {stage8_9[0]}
   );
   gpc1_1 gpc183 (
      {stage7_10[0]},
      {stage8_10[0]}
   );
   gpc1_1 gpc184 (
      {stage7_11[0]},
      {stage8_11[0]}
   );
   gpc1_1 gpc185 (
      {stage7_12[0]},
      {stage8_12[0]}
   );
   gpc1_1 gpc186 (
      {stage7_13[0]},
      {stage8_13[0]}
   );
   gpc1_1 gpc187 (
      {stage7_14[0]},
      {stage8_14[0]}
   );
   gpc1_1 gpc188 (
      {stage7_15[0]},
      {stage8_15[0]}
   );
   gpc1_1 gpc189 (
      {stage7_16[0]},
      {stage8_16[0]}
   );
   gpc1_1 gpc190 (
      {stage7_17[0]},
      {stage8_17[0]}
   );
   gpc1_1 gpc191 (
      {stage8_0[0]},
      {stage9_0[0]}
   );
   gpc1_1 gpc192 (
      {stage8_1[0]},
      {stage9_1[0]}
   );
   gpc1_1 gpc193 (
      {stage8_2[0]},
      {stage9_2[0]}
   );
   gpc1_1 gpc194 (
      {stage8_3[0]},
      {stage9_3[0]}
   );
   gpc1_1 gpc195 (
      {stage8_4[0]},
      {stage9_4[0]}
   );
   gpc1_1 gpc196 (
      {stage8_5[0]},
      {stage9_5[0]}
   );
   gpc1_1 gpc197 (
      {stage8_6[0]},
      {stage9_6[0]}
   );
   gpc1_1 gpc198 (
      {stage8_7[0]},
      {stage9_7[0]}
   );
   gpc1_1 gpc199 (
      {stage8_8[0]},
      {stage9_8[0]}
   );
   gpc1_1 gpc200 (
      {stage8_9[0]},
      {stage9_9[0]}
   );
   gpc1_1 gpc201 (
      {stage8_10[0]},
      {stage9_10[0]}
   );
   gpc1_1 gpc202 (
      {stage8_11[0]},
      {stage9_11[0]}
   );
   gpc1_1 gpc203 (
      {stage8_12[0]},
      {stage9_12[0]}
   );
   gpc1_1 gpc204 (
      {stage8_13[0]},
      {stage9_13[0]}
   );
   gpc1_1 gpc205 (
      {stage8_14[0]},
      {stage9_14[0]}
   );
   gpc1_1 gpc206 (
      {stage8_15[0]},
      {stage9_15[0]}
   );
   gpc1_1 gpc207 (
      {stage8_16[0]},
      {stage9_16[0]}
   );
   gpc1_1 gpc208 (
      {stage8_17[0]},
      {stage9_17[0]}
   );
endmodule
