module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24);
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    compressor2_1_486_16 compressor2_1_486_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24));
    initial begin
        src0 <= 486'h0;
        src1 <= 486'h0;
        src2 <= 486'h0;
        src3 <= 486'h0;
        src4 <= 486'h0;
        src5 <= 486'h0;
        src6 <= 486'h0;
        src7 <= 486'h0;
        src8 <= 486'h0;
        src9 <= 486'h0;
        src10 <= 486'h0;
        src11 <= 486'h0;
        src12 <= 486'h0;
        src13 <= 486'h0;
        src14 <= 486'h0;
        src15 <= 486'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor2_1_486_16(
    input [485:0]src0,
    input [485:0]src1,
    input [485:0]src2,
    input [485:0]src3,
    input [485:0]src4,
    input [485:0]src5,
    input [485:0]src6,
    input [485:0]src7,
    input [485:0]src8,
    input [485:0]src9,
    input [485:0]src10,
    input [485:0]src11,
    input [485:0]src12,
    input [485:0]src13,
    input [485:0]src14,
    input [485:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [0:0] comp_out24;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24)
    );
    rowadder2_1_25 rowadder2_1inst(
        .src0({comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [485:0] src0,
      input wire [485:0] src1,
      input wire [485:0] src2,
      input wire [485:0] src3,
      input wire [485:0] src4,
      input wire [485:0] src5,
      input wire [485:0] src6,
      input wire [485:0] src7,
      input wire [485:0] src8,
      input wire [485:0] src9,
      input wire [485:0] src10,
      input wire [485:0] src11,
      input wire [485:0] src12,
      input wire [485:0] src13,
      input wire [485:0] src14,
      input wire [485:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [0:0] dst24);

   wire [485:0] stage0_0;
   wire [485:0] stage0_1;
   wire [485:0] stage0_2;
   wire [485:0] stage0_3;
   wire [485:0] stage0_4;
   wire [485:0] stage0_5;
   wire [485:0] stage0_6;
   wire [485:0] stage0_7;
   wire [485:0] stage0_8;
   wire [485:0] stage0_9;
   wire [485:0] stage0_10;
   wire [485:0] stage0_11;
   wire [485:0] stage0_12;
   wire [485:0] stage0_13;
   wire [485:0] stage0_14;
   wire [485:0] stage0_15;
   wire [147:0] stage1_0;
   wire [134:0] stage1_1;
   wire [167:0] stage1_2;
   wire [243:0] stage1_3;
   wire [222:0] stage1_4;
   wire [336:0] stage1_5;
   wire [196:0] stage1_6;
   wire [216:0] stage1_7;
   wire [195:0] stage1_8;
   wire [210:0] stage1_9;
   wire [281:0] stage1_10;
   wire [213:0] stage1_11;
   wire [201:0] stage1_12;
   wire [234:0] stage1_13;
   wire [182:0] stage1_14;
   wire [154:0] stage1_15;
   wire [150:0] stage1_16;
   wire [80:0] stage1_17;
   wire [37:0] stage2_0;
   wire [62:0] stage2_1;
   wire [53:0] stage2_2;
   wire [85:0] stage2_3;
   wire [106:0] stage2_4;
   wire [107:0] stage2_5;
   wire [89:0] stage2_6;
   wire [102:0] stage2_7;
   wire [105:0] stage2_8;
   wire [80:0] stage2_9;
   wire [89:0] stage2_10;
   wire [106:0] stage2_11;
   wire [93:0] stage2_12;
   wire [85:0] stage2_13;
   wire [101:0] stage2_14;
   wire [74:0] stage2_15;
   wire [76:0] stage2_16;
   wire [95:0] stage2_17;
   wire [25:0] stage2_18;
   wire [4:0] stage2_19;
   wire [19:0] stage3_0;
   wire [14:0] stage3_1;
   wire [18:0] stage3_2;
   wire [40:0] stage3_3;
   wire [38:0] stage3_4;
   wire [39:0] stage3_5;
   wire [49:0] stage3_6;
   wire [35:0] stage3_7;
   wire [47:0] stage3_8;
   wire [42:0] stage3_9;
   wire [43:0] stage3_10;
   wire [37:0] stage3_11;
   wire [46:0] stage3_12;
   wire [39:0] stage3_13;
   wire [31:0] stage3_14;
   wire [43:0] stage3_15;
   wire [44:0] stage3_16;
   wire [29:0] stage3_17;
   wire [25:0] stage3_18;
   wire [18:0] stage3_19;
   wire [4:0] stage3_20;
   wire [0:0] stage3_21;
   wire [9:0] stage4_0;
   wire [5:0] stage4_1;
   wire [8:0] stage4_2;
   wire [9:0] stage4_3;
   wire [16:0] stage4_4;
   wire [14:0] stage4_5;
   wire [15:0] stage4_6;
   wire [20:0] stage4_7;
   wire [19:0] stage4_8;
   wire [15:0] stage4_9;
   wire [17:0] stage4_10;
   wire [18:0] stage4_11;
   wire [23:0] stage4_12;
   wire [16:0] stage4_13;
   wire [19:0] stage4_14;
   wire [27:0] stage4_15;
   wire [18:0] stage4_16;
   wire [12:0] stage4_17;
   wire [24:0] stage4_18;
   wire [13:0] stage4_19;
   wire [8:0] stage4_20;
   wire [2:0] stage4_21;
   wire [9:0] stage5_0;
   wire [5:0] stage5_1;
   wire [8:0] stage5_2;
   wire [5:0] stage5_3;
   wire [4:0] stage5_4;
   wire [3:0] stage5_5;
   wire [8:0] stage5_6;
   wire [8:0] stage5_7;
   wire [13:0] stage5_8;
   wire [8:0] stage5_9;
   wire [7:0] stage5_10;
   wire [6:0] stage5_11;
   wire [6:0] stage5_12;
   wire [9:0] stage5_13;
   wire [7:0] stage5_14;
   wire [9:0] stage5_15;
   wire [9:0] stage5_16;
   wire [7:0] stage5_17;
   wire [6:0] stage5_18;
   wire [10:0] stage5_19;
   wire [11:0] stage5_20;
   wire [3:0] stage5_21;
   wire [0:0] stage5_22;
   wire [5:0] stage6_0;
   wire [3:0] stage6_1;
   wire [4:0] stage6_2;
   wire [2:0] stage6_3;
   wire [5:0] stage6_4;
   wire [4:0] stage6_5;
   wire [2:0] stage6_6;
   wire [3:0] stage6_7;
   wire [3:0] stage6_8;
   wire [5:0] stage6_9;
   wire [4:0] stage6_10;
   wire [2:0] stage6_11;
   wire [1:0] stage6_12;
   wire [6:0] stage6_13;
   wire [3:0] stage6_14;
   wire [2:0] stage6_15;
   wire [5:0] stage6_16;
   wire [2:0] stage6_17;
   wire [5:0] stage6_18;
   wire [3:0] stage6_19;
   wire [4:0] stage6_20;
   wire [2:0] stage6_21;
   wire [2:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage7_0;
   wire [1:0] stage7_1;
   wire [1:0] stage7_2;
   wire [1:0] stage7_3;
   wire [1:0] stage7_4;
   wire [1:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [1:0] stage7_19;
   wire [1:0] stage7_20;
   wire [1:0] stage7_21;
   wire [1:0] stage7_22;
   wire [1:0] stage7_23;
   wire [0:0] stage7_24;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;
   assign dst21 = stage7_21;
   assign dst22 = stage7_22;
   assign dst23 = stage7_23;
   assign dst24 = stage7_24;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[10]},
      {stage0_3[20], stage0_3[21]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc2135_5 gpc11 (
      {stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59]},
      {stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[11]},
      {stage0_3[22], stage0_3[23]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[12]},
      {stage0_3[24]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[63], stage0_0[64], stage0_0[65]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[13]},
      {stage0_3[25]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[14]},
      {stage0_3[26]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[69], stage0_0[70], stage0_0[71]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[15]},
      {stage0_3[27]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[16]},
      {stage0_3[28]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[75], stage0_0[76], stage0_0[77]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[17]},
      {stage0_3[29]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_2[18]},
      {stage0_3[30]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_2[19]},
      {stage0_3[31]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_2[20]},
      {stage0_3[32]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[87], stage0_0[88], stage0_0[89]},
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_2[21]},
      {stage0_3[33]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_2[22]},
      {stage0_3[34]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[93], stage0_0[94], stage0_0[95]},
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_2[23]},
      {stage0_3[35]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_2[24]},
      {stage0_3[36]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[99], stage0_0[100], stage0_0[101]},
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_2[25]},
      {stage0_3[37]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_2[26]},
      {stage0_3[38]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[105], stage0_0[106], stage0_0[107]},
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_2[27]},
      {stage0_3[39]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_2[28]},
      {stage0_3[40]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[111], stage0_0[112], stage0_0[113]},
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_2[29]},
      {stage0_3[41]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_2[30]},
      {stage0_3[42]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[117], stage0_0[118], stage0_0[119]},
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_2[31]},
      {stage0_3[43]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[120], stage0_0[121], stage0_0[122]},
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_2[32]},
      {stage0_3[44]},
      {stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[123], stage0_0[124], stage0_0[125]},
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_2[33]},
      {stage0_3[45]},
      {stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[126], stage0_0[127], stage0_0[128]},
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_2[34]},
      {stage0_3[46]},
      {stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[129], stage0_0[130], stage0_0[131]},
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_2[35]},
      {stage0_3[47]},
      {stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[132], stage0_0[133], stage0_0[134]},
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_2[36]},
      {stage0_3[48]},
      {stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[159], stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163], stage0_0[164]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[165], stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169], stage0_0[170]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[171], stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175], stage0_0[176]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[177], stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[183], stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[189], stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200]},
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206]},
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212]},
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218]},
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224]},
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[225], stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230]},
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132]},
      {stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[231], stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236]},
      {stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138]},
      {stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[237], stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242]},
      {stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage1_4[54],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248]},
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150]},
      {stage1_4[55],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[249], stage0_0[250], stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254]},
      {stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage1_4[56],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[255], stage0_0[256], stage0_0[257], stage0_0[258], stage0_0[259], stage0_0[260]},
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162]},
      {stage1_4[57],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[261], stage0_0[262], stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266]},
      {stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168]},
      {stage1_4[58],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[267], stage0_0[268], stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272]},
      {stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174]},
      {stage1_4[59],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[273], stage0_0[274], stage0_0[275], stage0_0[276], stage0_0[277], stage0_0[278]},
      {stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180]},
      {stage1_4[60],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[279], stage0_0[280], stage0_0[281], stage0_0[282], stage0_0[283], stage0_0[284]},
      {stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186]},
      {stage1_4[61],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[285], stage0_0[286], stage0_0[287], stage0_0[288], stage0_0[289], stage0_0[290]},
      {stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192]},
      {stage1_4[62],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[291], stage0_0[292], stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296]},
      {stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198]},
      {stage1_4[63],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[297], stage0_0[298], stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302]},
      {stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204]},
      {stage1_4[64],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[303], stage0_0[304], stage0_0[305], stage0_0[306], stage0_0[307], stage0_0[308]},
      {stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210]},
      {stage1_4[65],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[309], stage0_0[310], stage0_0[311], stage0_0[312], stage0_0[313], stage0_0[314]},
      {stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216]},
      {stage1_4[66],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[315], stage0_0[316], stage0_0[317], stage0_0[318], stage0_0[319], stage0_0[320]},
      {stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222]},
      {stage1_4[67],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[321], stage0_0[322], stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326]},
      {stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228]},
      {stage1_4[68],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[327], stage0_0[328], stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332]},
      {stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234]},
      {stage1_4[69],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[333], stage0_0[334], stage0_0[335], stage0_0[336], stage0_0[337], stage0_0[338]},
      {stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240]},
      {stage1_4[70],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[339], stage0_0[340], stage0_0[341], stage0_0[342], stage0_0[343], stage0_0[344]},
      {stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246]},
      {stage1_4[71],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[345], stage0_0[346], stage0_0[347], stage0_0[348], stage0_0[349], stage0_0[350]},
      {stage0_2[247], stage0_2[248], stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252]},
      {stage1_4[72],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[351], stage0_0[352], stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356]},
      {stage0_2[253], stage0_2[254], stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258]},
      {stage1_4[73],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[357], stage0_0[358], stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362]},
      {stage0_2[259], stage0_2[260], stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264]},
      {stage1_4[74],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[363], stage0_0[364], stage0_0[365], stage0_0[366], stage0_0[367], stage0_0[368]},
      {stage0_2[265], stage0_2[266], stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270]},
      {stage1_4[75],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[369], stage0_0[370], stage0_0[371], stage0_0[372], stage0_0[373], stage0_0[374]},
      {stage0_2[271], stage0_2[272], stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276]},
      {stage1_4[76],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[375], stage0_0[376], stage0_0[377], stage0_0[378], stage0_0[379], stage0_0[380]},
      {stage0_2[277], stage0_2[278], stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282]},
      {stage1_4[77],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[381], stage0_0[382], stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386]},
      {stage0_2[283], stage0_2[284], stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288]},
      {stage1_4[78],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[387], stage0_0[388], stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392]},
      {stage0_2[289], stage0_2[290], stage0_2[291], stage0_2[292], stage0_2[293], stage0_2[294]},
      {stage1_4[79],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[393], stage0_0[394], stage0_0[395], stage0_0[396], stage0_0[397], stage0_0[398]},
      {stage0_2[295], stage0_2[296], stage0_2[297], stage0_2[298], stage0_2[299], stage0_2[300]},
      {stage1_4[80],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[399], stage0_0[400], stage0_0[401], stage0_0[402], stage0_0[403], stage0_0[404]},
      {stage0_2[301], stage0_2[302], stage0_2[303], stage0_2[304], stage0_2[305], stage0_2[306]},
      {stage1_4[81],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[405], stage0_0[406], stage0_0[407], stage0_0[408], stage0_0[409], stage0_0[410]},
      {stage0_2[307], stage0_2[308], stage0_2[309], stage0_2[310], stage0_2[311], stage0_2[312]},
      {stage1_4[82],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[411], stage0_0[412], stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416]},
      {stage0_2[313], stage0_2[314], stage0_2[315], stage0_2[316], stage0_2[317], stage0_2[318]},
      {stage1_4[83],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[417], stage0_0[418], stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422]},
      {stage0_2[319], stage0_2[320], stage0_2[321], stage0_2[322], stage0_2[323], stage0_2[324]},
      {stage1_4[84],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage1_5[0],stage1_4[85],stage1_3[85],stage1_2[85],stage1_1[85]}
   );
   gpc606_5 gpc86 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60]},
      {stage1_5[1],stage1_4[86],stage1_3[86],stage1_2[86],stage1_1[86]}
   );
   gpc606_5 gpc87 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66]},
      {stage1_5[2],stage1_4[87],stage1_3[87],stage1_2[87],stage1_1[87]}
   );
   gpc606_5 gpc88 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72]},
      {stage1_5[3],stage1_4[88],stage1_3[88],stage1_2[88],stage1_1[88]}
   );
   gpc606_5 gpc89 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78]},
      {stage1_5[4],stage1_4[89],stage1_3[89],stage1_2[89],stage1_1[89]}
   );
   gpc606_5 gpc90 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84]},
      {stage1_5[5],stage1_4[90],stage1_3[90],stage1_2[90],stage1_1[90]}
   );
   gpc606_5 gpc91 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90]},
      {stage1_5[6],stage1_4[91],stage1_3[91],stage1_2[91],stage1_1[91]}
   );
   gpc606_5 gpc92 (
      {stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233]},
      {stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage1_5[7],stage1_4[92],stage1_3[92],stage1_2[92],stage1_1[92]}
   );
   gpc606_5 gpc93 (
      {stage0_1[234], stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239]},
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102]},
      {stage1_5[8],stage1_4[93],stage1_3[93],stage1_2[93],stage1_1[93]}
   );
   gpc606_5 gpc94 (
      {stage0_1[240], stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245]},
      {stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108]},
      {stage1_5[9],stage1_4[94],stage1_3[94],stage1_2[94],stage1_1[94]}
   );
   gpc606_5 gpc95 (
      {stage0_1[246], stage0_1[247], stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251]},
      {stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114]},
      {stage1_5[10],stage1_4[95],stage1_3[95],stage1_2[95],stage1_1[95]}
   );
   gpc606_5 gpc96 (
      {stage0_1[252], stage0_1[253], stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257]},
      {stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120]},
      {stage1_5[11],stage1_4[96],stage1_3[96],stage1_2[96],stage1_1[96]}
   );
   gpc606_5 gpc97 (
      {stage0_1[258], stage0_1[259], stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263]},
      {stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126]},
      {stage1_5[12],stage1_4[97],stage1_3[97],stage1_2[97],stage1_1[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[264], stage0_1[265], stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269]},
      {stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132]},
      {stage1_5[13],stage1_4[98],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[270], stage0_1[271], stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275]},
      {stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138]},
      {stage1_5[14],stage1_4[99],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[276], stage0_1[277], stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281]},
      {stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144]},
      {stage1_5[15],stage1_4[100],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[282], stage0_1[283], stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287]},
      {stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150]},
      {stage1_5[16],stage1_4[101],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[288], stage0_1[289], stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293]},
      {stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156]},
      {stage1_5[17],stage1_4[102],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[294], stage0_1[295], stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299]},
      {stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162]},
      {stage1_5[18],stage1_4[103],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[300], stage0_1[301], stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305]},
      {stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168]},
      {stage1_5[19],stage1_4[104],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[306], stage0_1[307], stage0_1[308], stage0_1[309], stage0_1[310], stage0_1[311]},
      {stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174]},
      {stage1_5[20],stage1_4[105],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[312], stage0_1[313], stage0_1[314], stage0_1[315], stage0_1[316], stage0_1[317]},
      {stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180]},
      {stage1_5[21],stage1_4[106],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[318], stage0_1[319], stage0_1[320], stage0_1[321], stage0_1[322], stage0_1[323]},
      {stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186]},
      {stage1_5[22],stage1_4[107],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[324], stage0_1[325], stage0_1[326], stage0_1[327], stage0_1[328], stage0_1[329]},
      {stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192]},
      {stage1_5[23],stage1_4[108],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[330], stage0_1[331], stage0_1[332], stage0_1[333], stage0_1[334], stage0_1[335]},
      {stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198]},
      {stage1_5[24],stage1_4[109],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[336], stage0_1[337], stage0_1[338], stage0_1[339], stage0_1[340], stage0_1[341]},
      {stage0_3[199], stage0_3[200], stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204]},
      {stage1_5[25],stage1_4[110],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[342], stage0_1[343], stage0_1[344], stage0_1[345], stage0_1[346], stage0_1[347]},
      {stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210]},
      {stage1_5[26],stage1_4[111],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[348], stage0_1[349], stage0_1[350], stage0_1[351], stage0_1[352], stage0_1[353]},
      {stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216]},
      {stage1_5[27],stage1_4[112],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[354], stage0_1[355], stage0_1[356], stage0_1[357], stage0_1[358], stage0_1[359]},
      {stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220], stage0_3[221], stage0_3[222]},
      {stage1_5[28],stage1_4[113],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[360], stage0_1[361], stage0_1[362], stage0_1[363], stage0_1[364], stage0_1[365]},
      {stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226], stage0_3[227], stage0_3[228]},
      {stage1_5[29],stage1_4[114],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[366], stage0_1[367], stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371]},
      {stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234]},
      {stage1_5[30],stage1_4[115],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[372], stage0_1[373], stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377]},
      {stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240]},
      {stage1_5[31],stage1_4[116],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[378], stage0_1[379], stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383]},
      {stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246]},
      {stage1_5[32],stage1_4[117],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[384], stage0_1[385], stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389]},
      {stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250], stage0_3[251], stage0_3[252]},
      {stage1_5[33],stage1_4[118],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[390], stage0_1[391], stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395]},
      {stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256], stage0_3[257], stage0_3[258]},
      {stage1_5[34],stage1_4[119],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[396], stage0_1[397], stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401]},
      {stage0_3[259], stage0_3[260], stage0_3[261], stage0_3[262], stage0_3[263], stage0_3[264]},
      {stage1_5[35],stage1_4[120],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[402], stage0_1[403], stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407]},
      {stage0_3[265], stage0_3[266], stage0_3[267], stage0_3[268], stage0_3[269], stage0_3[270]},
      {stage1_5[36],stage1_4[121],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[408], stage0_1[409], stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413]},
      {stage0_3[271], stage0_3[272], stage0_3[273], stage0_3[274], stage0_3[275], stage0_3[276]},
      {stage1_5[37],stage1_4[122],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[414], stage0_1[415], stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419]},
      {stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280], stage0_3[281], stage0_3[282]},
      {stage1_5[38],stage1_4[123],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[420], stage0_1[421], stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425]},
      {stage0_3[283], stage0_3[284], stage0_3[285], stage0_3[286], stage0_3[287], stage0_3[288]},
      {stage1_5[39],stage1_4[124],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[426], stage0_1[427], stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431]},
      {stage0_3[289], stage0_3[290], stage0_3[291], stage0_3[292], stage0_3[293], stage0_3[294]},
      {stage1_5[40],stage1_4[125],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[432], stage0_1[433], stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437]},
      {stage0_3[295], stage0_3[296], stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300]},
      {stage1_5[41],stage1_4[126],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[438], stage0_1[439], stage0_1[440], stage0_1[441], stage0_1[442], stage0_1[443]},
      {stage0_3[301], stage0_3[302], stage0_3[303], stage0_3[304], stage0_3[305], stage0_3[306]},
      {stage1_5[42],stage1_4[127],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[444], stage0_1[445], stage0_1[446], stage0_1[447], stage0_1[448], stage0_1[449]},
      {stage0_3[307], stage0_3[308], stage0_3[309], stage0_3[310], stage0_3[311], stage0_3[312]},
      {stage1_5[43],stage1_4[128],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[450], stage0_1[451], stage0_1[452], stage0_1[453], stage0_1[454], stage0_1[455]},
      {stage0_3[313], stage0_3[314], stage0_3[315], stage0_3[316], stage0_3[317], stage0_3[318]},
      {stage1_5[44],stage1_4[129],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[456], stage0_1[457], stage0_1[458], stage0_1[459], stage0_1[460], stage0_1[461]},
      {stage0_3[319], stage0_3[320], stage0_3[321], stage0_3[322], stage0_3[323], stage0_3[324]},
      {stage1_5[45],stage1_4[130],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[462], stage0_1[463], stage0_1[464], stage0_1[465], stage0_1[466], stage0_1[467]},
      {stage0_3[325], stage0_3[326], stage0_3[327], stage0_3[328], stage0_3[329], stage0_3[330]},
      {stage1_5[46],stage1_4[131],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[468], stage0_1[469], stage0_1[470], stage0_1[471], stage0_1[472], stage0_1[473]},
      {stage0_3[331], stage0_3[332], stage0_3[333], stage0_3[334], stage0_3[335], stage0_3[336]},
      {stage1_5[47],stage1_4[132],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[474], stage0_1[475], stage0_1[476], stage0_1[477], stage0_1[478], stage0_1[479]},
      {stage0_3[337], stage0_3[338], stage0_3[339], stage0_3[340], stage0_3[341], stage0_3[342]},
      {stage1_5[48],stage1_4[133],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[480], stage0_1[481], stage0_1[482], stage0_1[483], stage0_1[484], stage0_1[485]},
      {stage0_3[343], stage0_3[344], stage0_3[345], stage0_3[346], stage0_3[347], stage0_3[348]},
      {stage1_5[49],stage1_4[134],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_2[325], stage0_2[326], stage0_2[327], stage0_2[328], stage0_2[329], stage0_2[330]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[50],stage1_4[135],stage1_3[135],stage1_2[135]}
   );
   gpc606_5 gpc136 (
      {stage0_2[331], stage0_2[332], stage0_2[333], stage0_2[334], stage0_2[335], stage0_2[336]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[51],stage1_4[136],stage1_3[136],stage1_2[136]}
   );
   gpc606_5 gpc137 (
      {stage0_2[337], stage0_2[338], stage0_2[339], stage0_2[340], stage0_2[341], stage0_2[342]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[52],stage1_4[137],stage1_3[137],stage1_2[137]}
   );
   gpc606_5 gpc138 (
      {stage0_2[343], stage0_2[344], stage0_2[345], stage0_2[346], stage0_2[347], stage0_2[348]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[53],stage1_4[138],stage1_3[138],stage1_2[138]}
   );
   gpc615_5 gpc139 (
      {stage0_2[349], stage0_2[350], stage0_2[351], stage0_2[352], stage0_2[353]},
      {stage0_3[349]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[54],stage1_4[139],stage1_3[139],stage1_2[139]}
   );
   gpc615_5 gpc140 (
      {stage0_2[354], stage0_2[355], stage0_2[356], stage0_2[357], stage0_2[358]},
      {stage0_3[350]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[55],stage1_4[140],stage1_3[140],stage1_2[140]}
   );
   gpc615_5 gpc141 (
      {stage0_2[359], stage0_2[360], stage0_2[361], stage0_2[362], stage0_2[363]},
      {stage0_3[351]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[56],stage1_4[141],stage1_3[141],stage1_2[141]}
   );
   gpc615_5 gpc142 (
      {stage0_2[364], stage0_2[365], stage0_2[366], stage0_2[367], stage0_2[368]},
      {stage0_3[352]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[57],stage1_4[142],stage1_3[142],stage1_2[142]}
   );
   gpc615_5 gpc143 (
      {stage0_2[369], stage0_2[370], stage0_2[371], stage0_2[372], stage0_2[373]},
      {stage0_3[353]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[58],stage1_4[143],stage1_3[143],stage1_2[143]}
   );
   gpc615_5 gpc144 (
      {stage0_2[374], stage0_2[375], stage0_2[376], stage0_2[377], stage0_2[378]},
      {stage0_3[354]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[59],stage1_4[144],stage1_3[144],stage1_2[144]}
   );
   gpc615_5 gpc145 (
      {stage0_2[379], stage0_2[380], stage0_2[381], stage0_2[382], stage0_2[383]},
      {stage0_3[355]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[60],stage1_4[145],stage1_3[145],stage1_2[145]}
   );
   gpc615_5 gpc146 (
      {stage0_2[384], stage0_2[385], stage0_2[386], stage0_2[387], stage0_2[388]},
      {stage0_3[356]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[61],stage1_4[146],stage1_3[146],stage1_2[146]}
   );
   gpc615_5 gpc147 (
      {stage0_2[389], stage0_2[390], stage0_2[391], stage0_2[392], stage0_2[393]},
      {stage0_3[357]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[62],stage1_4[147],stage1_3[147],stage1_2[147]}
   );
   gpc615_5 gpc148 (
      {stage0_2[394], stage0_2[395], stage0_2[396], stage0_2[397], stage0_2[398]},
      {stage0_3[358]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[63],stage1_4[148],stage1_3[148],stage1_2[148]}
   );
   gpc615_5 gpc149 (
      {stage0_2[399], stage0_2[400], stage0_2[401], stage0_2[402], stage0_2[403]},
      {stage0_3[359]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[64],stage1_4[149],stage1_3[149],stage1_2[149]}
   );
   gpc615_5 gpc150 (
      {stage0_2[404], stage0_2[405], stage0_2[406], stage0_2[407], stage0_2[408]},
      {stage0_3[360]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[65],stage1_4[150],stage1_3[150],stage1_2[150]}
   );
   gpc615_5 gpc151 (
      {stage0_2[409], stage0_2[410], stage0_2[411], stage0_2[412], stage0_2[413]},
      {stage0_3[361]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[66],stage1_4[151],stage1_3[151],stage1_2[151]}
   );
   gpc615_5 gpc152 (
      {stage0_2[414], stage0_2[415], stage0_2[416], stage0_2[417], stage0_2[418]},
      {stage0_3[362]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[67],stage1_4[152],stage1_3[152],stage1_2[152]}
   );
   gpc615_5 gpc153 (
      {stage0_2[419], stage0_2[420], stage0_2[421], stage0_2[422], stage0_2[423]},
      {stage0_3[363]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage1_6[18],stage1_5[68],stage1_4[153],stage1_3[153],stage1_2[153]}
   );
   gpc615_5 gpc154 (
      {stage0_2[424], stage0_2[425], stage0_2[426], stage0_2[427], stage0_2[428]},
      {stage0_3[364]},
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage1_6[19],stage1_5[69],stage1_4[154],stage1_3[154],stage1_2[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[429], stage0_2[430], stage0_2[431], stage0_2[432], stage0_2[433]},
      {stage0_3[365]},
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage1_6[20],stage1_5[70],stage1_4[155],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[434], stage0_2[435], stage0_2[436], stage0_2[437], stage0_2[438]},
      {stage0_3[366]},
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage1_6[21],stage1_5[71],stage1_4[156],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_2[439], stage0_2[440], stage0_2[441], stage0_2[442], stage0_2[443]},
      {stage0_3[367]},
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage1_6[22],stage1_5[72],stage1_4[157],stage1_3[157],stage1_2[157]}
   );
   gpc615_5 gpc158 (
      {stage0_2[444], stage0_2[445], stage0_2[446], stage0_2[447], stage0_2[448]},
      {stage0_3[368]},
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage1_6[23],stage1_5[73],stage1_4[158],stage1_3[158],stage1_2[158]}
   );
   gpc615_5 gpc159 (
      {stage0_2[449], stage0_2[450], stage0_2[451], stage0_2[452], stage0_2[453]},
      {stage0_3[369]},
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage1_6[24],stage1_5[74],stage1_4[159],stage1_3[159],stage1_2[159]}
   );
   gpc615_5 gpc160 (
      {stage0_2[454], stage0_2[455], stage0_2[456], stage0_2[457], stage0_2[458]},
      {stage0_3[370]},
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage1_6[25],stage1_5[75],stage1_4[160],stage1_3[160],stage1_2[160]}
   );
   gpc615_5 gpc161 (
      {stage0_2[459], stage0_2[460], stage0_2[461], stage0_2[462], stage0_2[463]},
      {stage0_3[371]},
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage1_6[26],stage1_5[76],stage1_4[161],stage1_3[161],stage1_2[161]}
   );
   gpc615_5 gpc162 (
      {stage0_2[464], stage0_2[465], stage0_2[466], stage0_2[467], stage0_2[468]},
      {stage0_3[372]},
      {stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167]},
      {stage1_6[27],stage1_5[77],stage1_4[162],stage1_3[162],stage1_2[162]}
   );
   gpc615_5 gpc163 (
      {stage0_2[469], stage0_2[470], stage0_2[471], stage0_2[472], stage0_2[473]},
      {stage0_3[373]},
      {stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173]},
      {stage1_6[28],stage1_5[78],stage1_4[163],stage1_3[163],stage1_2[163]}
   );
   gpc615_5 gpc164 (
      {stage0_2[474], stage0_2[475], stage0_2[476], stage0_2[477], stage0_2[478]},
      {stage0_3[374]},
      {stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178], stage0_4[179]},
      {stage1_6[29],stage1_5[79],stage1_4[164],stage1_3[164],stage1_2[164]}
   );
   gpc615_5 gpc165 (
      {stage0_2[479], stage0_2[480], stage0_2[481], stage0_2[482], stage0_2[483]},
      {stage0_3[375]},
      {stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184], stage0_4[185]},
      {stage1_6[30],stage1_5[80],stage1_4[165],stage1_3[165],stage1_2[165]}
   );
   gpc615_5 gpc166 (
      {stage0_3[376], stage0_3[377], stage0_3[378], stage0_3[379], stage0_3[380]},
      {stage0_4[186]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[31],stage1_5[81],stage1_4[166],stage1_3[166]}
   );
   gpc615_5 gpc167 (
      {stage0_3[381], stage0_3[382], stage0_3[383], stage0_3[384], stage0_3[385]},
      {stage0_4[187]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[32],stage1_5[82],stage1_4[167],stage1_3[167]}
   );
   gpc615_5 gpc168 (
      {stage0_3[386], stage0_3[387], stage0_3[388], stage0_3[389], stage0_3[390]},
      {stage0_4[188]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[33],stage1_5[83],stage1_4[168],stage1_3[168]}
   );
   gpc615_5 gpc169 (
      {stage0_3[391], stage0_3[392], stage0_3[393], stage0_3[394], stage0_3[395]},
      {stage0_4[189]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[34],stage1_5[84],stage1_4[169],stage1_3[169]}
   );
   gpc615_5 gpc170 (
      {stage0_3[396], stage0_3[397], stage0_3[398], stage0_3[399], stage0_3[400]},
      {stage0_4[190]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[35],stage1_5[85],stage1_4[170],stage1_3[170]}
   );
   gpc615_5 gpc171 (
      {stage0_3[401], stage0_3[402], stage0_3[403], stage0_3[404], stage0_3[405]},
      {stage0_4[191]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[36],stage1_5[86],stage1_4[171],stage1_3[171]}
   );
   gpc615_5 gpc172 (
      {stage0_3[406], stage0_3[407], stage0_3[408], stage0_3[409], stage0_3[410]},
      {stage0_4[192]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[37],stage1_5[87],stage1_4[172],stage1_3[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[411], stage0_3[412], stage0_3[413], stage0_3[414], stage0_3[415]},
      {stage0_4[193]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[38],stage1_5[88],stage1_4[173],stage1_3[173]}
   );
   gpc606_5 gpc174 (
      {stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[8],stage1_6[39],stage1_5[89],stage1_4[174]}
   );
   gpc606_5 gpc175 (
      {stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[9],stage1_6[40],stage1_5[90],stage1_4[175]}
   );
   gpc606_5 gpc176 (
      {stage0_4[206], stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[10],stage1_6[41],stage1_5[91],stage1_4[176]}
   );
   gpc606_5 gpc177 (
      {stage0_4[212], stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[11],stage1_6[42],stage1_5[92],stage1_4[177]}
   );
   gpc606_5 gpc178 (
      {stage0_4[218], stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[12],stage1_6[43],stage1_5[93],stage1_4[178]}
   );
   gpc606_5 gpc179 (
      {stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[13],stage1_6[44],stage1_5[94],stage1_4[179]}
   );
   gpc606_5 gpc180 (
      {stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[14],stage1_6[45],stage1_5[95],stage1_4[180]}
   );
   gpc606_5 gpc181 (
      {stage0_4[236], stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[15],stage1_6[46],stage1_5[96],stage1_4[181]}
   );
   gpc606_5 gpc182 (
      {stage0_4[242], stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[16],stage1_6[47],stage1_5[97],stage1_4[182]}
   );
   gpc606_5 gpc183 (
      {stage0_4[248], stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[17],stage1_6[48],stage1_5[98],stage1_4[183]}
   );
   gpc606_5 gpc184 (
      {stage0_4[254], stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258], stage0_4[259]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[18],stage1_6[49],stage1_5[99],stage1_4[184]}
   );
   gpc606_5 gpc185 (
      {stage0_4[260], stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264], stage0_4[265]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[19],stage1_6[50],stage1_5[100],stage1_4[185]}
   );
   gpc606_5 gpc186 (
      {stage0_4[266], stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270], stage0_4[271]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[20],stage1_6[51],stage1_5[101],stage1_4[186]}
   );
   gpc606_5 gpc187 (
      {stage0_4[272], stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276], stage0_4[277]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[21],stage1_6[52],stage1_5[102],stage1_4[187]}
   );
   gpc606_5 gpc188 (
      {stage0_4[278], stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282], stage0_4[283]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[22],stage1_6[53],stage1_5[103],stage1_4[188]}
   );
   gpc606_5 gpc189 (
      {stage0_4[284], stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288], stage0_4[289]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[23],stage1_6[54],stage1_5[104],stage1_4[189]}
   );
   gpc606_5 gpc190 (
      {stage0_4[290], stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294], stage0_4[295]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[24],stage1_6[55],stage1_5[105],stage1_4[190]}
   );
   gpc606_5 gpc191 (
      {stage0_4[296], stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300], stage0_4[301]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[25],stage1_6[56],stage1_5[106],stage1_4[191]}
   );
   gpc606_5 gpc192 (
      {stage0_4[302], stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306], stage0_4[307]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[26],stage1_6[57],stage1_5[107],stage1_4[192]}
   );
   gpc606_5 gpc193 (
      {stage0_4[308], stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312], stage0_4[313]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[27],stage1_6[58],stage1_5[108],stage1_4[193]}
   );
   gpc606_5 gpc194 (
      {stage0_4[314], stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318], stage0_4[319]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[28],stage1_6[59],stage1_5[109],stage1_4[194]}
   );
   gpc606_5 gpc195 (
      {stage0_4[320], stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324], stage0_4[325]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[29],stage1_6[60],stage1_5[110],stage1_4[195]}
   );
   gpc606_5 gpc196 (
      {stage0_4[326], stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330], stage0_4[331]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[30],stage1_6[61],stage1_5[111],stage1_4[196]}
   );
   gpc606_5 gpc197 (
      {stage0_4[332], stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336], stage0_4[337]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[31],stage1_6[62],stage1_5[112],stage1_4[197]}
   );
   gpc606_5 gpc198 (
      {stage0_4[338], stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342], stage0_4[343]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[32],stage1_6[63],stage1_5[113],stage1_4[198]}
   );
   gpc606_5 gpc199 (
      {stage0_4[344], stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348], stage0_4[349]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[33],stage1_6[64],stage1_5[114],stage1_4[199]}
   );
   gpc606_5 gpc200 (
      {stage0_4[350], stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354], stage0_4[355]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[34],stage1_6[65],stage1_5[115],stage1_4[200]}
   );
   gpc606_5 gpc201 (
      {stage0_4[356], stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360], stage0_4[361]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[35],stage1_6[66],stage1_5[116],stage1_4[201]}
   );
   gpc606_5 gpc202 (
      {stage0_4[362], stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366], stage0_4[367]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[36],stage1_6[67],stage1_5[117],stage1_4[202]}
   );
   gpc606_5 gpc203 (
      {stage0_4[368], stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372], stage0_4[373]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[37],stage1_6[68],stage1_5[118],stage1_4[203]}
   );
   gpc606_5 gpc204 (
      {stage0_4[374], stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378], stage0_4[379]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[38],stage1_6[69],stage1_5[119],stage1_4[204]}
   );
   gpc606_5 gpc205 (
      {stage0_4[380], stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384], stage0_4[385]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[39],stage1_6[70],stage1_5[120],stage1_4[205]}
   );
   gpc606_5 gpc206 (
      {stage0_4[386], stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390], stage0_4[391]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[40],stage1_6[71],stage1_5[121],stage1_4[206]}
   );
   gpc606_5 gpc207 (
      {stage0_4[392], stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396], stage0_4[397]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[41],stage1_6[72],stage1_5[122],stage1_4[207]}
   );
   gpc606_5 gpc208 (
      {stage0_4[398], stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402], stage0_4[403]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[42],stage1_6[73],stage1_5[123],stage1_4[208]}
   );
   gpc606_5 gpc209 (
      {stage0_4[404], stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408], stage0_4[409]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[43],stage1_6[74],stage1_5[124],stage1_4[209]}
   );
   gpc606_5 gpc210 (
      {stage0_4[410], stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414], stage0_4[415]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[44],stage1_6[75],stage1_5[125],stage1_4[210]}
   );
   gpc606_5 gpc211 (
      {stage0_4[416], stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420], stage0_4[421]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[45],stage1_6[76],stage1_5[126],stage1_4[211]}
   );
   gpc606_5 gpc212 (
      {stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426], stage0_4[427]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[46],stage1_6[77],stage1_5[127],stage1_4[212]}
   );
   gpc606_5 gpc213 (
      {stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431], stage0_4[432], stage0_4[433]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[47],stage1_6[78],stage1_5[128],stage1_4[213]}
   );
   gpc606_5 gpc214 (
      {stage0_4[434], stage0_4[435], stage0_4[436], stage0_4[437], stage0_4[438], stage0_4[439]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[48],stage1_6[79],stage1_5[129],stage1_4[214]}
   );
   gpc606_5 gpc215 (
      {stage0_4[440], stage0_4[441], stage0_4[442], stage0_4[443], stage0_4[444], stage0_4[445]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[49],stage1_6[80],stage1_5[130],stage1_4[215]}
   );
   gpc606_5 gpc216 (
      {stage0_4[446], stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450], stage0_4[451]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[50],stage1_6[81],stage1_5[131],stage1_4[216]}
   );
   gpc606_5 gpc217 (
      {stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455], stage0_4[456], stage0_4[457]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[51],stage1_6[82],stage1_5[132],stage1_4[217]}
   );
   gpc606_5 gpc218 (
      {stage0_4[458], stage0_4[459], stage0_4[460], stage0_4[461], stage0_4[462], stage0_4[463]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[52],stage1_6[83],stage1_5[133],stage1_4[218]}
   );
   gpc606_5 gpc219 (
      {stage0_4[464], stage0_4[465], stage0_4[466], stage0_4[467], stage0_4[468], stage0_4[469]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[53],stage1_6[84],stage1_5[134],stage1_4[219]}
   );
   gpc606_5 gpc220 (
      {stage0_4[470], stage0_4[471], stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[54],stage1_6[85],stage1_5[135],stage1_4[220]}
   );
   gpc615_5 gpc221 (
      {stage0_4[476], stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480]},
      {stage0_5[48]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[55],stage1_6[86],stage1_5[136],stage1_4[221]}
   );
   gpc615_5 gpc222 (
      {stage0_4[481], stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485]},
      {stage0_5[49]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[56],stage1_6[87],stage1_5[137],stage1_4[222]}
   );
   gpc606_5 gpc223 (
      {stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53], stage0_5[54], stage0_5[55]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[49],stage1_7[57],stage1_6[88],stage1_5[138]}
   );
   gpc606_5 gpc224 (
      {stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60], stage0_5[61]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[50],stage1_7[58],stage1_6[89],stage1_5[139]}
   );
   gpc606_5 gpc225 (
      {stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65], stage0_5[66], stage0_5[67]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[51],stage1_7[59],stage1_6[90],stage1_5[140]}
   );
   gpc606_5 gpc226 (
      {stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71], stage0_5[72], stage0_5[73]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[52],stage1_7[60],stage1_6[91],stage1_5[141]}
   );
   gpc606_5 gpc227 (
      {stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77], stage0_5[78], stage0_5[79]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[53],stage1_7[61],stage1_6[92],stage1_5[142]}
   );
   gpc606_5 gpc228 (
      {stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83], stage0_5[84], stage0_5[85]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[54],stage1_7[62],stage1_6[93],stage1_5[143]}
   );
   gpc606_5 gpc229 (
      {stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89], stage0_5[90], stage0_5[91]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[55],stage1_7[63],stage1_6[94],stage1_5[144]}
   );
   gpc606_5 gpc230 (
      {stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95], stage0_5[96], stage0_5[97]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[56],stage1_7[64],stage1_6[95],stage1_5[145]}
   );
   gpc606_5 gpc231 (
      {stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102], stage0_5[103]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[57],stage1_7[65],stage1_6[96],stage1_5[146]}
   );
   gpc606_5 gpc232 (
      {stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107], stage0_5[108], stage0_5[109]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[58],stage1_7[66],stage1_6[97],stage1_5[147]}
   );
   gpc606_5 gpc233 (
      {stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113], stage0_5[114], stage0_5[115]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[59],stage1_7[67],stage1_6[98],stage1_5[148]}
   );
   gpc606_5 gpc234 (
      {stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119], stage0_5[120], stage0_5[121]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[60],stage1_7[68],stage1_6[99],stage1_5[149]}
   );
   gpc606_5 gpc235 (
      {stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126], stage0_5[127]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[61],stage1_7[69],stage1_6[100],stage1_5[150]}
   );
   gpc606_5 gpc236 (
      {stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131], stage0_5[132], stage0_5[133]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[62],stage1_7[70],stage1_6[101],stage1_5[151]}
   );
   gpc606_5 gpc237 (
      {stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137], stage0_5[138], stage0_5[139]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[63],stage1_7[71],stage1_6[102],stage1_5[152]}
   );
   gpc606_5 gpc238 (
      {stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143], stage0_5[144], stage0_5[145]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[64],stage1_7[72],stage1_6[103],stage1_5[153]}
   );
   gpc606_5 gpc239 (
      {stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150], stage0_5[151]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[65],stage1_7[73],stage1_6[104],stage1_5[154]}
   );
   gpc606_5 gpc240 (
      {stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156], stage0_5[157]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[66],stage1_7[74],stage1_6[105],stage1_5[155]}
   );
   gpc606_5 gpc241 (
      {stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161], stage0_5[162], stage0_5[163]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[67],stage1_7[75],stage1_6[106],stage1_5[156]}
   );
   gpc606_5 gpc242 (
      {stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167], stage0_5[168], stage0_5[169]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[68],stage1_7[76],stage1_6[107],stage1_5[157]}
   );
   gpc606_5 gpc243 (
      {stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173], stage0_5[174], stage0_5[175]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[69],stage1_7[77],stage1_6[108],stage1_5[158]}
   );
   gpc606_5 gpc244 (
      {stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179], stage0_5[180], stage0_5[181]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[70],stage1_7[78],stage1_6[109],stage1_5[159]}
   );
   gpc606_5 gpc245 (
      {stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186], stage0_5[187]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[71],stage1_7[79],stage1_6[110],stage1_5[160]}
   );
   gpc606_5 gpc246 (
      {stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192], stage0_5[193]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[72],stage1_7[80],stage1_6[111],stage1_5[161]}
   );
   gpc606_5 gpc247 (
      {stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198], stage0_5[199]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[73],stage1_7[81],stage1_6[112],stage1_5[162]}
   );
   gpc606_5 gpc248 (
      {stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204], stage0_5[205]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[74],stage1_7[82],stage1_6[113],stage1_5[163]}
   );
   gpc606_5 gpc249 (
      {stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210], stage0_5[211]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[75],stage1_7[83],stage1_6[114],stage1_5[164]}
   );
   gpc606_5 gpc250 (
      {stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216], stage0_5[217]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[76],stage1_7[84],stage1_6[115],stage1_5[165]}
   );
   gpc606_5 gpc251 (
      {stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222], stage0_5[223]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[77],stage1_7[85],stage1_6[116],stage1_5[166]}
   );
   gpc606_5 gpc252 (
      {stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228], stage0_5[229]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[78],stage1_7[86],stage1_6[117],stage1_5[167]}
   );
   gpc606_5 gpc253 (
      {stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234], stage0_5[235]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[79],stage1_7[87],stage1_6[118],stage1_5[168]}
   );
   gpc606_5 gpc254 (
      {stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239], stage0_5[240], stage0_5[241]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[80],stage1_7[88],stage1_6[119],stage1_5[169]}
   );
   gpc606_5 gpc255 (
      {stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245], stage0_5[246], stage0_5[247]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[81],stage1_7[89],stage1_6[120],stage1_5[170]}
   );
   gpc606_5 gpc256 (
      {stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251], stage0_5[252], stage0_5[253]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[82],stage1_7[90],stage1_6[121],stage1_5[171]}
   );
   gpc606_5 gpc257 (
      {stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257], stage0_5[258], stage0_5[259]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[83],stage1_7[91],stage1_6[122],stage1_5[172]}
   );
   gpc606_5 gpc258 (
      {stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263], stage0_5[264], stage0_5[265]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[84],stage1_7[92],stage1_6[123],stage1_5[173]}
   );
   gpc606_5 gpc259 (
      {stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269], stage0_5[270], stage0_5[271]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[85],stage1_7[93],stage1_6[124],stage1_5[174]}
   );
   gpc615_5 gpc260 (
      {stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275], stage0_5[276]},
      {stage0_6[294]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[86],stage1_7[94],stage1_6[125],stage1_5[175]}
   );
   gpc615_5 gpc261 (
      {stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281]},
      {stage0_6[295]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[87],stage1_7[95],stage1_6[126],stage1_5[176]}
   );
   gpc615_5 gpc262 (
      {stage0_5[282], stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286]},
      {stage0_6[296]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[88],stage1_7[96],stage1_6[127],stage1_5[177]}
   );
   gpc615_5 gpc263 (
      {stage0_5[287], stage0_5[288], stage0_5[289], stage0_5[290], stage0_5[291]},
      {stage0_6[297]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[89],stage1_7[97],stage1_6[128],stage1_5[178]}
   );
   gpc615_5 gpc264 (
      {stage0_5[292], stage0_5[293], stage0_5[294], stage0_5[295], stage0_5[296]},
      {stage0_6[298]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[90],stage1_7[98],stage1_6[129],stage1_5[179]}
   );
   gpc615_5 gpc265 (
      {stage0_5[297], stage0_5[298], stage0_5[299], stage0_5[300], stage0_5[301]},
      {stage0_6[299]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[91],stage1_7[99],stage1_6[130],stage1_5[180]}
   );
   gpc615_5 gpc266 (
      {stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305], stage0_5[306]},
      {stage0_6[300]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[92],stage1_7[100],stage1_6[131],stage1_5[181]}
   );
   gpc615_5 gpc267 (
      {stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311]},
      {stage0_6[301]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[93],stage1_7[101],stage1_6[132],stage1_5[182]}
   );
   gpc615_5 gpc268 (
      {stage0_5[312], stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316]},
      {stage0_6[302]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[94],stage1_7[102],stage1_6[133],stage1_5[183]}
   );
   gpc615_5 gpc269 (
      {stage0_5[317], stage0_5[318], stage0_5[319], stage0_5[320], stage0_5[321]},
      {stage0_6[303]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[95],stage1_7[103],stage1_6[134],stage1_5[184]}
   );
   gpc615_5 gpc270 (
      {stage0_5[322], stage0_5[323], stage0_5[324], stage0_5[325], stage0_5[326]},
      {stage0_6[304]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[96],stage1_7[104],stage1_6[135],stage1_5[185]}
   );
   gpc615_5 gpc271 (
      {stage0_5[327], stage0_5[328], stage0_5[329], stage0_5[330], stage0_5[331]},
      {stage0_6[305]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[97],stage1_7[105],stage1_6[136],stage1_5[186]}
   );
   gpc615_5 gpc272 (
      {stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335], stage0_5[336]},
      {stage0_6[306]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[98],stage1_7[106],stage1_6[137],stage1_5[187]}
   );
   gpc615_5 gpc273 (
      {stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage0_7[300]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[50],stage1_8[99],stage1_7[107],stage1_6[138]}
   );
   gpc615_5 gpc274 (
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316]},
      {stage0_7[301]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[51],stage1_8[100],stage1_7[108],stage1_6[139]}
   );
   gpc615_5 gpc275 (
      {stage0_6[317], stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321]},
      {stage0_7[302]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[52],stage1_8[101],stage1_7[109],stage1_6[140]}
   );
   gpc615_5 gpc276 (
      {stage0_6[322], stage0_6[323], stage0_6[324], stage0_6[325], stage0_6[326]},
      {stage0_7[303]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[53],stage1_8[102],stage1_7[110],stage1_6[141]}
   );
   gpc615_5 gpc277 (
      {stage0_6[327], stage0_6[328], stage0_6[329], stage0_6[330], stage0_6[331]},
      {stage0_7[304]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[54],stage1_8[103],stage1_7[111],stage1_6[142]}
   );
   gpc615_5 gpc278 (
      {stage0_6[332], stage0_6[333], stage0_6[334], stage0_6[335], stage0_6[336]},
      {stage0_7[305]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[55],stage1_8[104],stage1_7[112],stage1_6[143]}
   );
   gpc615_5 gpc279 (
      {stage0_6[337], stage0_6[338], stage0_6[339], stage0_6[340], stage0_6[341]},
      {stage0_7[306]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[56],stage1_8[105],stage1_7[113],stage1_6[144]}
   );
   gpc615_5 gpc280 (
      {stage0_6[342], stage0_6[343], stage0_6[344], stage0_6[345], stage0_6[346]},
      {stage0_7[307]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[57],stage1_8[106],stage1_7[114],stage1_6[145]}
   );
   gpc615_5 gpc281 (
      {stage0_6[347], stage0_6[348], stage0_6[349], stage0_6[350], stage0_6[351]},
      {stage0_7[308]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[58],stage1_8[107],stage1_7[115],stage1_6[146]}
   );
   gpc615_5 gpc282 (
      {stage0_6[352], stage0_6[353], stage0_6[354], stage0_6[355], stage0_6[356]},
      {stage0_7[309]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[59],stage1_8[108],stage1_7[116],stage1_6[147]}
   );
   gpc615_5 gpc283 (
      {stage0_6[357], stage0_6[358], stage0_6[359], stage0_6[360], stage0_6[361]},
      {stage0_7[310]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[60],stage1_8[109],stage1_7[117],stage1_6[148]}
   );
   gpc615_5 gpc284 (
      {stage0_6[362], stage0_6[363], stage0_6[364], stage0_6[365], stage0_6[366]},
      {stage0_7[311]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[61],stage1_8[110],stage1_7[118],stage1_6[149]}
   );
   gpc615_5 gpc285 (
      {stage0_6[367], stage0_6[368], stage0_6[369], stage0_6[370], stage0_6[371]},
      {stage0_7[312]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[62],stage1_8[111],stage1_7[119],stage1_6[150]}
   );
   gpc615_5 gpc286 (
      {stage0_6[372], stage0_6[373], stage0_6[374], stage0_6[375], stage0_6[376]},
      {stage0_7[313]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[63],stage1_8[112],stage1_7[120],stage1_6[151]}
   );
   gpc615_5 gpc287 (
      {stage0_6[377], stage0_6[378], stage0_6[379], stage0_6[380], stage0_6[381]},
      {stage0_7[314]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[64],stage1_8[113],stage1_7[121],stage1_6[152]}
   );
   gpc615_5 gpc288 (
      {stage0_6[382], stage0_6[383], stage0_6[384], stage0_6[385], stage0_6[386]},
      {stage0_7[315]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[65],stage1_8[114],stage1_7[122],stage1_6[153]}
   );
   gpc615_5 gpc289 (
      {stage0_6[387], stage0_6[388], stage0_6[389], stage0_6[390], stage0_6[391]},
      {stage0_7[316]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[66],stage1_8[115],stage1_7[123],stage1_6[154]}
   );
   gpc615_5 gpc290 (
      {stage0_6[392], stage0_6[393], stage0_6[394], stage0_6[395], stage0_6[396]},
      {stage0_7[317]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[67],stage1_8[116],stage1_7[124],stage1_6[155]}
   );
   gpc615_5 gpc291 (
      {stage0_6[397], stage0_6[398], stage0_6[399], stage0_6[400], stage0_6[401]},
      {stage0_7[318]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[68],stage1_8[117],stage1_7[125],stage1_6[156]}
   );
   gpc615_5 gpc292 (
      {stage0_6[402], stage0_6[403], stage0_6[404], stage0_6[405], stage0_6[406]},
      {stage0_7[319]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[69],stage1_8[118],stage1_7[126],stage1_6[157]}
   );
   gpc615_5 gpc293 (
      {stage0_6[407], stage0_6[408], stage0_6[409], stage0_6[410], stage0_6[411]},
      {stage0_7[320]},
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage1_10[20],stage1_9[70],stage1_8[119],stage1_7[127],stage1_6[158]}
   );
   gpc615_5 gpc294 (
      {stage0_6[412], stage0_6[413], stage0_6[414], stage0_6[415], stage0_6[416]},
      {stage0_7[321]},
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage1_10[21],stage1_9[71],stage1_8[120],stage1_7[128],stage1_6[159]}
   );
   gpc615_5 gpc295 (
      {stage0_6[417], stage0_6[418], stage0_6[419], stage0_6[420], stage0_6[421]},
      {stage0_7[322]},
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage1_10[22],stage1_9[72],stage1_8[121],stage1_7[129],stage1_6[160]}
   );
   gpc615_5 gpc296 (
      {stage0_6[422], stage0_6[423], stage0_6[424], stage0_6[425], stage0_6[426]},
      {stage0_7[323]},
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage1_10[23],stage1_9[73],stage1_8[122],stage1_7[130],stage1_6[161]}
   );
   gpc615_5 gpc297 (
      {stage0_6[427], stage0_6[428], stage0_6[429], stage0_6[430], stage0_6[431]},
      {stage0_7[324]},
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage1_10[24],stage1_9[74],stage1_8[123],stage1_7[131],stage1_6[162]}
   );
   gpc615_5 gpc298 (
      {stage0_6[432], stage0_6[433], stage0_6[434], stage0_6[435], stage0_6[436]},
      {stage0_7[325]},
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage1_10[25],stage1_9[75],stage1_8[124],stage1_7[132],stage1_6[163]}
   );
   gpc615_5 gpc299 (
      {stage0_6[437], stage0_6[438], stage0_6[439], stage0_6[440], stage0_6[441]},
      {stage0_7[326]},
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage1_10[26],stage1_9[76],stage1_8[125],stage1_7[133],stage1_6[164]}
   );
   gpc615_5 gpc300 (
      {stage0_6[442], stage0_6[443], stage0_6[444], stage0_6[445], stage0_6[446]},
      {stage0_7[327]},
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage1_10[27],stage1_9[77],stage1_8[126],stage1_7[134],stage1_6[165]}
   );
   gpc615_5 gpc301 (
      {stage0_6[447], stage0_6[448], stage0_6[449], stage0_6[450], stage0_6[451]},
      {stage0_7[328]},
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage1_10[28],stage1_9[78],stage1_8[127],stage1_7[135],stage1_6[166]}
   );
   gpc615_5 gpc302 (
      {stage0_6[452], stage0_6[453], stage0_6[454], stage0_6[455], stage0_6[456]},
      {stage0_7[329]},
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage1_10[29],stage1_9[79],stage1_8[128],stage1_7[136],stage1_6[167]}
   );
   gpc615_5 gpc303 (
      {stage0_7[330], stage0_7[331], stage0_7[332], stage0_7[333], stage0_7[334]},
      {stage0_8[180]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[30],stage1_9[80],stage1_8[129],stage1_7[137]}
   );
   gpc615_5 gpc304 (
      {stage0_7[335], stage0_7[336], stage0_7[337], stage0_7[338], stage0_7[339]},
      {stage0_8[181]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[31],stage1_9[81],stage1_8[130],stage1_7[138]}
   );
   gpc615_5 gpc305 (
      {stage0_7[340], stage0_7[341], stage0_7[342], stage0_7[343], stage0_7[344]},
      {stage0_8[182]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[32],stage1_9[82],stage1_8[131],stage1_7[139]}
   );
   gpc615_5 gpc306 (
      {stage0_7[345], stage0_7[346], stage0_7[347], stage0_7[348], stage0_7[349]},
      {stage0_8[183]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[33],stage1_9[83],stage1_8[132],stage1_7[140]}
   );
   gpc615_5 gpc307 (
      {stage0_7[350], stage0_7[351], stage0_7[352], stage0_7[353], stage0_7[354]},
      {stage0_8[184]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[34],stage1_9[84],stage1_8[133],stage1_7[141]}
   );
   gpc615_5 gpc308 (
      {stage0_7[355], stage0_7[356], stage0_7[357], stage0_7[358], stage0_7[359]},
      {stage0_8[185]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[35],stage1_9[85],stage1_8[134],stage1_7[142]}
   );
   gpc615_5 gpc309 (
      {stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364]},
      {stage0_8[186]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[36],stage1_9[86],stage1_8[135],stage1_7[143]}
   );
   gpc615_5 gpc310 (
      {stage0_7[365], stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369]},
      {stage0_8[187]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[37],stage1_9[87],stage1_8[136],stage1_7[144]}
   );
   gpc615_5 gpc311 (
      {stage0_7[370], stage0_7[371], stage0_7[372], stage0_7[373], stage0_7[374]},
      {stage0_8[188]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[38],stage1_9[88],stage1_8[137],stage1_7[145]}
   );
   gpc615_5 gpc312 (
      {stage0_7[375], stage0_7[376], stage0_7[377], stage0_7[378], stage0_7[379]},
      {stage0_8[189]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[39],stage1_9[89],stage1_8[138],stage1_7[146]}
   );
   gpc615_5 gpc313 (
      {stage0_7[380], stage0_7[381], stage0_7[382], stage0_7[383], stage0_7[384]},
      {stage0_8[190]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[40],stage1_9[90],stage1_8[139],stage1_7[147]}
   );
   gpc615_5 gpc314 (
      {stage0_7[385], stage0_7[386], stage0_7[387], stage0_7[388], stage0_7[389]},
      {stage0_8[191]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[41],stage1_9[91],stage1_8[140],stage1_7[148]}
   );
   gpc615_5 gpc315 (
      {stage0_7[390], stage0_7[391], stage0_7[392], stage0_7[393], stage0_7[394]},
      {stage0_8[192]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[42],stage1_9[92],stage1_8[141],stage1_7[149]}
   );
   gpc615_5 gpc316 (
      {stage0_7[395], stage0_7[396], stage0_7[397], stage0_7[398], stage0_7[399]},
      {stage0_8[193]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[43],stage1_9[93],stage1_8[142],stage1_7[150]}
   );
   gpc615_5 gpc317 (
      {stage0_7[400], stage0_7[401], stage0_7[402], stage0_7[403], stage0_7[404]},
      {stage0_8[194]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[44],stage1_9[94],stage1_8[143],stage1_7[151]}
   );
   gpc615_5 gpc318 (
      {stage0_7[405], stage0_7[406], stage0_7[407], stage0_7[408], stage0_7[409]},
      {stage0_8[195]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[45],stage1_9[95],stage1_8[144],stage1_7[152]}
   );
   gpc615_5 gpc319 (
      {stage0_7[410], stage0_7[411], stage0_7[412], stage0_7[413], stage0_7[414]},
      {stage0_8[196]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[46],stage1_9[96],stage1_8[145],stage1_7[153]}
   );
   gpc615_5 gpc320 (
      {stage0_7[415], stage0_7[416], stage0_7[417], stage0_7[418], stage0_7[419]},
      {stage0_8[197]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[47],stage1_9[97],stage1_8[146],stage1_7[154]}
   );
   gpc615_5 gpc321 (
      {stage0_7[420], stage0_7[421], stage0_7[422], stage0_7[423], stage0_7[424]},
      {stage0_8[198]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[48],stage1_9[98],stage1_8[147],stage1_7[155]}
   );
   gpc606_5 gpc322 (
      {stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[19],stage1_10[49],stage1_9[99],stage1_8[148]}
   );
   gpc606_5 gpc323 (
      {stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209], stage0_8[210]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[20],stage1_10[50],stage1_9[100],stage1_8[149]}
   );
   gpc606_5 gpc324 (
      {stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[21],stage1_10[51],stage1_9[101],stage1_8[150]}
   );
   gpc606_5 gpc325 (
      {stage0_8[217], stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[22],stage1_10[52],stage1_9[102],stage1_8[151]}
   );
   gpc606_5 gpc326 (
      {stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[23],stage1_10[53],stage1_9[103],stage1_8[152]}
   );
   gpc606_5 gpc327 (
      {stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[24],stage1_10[54],stage1_9[104],stage1_8[153]}
   );
   gpc606_5 gpc328 (
      {stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239], stage0_8[240]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[25],stage1_10[55],stage1_9[105],stage1_8[154]}
   );
   gpc606_5 gpc329 (
      {stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245], stage0_8[246]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[26],stage1_10[56],stage1_9[106],stage1_8[155]}
   );
   gpc606_5 gpc330 (
      {stage0_8[247], stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251], stage0_8[252]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[27],stage1_10[57],stage1_9[107],stage1_8[156]}
   );
   gpc606_5 gpc331 (
      {stage0_8[253], stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257], stage0_8[258]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[28],stage1_10[58],stage1_9[108],stage1_8[157]}
   );
   gpc606_5 gpc332 (
      {stage0_8[259], stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[29],stage1_10[59],stage1_9[109],stage1_8[158]}
   );
   gpc606_5 gpc333 (
      {stage0_8[265], stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[30],stage1_10[60],stage1_9[110],stage1_8[159]}
   );
   gpc606_5 gpc334 (
      {stage0_8[271], stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[31],stage1_10[61],stage1_9[111],stage1_8[160]}
   );
   gpc606_5 gpc335 (
      {stage0_8[277], stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[32],stage1_10[62],stage1_9[112],stage1_8[161]}
   );
   gpc606_5 gpc336 (
      {stage0_8[283], stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[33],stage1_10[63],stage1_9[113],stage1_8[162]}
   );
   gpc606_5 gpc337 (
      {stage0_8[289], stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[34],stage1_10[64],stage1_9[114],stage1_8[163]}
   );
   gpc606_5 gpc338 (
      {stage0_8[295], stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[35],stage1_10[65],stage1_9[115],stage1_8[164]}
   );
   gpc606_5 gpc339 (
      {stage0_8[301], stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[36],stage1_10[66],stage1_9[116],stage1_8[165]}
   );
   gpc606_5 gpc340 (
      {stage0_8[307], stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[37],stage1_10[67],stage1_9[117],stage1_8[166]}
   );
   gpc606_5 gpc341 (
      {stage0_8[313], stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[38],stage1_10[68],stage1_9[118],stage1_8[167]}
   );
   gpc606_5 gpc342 (
      {stage0_8[319], stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[39],stage1_10[69],stage1_9[119],stage1_8[168]}
   );
   gpc606_5 gpc343 (
      {stage0_8[325], stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[40],stage1_10[70],stage1_9[120],stage1_8[169]}
   );
   gpc606_5 gpc344 (
      {stage0_8[331], stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[41],stage1_10[71],stage1_9[121],stage1_8[170]}
   );
   gpc606_5 gpc345 (
      {stage0_8[337], stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341], stage0_8[342]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[42],stage1_10[72],stage1_9[122],stage1_8[171]}
   );
   gpc606_5 gpc346 (
      {stage0_8[343], stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347], stage0_8[348]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[43],stage1_10[73],stage1_9[123],stage1_8[172]}
   );
   gpc606_5 gpc347 (
      {stage0_8[349], stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353], stage0_8[354]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[44],stage1_10[74],stage1_9[124],stage1_8[173]}
   );
   gpc606_5 gpc348 (
      {stage0_8[355], stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[45],stage1_10[75],stage1_9[125],stage1_8[174]}
   );
   gpc606_5 gpc349 (
      {stage0_8[361], stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[46],stage1_10[76],stage1_9[126],stage1_8[175]}
   );
   gpc606_5 gpc350 (
      {stage0_8[367], stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371], stage0_8[372]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[47],stage1_10[77],stage1_9[127],stage1_8[176]}
   );
   gpc606_5 gpc351 (
      {stage0_8[373], stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377], stage0_8[378]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[48],stage1_10[78],stage1_9[128],stage1_8[177]}
   );
   gpc606_5 gpc352 (
      {stage0_8[379], stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383], stage0_8[384]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[49],stage1_10[79],stage1_9[129],stage1_8[178]}
   );
   gpc606_5 gpc353 (
      {stage0_8[385], stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389], stage0_8[390]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[50],stage1_10[80],stage1_9[130],stage1_8[179]}
   );
   gpc606_5 gpc354 (
      {stage0_8[391], stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395], stage0_8[396]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[51],stage1_10[81],stage1_9[131],stage1_8[180]}
   );
   gpc606_5 gpc355 (
      {stage0_8[397], stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401], stage0_8[402]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[52],stage1_10[82],stage1_9[132],stage1_8[181]}
   );
   gpc606_5 gpc356 (
      {stage0_8[403], stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407], stage0_8[408]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[53],stage1_10[83],stage1_9[133],stage1_8[182]}
   );
   gpc606_5 gpc357 (
      {stage0_8[409], stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413], stage0_8[414]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[54],stage1_10[84],stage1_9[134],stage1_8[183]}
   );
   gpc606_5 gpc358 (
      {stage0_8[415], stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419], stage0_8[420]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[55],stage1_10[85],stage1_9[135],stage1_8[184]}
   );
   gpc606_5 gpc359 (
      {stage0_8[421], stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425], stage0_8[426]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[56],stage1_10[86],stage1_9[136],stage1_8[185]}
   );
   gpc606_5 gpc360 (
      {stage0_8[427], stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431], stage0_8[432]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[57],stage1_10[87],stage1_9[137],stage1_8[186]}
   );
   gpc606_5 gpc361 (
      {stage0_8[433], stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437], stage0_8[438]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[58],stage1_10[88],stage1_9[138],stage1_8[187]}
   );
   gpc606_5 gpc362 (
      {stage0_8[439], stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443], stage0_8[444]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[59],stage1_10[89],stage1_9[139],stage1_8[188]}
   );
   gpc606_5 gpc363 (
      {stage0_8[445], stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449], stage0_8[450]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[60],stage1_10[90],stage1_9[140],stage1_8[189]}
   );
   gpc606_5 gpc364 (
      {stage0_8[451], stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455], stage0_8[456]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[61],stage1_10[91],stage1_9[141],stage1_8[190]}
   );
   gpc606_5 gpc365 (
      {stage0_8[457], stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461], stage0_8[462]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[62],stage1_10[92],stage1_9[142],stage1_8[191]}
   );
   gpc606_5 gpc366 (
      {stage0_8[463], stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467], stage0_8[468]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[63],stage1_10[93],stage1_9[143],stage1_8[192]}
   );
   gpc606_5 gpc367 (
      {stage0_8[469], stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473], stage0_8[474]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[64],stage1_10[94],stage1_9[144],stage1_8[193]}
   );
   gpc606_5 gpc368 (
      {stage0_8[475], stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479], stage0_8[480]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[65],stage1_10[95],stage1_9[145],stage1_8[194]}
   );
   gpc615_5 gpc369 (
      {stage0_8[481], stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485]},
      {stage0_9[114]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[66],stage1_10[96],stage1_9[146],stage1_8[195]}
   );
   gpc606_5 gpc370 (
      {stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[48],stage1_11[67],stage1_10[97],stage1_9[147]}
   );
   gpc606_5 gpc371 (
      {stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[49],stage1_11[68],stage1_10[98],stage1_9[148]}
   );
   gpc606_5 gpc372 (
      {stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131], stage0_9[132]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[50],stage1_11[69],stage1_10[99],stage1_9[149]}
   );
   gpc606_5 gpc373 (
      {stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137], stage0_9[138]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[51],stage1_11[70],stage1_10[100],stage1_9[150]}
   );
   gpc606_5 gpc374 (
      {stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143], stage0_9[144]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[52],stage1_11[71],stage1_10[101],stage1_9[151]}
   );
   gpc606_5 gpc375 (
      {stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[53],stage1_11[72],stage1_10[102],stage1_9[152]}
   );
   gpc606_5 gpc376 (
      {stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155], stage0_9[156]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[54],stage1_11[73],stage1_10[103],stage1_9[153]}
   );
   gpc606_5 gpc377 (
      {stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161], stage0_9[162]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[55],stage1_11[74],stage1_10[104],stage1_9[154]}
   );
   gpc606_5 gpc378 (
      {stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166], stage0_9[167], stage0_9[168]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[56],stage1_11[75],stage1_10[105],stage1_9[155]}
   );
   gpc606_5 gpc379 (
      {stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[57],stage1_11[76],stage1_10[106],stage1_9[156]}
   );
   gpc606_5 gpc380 (
      {stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[58],stage1_11[77],stage1_10[107],stage1_9[157]}
   );
   gpc606_5 gpc381 (
      {stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185], stage0_9[186]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[59],stage1_11[78],stage1_10[108],stage1_9[158]}
   );
   gpc606_5 gpc382 (
      {stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190], stage0_9[191], stage0_9[192]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[60],stage1_11[79],stage1_10[109],stage1_9[159]}
   );
   gpc606_5 gpc383 (
      {stage0_9[193], stage0_9[194], stage0_9[195], stage0_9[196], stage0_9[197], stage0_9[198]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[61],stage1_11[80],stage1_10[110],stage1_9[160]}
   );
   gpc606_5 gpc384 (
      {stage0_9[199], stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[62],stage1_11[81],stage1_10[111],stage1_9[161]}
   );
   gpc606_5 gpc385 (
      {stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[63],stage1_11[82],stage1_10[112],stage1_9[162]}
   );
   gpc606_5 gpc386 (
      {stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215], stage0_9[216]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[64],stage1_11[83],stage1_10[113],stage1_9[163]}
   );
   gpc606_5 gpc387 (
      {stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220], stage0_9[221], stage0_9[222]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[65],stage1_11[84],stage1_10[114],stage1_9[164]}
   );
   gpc606_5 gpc388 (
      {stage0_9[223], stage0_9[224], stage0_9[225], stage0_9[226], stage0_9[227], stage0_9[228]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[66],stage1_11[85],stage1_10[115],stage1_9[165]}
   );
   gpc606_5 gpc389 (
      {stage0_9[229], stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[67],stage1_11[86],stage1_10[116],stage1_9[166]}
   );
   gpc606_5 gpc390 (
      {stage0_9[235], stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[68],stage1_11[87],stage1_10[117],stage1_9[167]}
   );
   gpc606_5 gpc391 (
      {stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245], stage0_9[246]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[69],stage1_11[88],stage1_10[118],stage1_9[168]}
   );
   gpc606_5 gpc392 (
      {stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250], stage0_9[251], stage0_9[252]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[70],stage1_11[89],stage1_10[119],stage1_9[169]}
   );
   gpc606_5 gpc393 (
      {stage0_9[253], stage0_9[254], stage0_9[255], stage0_9[256], stage0_9[257], stage0_9[258]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[71],stage1_11[90],stage1_10[120],stage1_9[170]}
   );
   gpc606_5 gpc394 (
      {stage0_9[259], stage0_9[260], stage0_9[261], stage0_9[262], stage0_9[263], stage0_9[264]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[72],stage1_11[91],stage1_10[121],stage1_9[171]}
   );
   gpc606_5 gpc395 (
      {stage0_9[265], stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269], stage0_9[270]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[73],stage1_11[92],stage1_10[122],stage1_9[172]}
   );
   gpc606_5 gpc396 (
      {stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275], stage0_9[276]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[74],stage1_11[93],stage1_10[123],stage1_9[173]}
   );
   gpc606_5 gpc397 (
      {stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280], stage0_9[281], stage0_9[282]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[75],stage1_11[94],stage1_10[124],stage1_9[174]}
   );
   gpc606_5 gpc398 (
      {stage0_9[283], stage0_9[284], stage0_9[285], stage0_9[286], stage0_9[287], stage0_9[288]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[76],stage1_11[95],stage1_10[125],stage1_9[175]}
   );
   gpc606_5 gpc399 (
      {stage0_9[289], stage0_9[290], stage0_9[291], stage0_9[292], stage0_9[293], stage0_9[294]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[77],stage1_11[96],stage1_10[126],stage1_9[176]}
   );
   gpc606_5 gpc400 (
      {stage0_9[295], stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299], stage0_9[300]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[78],stage1_11[97],stage1_10[127],stage1_9[177]}
   );
   gpc606_5 gpc401 (
      {stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305], stage0_9[306]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[79],stage1_11[98],stage1_10[128],stage1_9[178]}
   );
   gpc606_5 gpc402 (
      {stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310], stage0_9[311], stage0_9[312]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[80],stage1_11[99],stage1_10[129],stage1_9[179]}
   );
   gpc606_5 gpc403 (
      {stage0_9[313], stage0_9[314], stage0_9[315], stage0_9[316], stage0_9[317], stage0_9[318]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[81],stage1_11[100],stage1_10[130],stage1_9[180]}
   );
   gpc606_5 gpc404 (
      {stage0_9[319], stage0_9[320], stage0_9[321], stage0_9[322], stage0_9[323], stage0_9[324]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[82],stage1_11[101],stage1_10[131],stage1_9[181]}
   );
   gpc606_5 gpc405 (
      {stage0_9[325], stage0_9[326], stage0_9[327], stage0_9[328], stage0_9[329], stage0_9[330]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[83],stage1_11[102],stage1_10[132],stage1_9[182]}
   );
   gpc606_5 gpc406 (
      {stage0_9[331], stage0_9[332], stage0_9[333], stage0_9[334], stage0_9[335], stage0_9[336]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[84],stage1_11[103],stage1_10[133],stage1_9[183]}
   );
   gpc606_5 gpc407 (
      {stage0_9[337], stage0_9[338], stage0_9[339], stage0_9[340], stage0_9[341], stage0_9[342]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[85],stage1_11[104],stage1_10[134],stage1_9[184]}
   );
   gpc606_5 gpc408 (
      {stage0_9[343], stage0_9[344], stage0_9[345], stage0_9[346], stage0_9[347], stage0_9[348]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[86],stage1_11[105],stage1_10[135],stage1_9[185]}
   );
   gpc606_5 gpc409 (
      {stage0_9[349], stage0_9[350], stage0_9[351], stage0_9[352], stage0_9[353], stage0_9[354]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[87],stage1_11[106],stage1_10[136],stage1_9[186]}
   );
   gpc606_5 gpc410 (
      {stage0_9[355], stage0_9[356], stage0_9[357], stage0_9[358], stage0_9[359], stage0_9[360]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[88],stage1_11[107],stage1_10[137],stage1_9[187]}
   );
   gpc606_5 gpc411 (
      {stage0_9[361], stage0_9[362], stage0_9[363], stage0_9[364], stage0_9[365], stage0_9[366]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[89],stage1_11[108],stage1_10[138],stage1_9[188]}
   );
   gpc606_5 gpc412 (
      {stage0_9[367], stage0_9[368], stage0_9[369], stage0_9[370], stage0_9[371], stage0_9[372]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[90],stage1_11[109],stage1_10[139],stage1_9[189]}
   );
   gpc606_5 gpc413 (
      {stage0_9[373], stage0_9[374], stage0_9[375], stage0_9[376], stage0_9[377], stage0_9[378]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[91],stage1_11[110],stage1_10[140],stage1_9[190]}
   );
   gpc606_5 gpc414 (
      {stage0_9[379], stage0_9[380], stage0_9[381], stage0_9[382], stage0_9[383], stage0_9[384]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[92],stage1_11[111],stage1_10[141],stage1_9[191]}
   );
   gpc606_5 gpc415 (
      {stage0_9[385], stage0_9[386], stage0_9[387], stage0_9[388], stage0_9[389], stage0_9[390]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[93],stage1_11[112],stage1_10[142],stage1_9[192]}
   );
   gpc606_5 gpc416 (
      {stage0_9[391], stage0_9[392], stage0_9[393], stage0_9[394], stage0_9[395], stage0_9[396]},
      {stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage1_13[46],stage1_12[94],stage1_11[113],stage1_10[143],stage1_9[193]}
   );
   gpc606_5 gpc417 (
      {stage0_9[397], stage0_9[398], stage0_9[399], stage0_9[400], stage0_9[401], stage0_9[402]},
      {stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage1_13[47],stage1_12[95],stage1_11[114],stage1_10[144],stage1_9[194]}
   );
   gpc606_5 gpc418 (
      {stage0_9[403], stage0_9[404], stage0_9[405], stage0_9[406], stage0_9[407], stage0_9[408]},
      {stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293]},
      {stage1_13[48],stage1_12[96],stage1_11[115],stage1_10[145],stage1_9[195]}
   );
   gpc606_5 gpc419 (
      {stage0_9[409], stage0_9[410], stage0_9[411], stage0_9[412], stage0_9[413], stage0_9[414]},
      {stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage1_13[49],stage1_12[97],stage1_11[116],stage1_10[146],stage1_9[196]}
   );
   gpc606_5 gpc420 (
      {stage0_9[415], stage0_9[416], stage0_9[417], stage0_9[418], stage0_9[419], stage0_9[420]},
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305]},
      {stage1_13[50],stage1_12[98],stage1_11[117],stage1_10[147],stage1_9[197]}
   );
   gpc615_5 gpc421 (
      {stage0_9[421], stage0_9[422], stage0_9[423], stage0_9[424], stage0_9[425]},
      {stage0_10[288]},
      {stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage1_13[51],stage1_12[99],stage1_11[118],stage1_10[148],stage1_9[198]}
   );
   gpc615_5 gpc422 (
      {stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429], stage0_9[430]},
      {stage0_10[289]},
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316], stage0_11[317]},
      {stage1_13[52],stage1_12[100],stage1_11[119],stage1_10[149],stage1_9[199]}
   );
   gpc615_5 gpc423 (
      {stage0_9[431], stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435]},
      {stage0_10[290]},
      {stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323]},
      {stage1_13[53],stage1_12[101],stage1_11[120],stage1_10[150],stage1_9[200]}
   );
   gpc615_5 gpc424 (
      {stage0_9[436], stage0_9[437], stage0_9[438], stage0_9[439], stage0_9[440]},
      {stage0_10[291]},
      {stage0_11[324], stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage1_13[54],stage1_12[102],stage1_11[121],stage1_10[151],stage1_9[201]}
   );
   gpc615_5 gpc425 (
      {stage0_9[441], stage0_9[442], stage0_9[443], stage0_9[444], stage0_9[445]},
      {stage0_10[292]},
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage1_13[55],stage1_12[103],stage1_11[122],stage1_10[152],stage1_9[202]}
   );
   gpc615_5 gpc426 (
      {stage0_9[446], stage0_9[447], stage0_9[448], stage0_9[449], stage0_9[450]},
      {stage0_10[293]},
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage1_13[56],stage1_12[104],stage1_11[123],stage1_10[153],stage1_9[203]}
   );
   gpc615_5 gpc427 (
      {stage0_9[451], stage0_9[452], stage0_9[453], stage0_9[454], stage0_9[455]},
      {stage0_10[294]},
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346], stage0_11[347]},
      {stage1_13[57],stage1_12[105],stage1_11[124],stage1_10[154],stage1_9[204]}
   );
   gpc615_5 gpc428 (
      {stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459], stage0_9[460]},
      {stage0_10[295]},
      {stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353]},
      {stage1_13[58],stage1_12[106],stage1_11[125],stage1_10[155],stage1_9[205]}
   );
   gpc615_5 gpc429 (
      {stage0_9[461], stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465]},
      {stage0_10[296]},
      {stage0_11[354], stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage1_13[59],stage1_12[107],stage1_11[126],stage1_10[156],stage1_9[206]}
   );
   gpc615_5 gpc430 (
      {stage0_9[466], stage0_9[467], stage0_9[468], stage0_9[469], stage0_9[470]},
      {stage0_10[297]},
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage1_13[60],stage1_12[108],stage1_11[127],stage1_10[157],stage1_9[207]}
   );
   gpc615_5 gpc431 (
      {stage0_9[471], stage0_9[472], stage0_9[473], stage0_9[474], stage0_9[475]},
      {stage0_10[298]},
      {stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369], stage0_11[370], stage0_11[371]},
      {stage1_13[61],stage1_12[109],stage1_11[128],stage1_10[158],stage1_9[208]}
   );
   gpc615_5 gpc432 (
      {stage0_9[476], stage0_9[477], stage0_9[478], stage0_9[479], stage0_9[480]},
      {stage0_10[299]},
      {stage0_11[372], stage0_11[373], stage0_11[374], stage0_11[375], stage0_11[376], stage0_11[377]},
      {stage1_13[62],stage1_12[110],stage1_11[129],stage1_10[159],stage1_9[209]}
   );
   gpc615_5 gpc433 (
      {stage0_9[481], stage0_9[482], stage0_9[483], stage0_9[484], stage0_9[485]},
      {stage0_10[300]},
      {stage0_11[378], stage0_11[379], stage0_11[380], stage0_11[381], stage0_11[382], stage0_11[383]},
      {stage1_13[63],stage1_12[111],stage1_11[130],stage1_10[160],stage1_9[210]}
   );
   gpc615_5 gpc434 (
      {stage0_10[301], stage0_10[302], stage0_10[303], stage0_10[304], stage0_10[305]},
      {stage0_11[384]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[64],stage1_12[112],stage1_11[131],stage1_10[161]}
   );
   gpc615_5 gpc435 (
      {stage0_10[306], stage0_10[307], stage0_10[308], stage0_10[309], stage0_10[310]},
      {stage0_11[385]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[65],stage1_12[113],stage1_11[132],stage1_10[162]}
   );
   gpc615_5 gpc436 (
      {stage0_10[311], stage0_10[312], stage0_10[313], stage0_10[314], stage0_10[315]},
      {stage0_11[386]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[66],stage1_12[114],stage1_11[133],stage1_10[163]}
   );
   gpc615_5 gpc437 (
      {stage0_10[316], stage0_10[317], stage0_10[318], stage0_10[319], stage0_10[320]},
      {stage0_11[387]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[67],stage1_12[115],stage1_11[134],stage1_10[164]}
   );
   gpc615_5 gpc438 (
      {stage0_10[321], stage0_10[322], stage0_10[323], stage0_10[324], stage0_10[325]},
      {stage0_11[388]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[68],stage1_12[116],stage1_11[135],stage1_10[165]}
   );
   gpc615_5 gpc439 (
      {stage0_10[326], stage0_10[327], stage0_10[328], stage0_10[329], stage0_10[330]},
      {stage0_11[389]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[69],stage1_12[117],stage1_11[136],stage1_10[166]}
   );
   gpc615_5 gpc440 (
      {stage0_10[331], stage0_10[332], stage0_10[333], stage0_10[334], stage0_10[335]},
      {stage0_11[390]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[70],stage1_12[118],stage1_11[137],stage1_10[167]}
   );
   gpc615_5 gpc441 (
      {stage0_10[336], stage0_10[337], stage0_10[338], stage0_10[339], stage0_10[340]},
      {stage0_11[391]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[71],stage1_12[119],stage1_11[138],stage1_10[168]}
   );
   gpc615_5 gpc442 (
      {stage0_10[341], stage0_10[342], stage0_10[343], stage0_10[344], stage0_10[345]},
      {stage0_11[392]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[72],stage1_12[120],stage1_11[139],stage1_10[169]}
   );
   gpc615_5 gpc443 (
      {stage0_10[346], stage0_10[347], stage0_10[348], stage0_10[349], stage0_10[350]},
      {stage0_11[393]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[73],stage1_12[121],stage1_11[140],stage1_10[170]}
   );
   gpc615_5 gpc444 (
      {stage0_10[351], stage0_10[352], stage0_10[353], stage0_10[354], stage0_10[355]},
      {stage0_11[394]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[74],stage1_12[122],stage1_11[141],stage1_10[171]}
   );
   gpc615_5 gpc445 (
      {stage0_10[356], stage0_10[357], stage0_10[358], stage0_10[359], stage0_10[360]},
      {stage0_11[395]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[75],stage1_12[123],stage1_11[142],stage1_10[172]}
   );
   gpc615_5 gpc446 (
      {stage0_10[361], stage0_10[362], stage0_10[363], stage0_10[364], stage0_10[365]},
      {stage0_11[396]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[76],stage1_12[124],stage1_11[143],stage1_10[173]}
   );
   gpc615_5 gpc447 (
      {stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369], stage0_10[370]},
      {stage0_11[397]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[77],stage1_12[125],stage1_11[144],stage1_10[174]}
   );
   gpc615_5 gpc448 (
      {stage0_10[371], stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375]},
      {stage0_11[398]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[78],stage1_12[126],stage1_11[145],stage1_10[175]}
   );
   gpc615_5 gpc449 (
      {stage0_10[376], stage0_10[377], stage0_10[378], stage0_10[379], stage0_10[380]},
      {stage0_11[399]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[79],stage1_12[127],stage1_11[146],stage1_10[176]}
   );
   gpc2135_5 gpc450 (
      {stage0_11[400], stage0_11[401], stage0_11[402], stage0_11[403], stage0_11[404]},
      {stage0_12[96], stage0_12[97], stage0_12[98]},
      {stage0_13[0]},
      {stage0_14[0], stage0_14[1]},
      {stage1_15[0],stage1_14[16],stage1_13[80],stage1_12[128],stage1_11[147]}
   );
   gpc606_5 gpc451 (
      {stage0_11[405], stage0_11[406], stage0_11[407], stage0_11[408], stage0_11[409], stage0_11[410]},
      {stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5], stage0_13[6]},
      {stage1_15[1],stage1_14[17],stage1_13[81],stage1_12[129],stage1_11[148]}
   );
   gpc606_5 gpc452 (
      {stage0_11[411], stage0_11[412], stage0_11[413], stage0_11[414], stage0_11[415], stage0_11[416]},
      {stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12]},
      {stage1_15[2],stage1_14[18],stage1_13[82],stage1_12[130],stage1_11[149]}
   );
   gpc606_5 gpc453 (
      {stage0_11[417], stage0_11[418], stage0_11[419], stage0_11[420], stage0_11[421], stage0_11[422]},
      {stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17], stage0_13[18]},
      {stage1_15[3],stage1_14[19],stage1_13[83],stage1_12[131],stage1_11[150]}
   );
   gpc606_5 gpc454 (
      {stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103], stage0_12[104]},
      {stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5], stage0_14[6], stage0_14[7]},
      {stage1_16[0],stage1_15[4],stage1_14[20],stage1_13[84],stage1_12[132]}
   );
   gpc606_5 gpc455 (
      {stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109], stage0_12[110]},
      {stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11], stage0_14[12], stage0_14[13]},
      {stage1_16[1],stage1_15[5],stage1_14[21],stage1_13[85],stage1_12[133]}
   );
   gpc606_5 gpc456 (
      {stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115], stage0_12[116]},
      {stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17], stage0_14[18], stage0_14[19]},
      {stage1_16[2],stage1_15[6],stage1_14[22],stage1_13[86],stage1_12[134]}
   );
   gpc606_5 gpc457 (
      {stage0_12[117], stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121], stage0_12[122]},
      {stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23], stage0_14[24], stage0_14[25]},
      {stage1_16[3],stage1_15[7],stage1_14[23],stage1_13[87],stage1_12[135]}
   );
   gpc606_5 gpc458 (
      {stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127], stage0_12[128]},
      {stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29], stage0_14[30], stage0_14[31]},
      {stage1_16[4],stage1_15[8],stage1_14[24],stage1_13[88],stage1_12[136]}
   );
   gpc606_5 gpc459 (
      {stage0_12[129], stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133], stage0_12[134]},
      {stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35], stage0_14[36], stage0_14[37]},
      {stage1_16[5],stage1_15[9],stage1_14[25],stage1_13[89],stage1_12[137]}
   );
   gpc606_5 gpc460 (
      {stage0_12[135], stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139], stage0_12[140]},
      {stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41], stage0_14[42], stage0_14[43]},
      {stage1_16[6],stage1_15[10],stage1_14[26],stage1_13[90],stage1_12[138]}
   );
   gpc606_5 gpc461 (
      {stage0_12[141], stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146]},
      {stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47], stage0_14[48], stage0_14[49]},
      {stage1_16[7],stage1_15[11],stage1_14[27],stage1_13[91],stage1_12[139]}
   );
   gpc606_5 gpc462 (
      {stage0_12[147], stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151], stage0_12[152]},
      {stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53], stage0_14[54], stage0_14[55]},
      {stage1_16[8],stage1_15[12],stage1_14[28],stage1_13[92],stage1_12[140]}
   );
   gpc606_5 gpc463 (
      {stage0_12[153], stage0_12[154], stage0_12[155], stage0_12[156], stage0_12[157], stage0_12[158]},
      {stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59], stage0_14[60], stage0_14[61]},
      {stage1_16[9],stage1_15[13],stage1_14[29],stage1_13[93],stage1_12[141]}
   );
   gpc606_5 gpc464 (
      {stage0_12[159], stage0_12[160], stage0_12[161], stage0_12[162], stage0_12[163], stage0_12[164]},
      {stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65], stage0_14[66], stage0_14[67]},
      {stage1_16[10],stage1_15[14],stage1_14[30],stage1_13[94],stage1_12[142]}
   );
   gpc606_5 gpc465 (
      {stage0_12[165], stage0_12[166], stage0_12[167], stage0_12[168], stage0_12[169], stage0_12[170]},
      {stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71], stage0_14[72], stage0_14[73]},
      {stage1_16[11],stage1_15[15],stage1_14[31],stage1_13[95],stage1_12[143]}
   );
   gpc606_5 gpc466 (
      {stage0_12[171], stage0_12[172], stage0_12[173], stage0_12[174], stage0_12[175], stage0_12[176]},
      {stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77], stage0_14[78], stage0_14[79]},
      {stage1_16[12],stage1_15[16],stage1_14[32],stage1_13[96],stage1_12[144]}
   );
   gpc606_5 gpc467 (
      {stage0_12[177], stage0_12[178], stage0_12[179], stage0_12[180], stage0_12[181], stage0_12[182]},
      {stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83], stage0_14[84], stage0_14[85]},
      {stage1_16[13],stage1_15[17],stage1_14[33],stage1_13[97],stage1_12[145]}
   );
   gpc606_5 gpc468 (
      {stage0_12[183], stage0_12[184], stage0_12[185], stage0_12[186], stage0_12[187], stage0_12[188]},
      {stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89], stage0_14[90], stage0_14[91]},
      {stage1_16[14],stage1_15[18],stage1_14[34],stage1_13[98],stage1_12[146]}
   );
   gpc606_5 gpc469 (
      {stage0_12[189], stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193], stage0_12[194]},
      {stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95], stage0_14[96], stage0_14[97]},
      {stage1_16[15],stage1_15[19],stage1_14[35],stage1_13[99],stage1_12[147]}
   );
   gpc606_5 gpc470 (
      {stage0_12[195], stage0_12[196], stage0_12[197], stage0_12[198], stage0_12[199], stage0_12[200]},
      {stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101], stage0_14[102], stage0_14[103]},
      {stage1_16[16],stage1_15[20],stage1_14[36],stage1_13[100],stage1_12[148]}
   );
   gpc606_5 gpc471 (
      {stage0_12[201], stage0_12[202], stage0_12[203], stage0_12[204], stage0_12[205], stage0_12[206]},
      {stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107], stage0_14[108], stage0_14[109]},
      {stage1_16[17],stage1_15[21],stage1_14[37],stage1_13[101],stage1_12[149]}
   );
   gpc606_5 gpc472 (
      {stage0_12[207], stage0_12[208], stage0_12[209], stage0_12[210], stage0_12[211], stage0_12[212]},
      {stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113], stage0_14[114], stage0_14[115]},
      {stage1_16[18],stage1_15[22],stage1_14[38],stage1_13[102],stage1_12[150]}
   );
   gpc606_5 gpc473 (
      {stage0_12[213], stage0_12[214], stage0_12[215], stage0_12[216], stage0_12[217], stage0_12[218]},
      {stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119], stage0_14[120], stage0_14[121]},
      {stage1_16[19],stage1_15[23],stage1_14[39],stage1_13[103],stage1_12[151]}
   );
   gpc606_5 gpc474 (
      {stage0_12[219], stage0_12[220], stage0_12[221], stage0_12[222], stage0_12[223], stage0_12[224]},
      {stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125], stage0_14[126], stage0_14[127]},
      {stage1_16[20],stage1_15[24],stage1_14[40],stage1_13[104],stage1_12[152]}
   );
   gpc606_5 gpc475 (
      {stage0_12[225], stage0_12[226], stage0_12[227], stage0_12[228], stage0_12[229], stage0_12[230]},
      {stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132], stage0_14[133]},
      {stage1_16[21],stage1_15[25],stage1_14[41],stage1_13[105],stage1_12[153]}
   );
   gpc606_5 gpc476 (
      {stage0_12[231], stage0_12[232], stage0_12[233], stage0_12[234], stage0_12[235], stage0_12[236]},
      {stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137], stage0_14[138], stage0_14[139]},
      {stage1_16[22],stage1_15[26],stage1_14[42],stage1_13[106],stage1_12[154]}
   );
   gpc606_5 gpc477 (
      {stage0_12[237], stage0_12[238], stage0_12[239], stage0_12[240], stage0_12[241], stage0_12[242]},
      {stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143], stage0_14[144], stage0_14[145]},
      {stage1_16[23],stage1_15[27],stage1_14[43],stage1_13[107],stage1_12[155]}
   );
   gpc606_5 gpc478 (
      {stage0_12[243], stage0_12[244], stage0_12[245], stage0_12[246], stage0_12[247], stage0_12[248]},
      {stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149], stage0_14[150], stage0_14[151]},
      {stage1_16[24],stage1_15[28],stage1_14[44],stage1_13[108],stage1_12[156]}
   );
   gpc606_5 gpc479 (
      {stage0_12[249], stage0_12[250], stage0_12[251], stage0_12[252], stage0_12[253], stage0_12[254]},
      {stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155], stage0_14[156], stage0_14[157]},
      {stage1_16[25],stage1_15[29],stage1_14[45],stage1_13[109],stage1_12[157]}
   );
   gpc606_5 gpc480 (
      {stage0_12[255], stage0_12[256], stage0_12[257], stage0_12[258], stage0_12[259], stage0_12[260]},
      {stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161], stage0_14[162], stage0_14[163]},
      {stage1_16[26],stage1_15[30],stage1_14[46],stage1_13[110],stage1_12[158]}
   );
   gpc606_5 gpc481 (
      {stage0_12[261], stage0_12[262], stage0_12[263], stage0_12[264], stage0_12[265], stage0_12[266]},
      {stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167], stage0_14[168], stage0_14[169]},
      {stage1_16[27],stage1_15[31],stage1_14[47],stage1_13[111],stage1_12[159]}
   );
   gpc606_5 gpc482 (
      {stage0_12[267], stage0_12[268], stage0_12[269], stage0_12[270], stage0_12[271], stage0_12[272]},
      {stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173], stage0_14[174], stage0_14[175]},
      {stage1_16[28],stage1_15[32],stage1_14[48],stage1_13[112],stage1_12[160]}
   );
   gpc606_5 gpc483 (
      {stage0_12[273], stage0_12[274], stage0_12[275], stage0_12[276], stage0_12[277], stage0_12[278]},
      {stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179], stage0_14[180], stage0_14[181]},
      {stage1_16[29],stage1_15[33],stage1_14[49],stage1_13[113],stage1_12[161]}
   );
   gpc606_5 gpc484 (
      {stage0_12[279], stage0_12[280], stage0_12[281], stage0_12[282], stage0_12[283], stage0_12[284]},
      {stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185], stage0_14[186], stage0_14[187]},
      {stage1_16[30],stage1_15[34],stage1_14[50],stage1_13[114],stage1_12[162]}
   );
   gpc606_5 gpc485 (
      {stage0_12[285], stage0_12[286], stage0_12[287], stage0_12[288], stage0_12[289], stage0_12[290]},
      {stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191], stage0_14[192], stage0_14[193]},
      {stage1_16[31],stage1_15[35],stage1_14[51],stage1_13[115],stage1_12[163]}
   );
   gpc606_5 gpc486 (
      {stage0_12[291], stage0_12[292], stage0_12[293], stage0_12[294], stage0_12[295], stage0_12[296]},
      {stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197], stage0_14[198], stage0_14[199]},
      {stage1_16[32],stage1_15[36],stage1_14[52],stage1_13[116],stage1_12[164]}
   );
   gpc606_5 gpc487 (
      {stage0_12[297], stage0_12[298], stage0_12[299], stage0_12[300], stage0_12[301], stage0_12[302]},
      {stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203], stage0_14[204], stage0_14[205]},
      {stage1_16[33],stage1_15[37],stage1_14[53],stage1_13[117],stage1_12[165]}
   );
   gpc606_5 gpc488 (
      {stage0_12[303], stage0_12[304], stage0_12[305], stage0_12[306], stage0_12[307], stage0_12[308]},
      {stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209], stage0_14[210], stage0_14[211]},
      {stage1_16[34],stage1_15[38],stage1_14[54],stage1_13[118],stage1_12[166]}
   );
   gpc606_5 gpc489 (
      {stage0_12[309], stage0_12[310], stage0_12[311], stage0_12[312], stage0_12[313], stage0_12[314]},
      {stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215], stage0_14[216], stage0_14[217]},
      {stage1_16[35],stage1_15[39],stage1_14[55],stage1_13[119],stage1_12[167]}
   );
   gpc606_5 gpc490 (
      {stage0_12[315], stage0_12[316], stage0_12[317], stage0_12[318], stage0_12[319], stage0_12[320]},
      {stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221], stage0_14[222], stage0_14[223]},
      {stage1_16[36],stage1_15[40],stage1_14[56],stage1_13[120],stage1_12[168]}
   );
   gpc615_5 gpc491 (
      {stage0_12[321], stage0_12[322], stage0_12[323], stage0_12[324], stage0_12[325]},
      {stage0_13[19]},
      {stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227], stage0_14[228], stage0_14[229]},
      {stage1_16[37],stage1_15[41],stage1_14[57],stage1_13[121],stage1_12[169]}
   );
   gpc615_5 gpc492 (
      {stage0_12[326], stage0_12[327], stage0_12[328], stage0_12[329], stage0_12[330]},
      {stage0_13[20]},
      {stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233], stage0_14[234], stage0_14[235]},
      {stage1_16[38],stage1_15[42],stage1_14[58],stage1_13[122],stage1_12[170]}
   );
   gpc615_5 gpc493 (
      {stage0_12[331], stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335]},
      {stage0_13[21]},
      {stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239], stage0_14[240], stage0_14[241]},
      {stage1_16[39],stage1_15[43],stage1_14[59],stage1_13[123],stage1_12[171]}
   );
   gpc615_5 gpc494 (
      {stage0_12[336], stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340]},
      {stage0_13[22]},
      {stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245], stage0_14[246], stage0_14[247]},
      {stage1_16[40],stage1_15[44],stage1_14[60],stage1_13[124],stage1_12[172]}
   );
   gpc615_5 gpc495 (
      {stage0_12[341], stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345]},
      {stage0_13[23]},
      {stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251], stage0_14[252], stage0_14[253]},
      {stage1_16[41],stage1_15[45],stage1_14[61],stage1_13[125],stage1_12[173]}
   );
   gpc615_5 gpc496 (
      {stage0_12[346], stage0_12[347], stage0_12[348], stage0_12[349], stage0_12[350]},
      {stage0_13[24]},
      {stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257], stage0_14[258], stage0_14[259]},
      {stage1_16[42],stage1_15[46],stage1_14[62],stage1_13[126],stage1_12[174]}
   );
   gpc615_5 gpc497 (
      {stage0_12[351], stage0_12[352], stage0_12[353], stage0_12[354], stage0_12[355]},
      {stage0_13[25]},
      {stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263], stage0_14[264], stage0_14[265]},
      {stage1_16[43],stage1_15[47],stage1_14[63],stage1_13[127],stage1_12[175]}
   );
   gpc615_5 gpc498 (
      {stage0_12[356], stage0_12[357], stage0_12[358], stage0_12[359], stage0_12[360]},
      {stage0_13[26]},
      {stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269], stage0_14[270], stage0_14[271]},
      {stage1_16[44],stage1_15[48],stage1_14[64],stage1_13[128],stage1_12[176]}
   );
   gpc615_5 gpc499 (
      {stage0_12[361], stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365]},
      {stage0_13[27]},
      {stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275], stage0_14[276], stage0_14[277]},
      {stage1_16[45],stage1_15[49],stage1_14[65],stage1_13[129],stage1_12[177]}
   );
   gpc615_5 gpc500 (
      {stage0_12[366], stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370]},
      {stage0_13[28]},
      {stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281], stage0_14[282], stage0_14[283]},
      {stage1_16[46],stage1_15[50],stage1_14[66],stage1_13[130],stage1_12[178]}
   );
   gpc615_5 gpc501 (
      {stage0_12[371], stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375]},
      {stage0_13[29]},
      {stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287], stage0_14[288], stage0_14[289]},
      {stage1_16[47],stage1_15[51],stage1_14[67],stage1_13[131],stage1_12[179]}
   );
   gpc615_5 gpc502 (
      {stage0_12[376], stage0_12[377], stage0_12[378], stage0_12[379], stage0_12[380]},
      {stage0_13[30]},
      {stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293], stage0_14[294], stage0_14[295]},
      {stage1_16[48],stage1_15[52],stage1_14[68],stage1_13[132],stage1_12[180]}
   );
   gpc615_5 gpc503 (
      {stage0_12[381], stage0_12[382], stage0_12[383], stage0_12[384], stage0_12[385]},
      {stage0_13[31]},
      {stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299], stage0_14[300], stage0_14[301]},
      {stage1_16[49],stage1_15[53],stage1_14[69],stage1_13[133],stage1_12[181]}
   );
   gpc615_5 gpc504 (
      {stage0_12[386], stage0_12[387], stage0_12[388], stage0_12[389], stage0_12[390]},
      {stage0_13[32]},
      {stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305], stage0_14[306], stage0_14[307]},
      {stage1_16[50],stage1_15[54],stage1_14[70],stage1_13[134],stage1_12[182]}
   );
   gpc615_5 gpc505 (
      {stage0_12[391], stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395]},
      {stage0_13[33]},
      {stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311], stage0_14[312], stage0_14[313]},
      {stage1_16[51],stage1_15[55],stage1_14[71],stage1_13[135],stage1_12[183]}
   );
   gpc615_5 gpc506 (
      {stage0_12[396], stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400]},
      {stage0_13[34]},
      {stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317], stage0_14[318], stage0_14[319]},
      {stage1_16[52],stage1_15[56],stage1_14[72],stage1_13[136],stage1_12[184]}
   );
   gpc615_5 gpc507 (
      {stage0_12[401], stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405]},
      {stage0_13[35]},
      {stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323], stage0_14[324], stage0_14[325]},
      {stage1_16[53],stage1_15[57],stage1_14[73],stage1_13[137],stage1_12[185]}
   );
   gpc615_5 gpc508 (
      {stage0_12[406], stage0_12[407], stage0_12[408], stage0_12[409], stage0_12[410]},
      {stage0_13[36]},
      {stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329], stage0_14[330], stage0_14[331]},
      {stage1_16[54],stage1_15[58],stage1_14[74],stage1_13[138],stage1_12[186]}
   );
   gpc615_5 gpc509 (
      {stage0_12[411], stage0_12[412], stage0_12[413], stage0_12[414], stage0_12[415]},
      {stage0_13[37]},
      {stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335], stage0_14[336], stage0_14[337]},
      {stage1_16[55],stage1_15[59],stage1_14[75],stage1_13[139],stage1_12[187]}
   );
   gpc615_5 gpc510 (
      {stage0_12[416], stage0_12[417], stage0_12[418], stage0_12[419], stage0_12[420]},
      {stage0_13[38]},
      {stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341], stage0_14[342], stage0_14[343]},
      {stage1_16[56],stage1_15[60],stage1_14[76],stage1_13[140],stage1_12[188]}
   );
   gpc615_5 gpc511 (
      {stage0_12[421], stage0_12[422], stage0_12[423], stage0_12[424], stage0_12[425]},
      {stage0_13[39]},
      {stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347], stage0_14[348], stage0_14[349]},
      {stage1_16[57],stage1_15[61],stage1_14[77],stage1_13[141],stage1_12[189]}
   );
   gpc615_5 gpc512 (
      {stage0_12[426], stage0_12[427], stage0_12[428], stage0_12[429], stage0_12[430]},
      {stage0_13[40]},
      {stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353], stage0_14[354], stage0_14[355]},
      {stage1_16[58],stage1_15[62],stage1_14[78],stage1_13[142],stage1_12[190]}
   );
   gpc615_5 gpc513 (
      {stage0_12[431], stage0_12[432], stage0_12[433], stage0_12[434], stage0_12[435]},
      {stage0_13[41]},
      {stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359], stage0_14[360], stage0_14[361]},
      {stage1_16[59],stage1_15[63],stage1_14[79],stage1_13[143],stage1_12[191]}
   );
   gpc615_5 gpc514 (
      {stage0_12[436], stage0_12[437], stage0_12[438], stage0_12[439], stage0_12[440]},
      {stage0_13[42]},
      {stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365], stage0_14[366], stage0_14[367]},
      {stage1_16[60],stage1_15[64],stage1_14[80],stage1_13[144],stage1_12[192]}
   );
   gpc615_5 gpc515 (
      {stage0_12[441], stage0_12[442], stage0_12[443], stage0_12[444], stage0_12[445]},
      {stage0_13[43]},
      {stage0_14[368], stage0_14[369], stage0_14[370], stage0_14[371], stage0_14[372], stage0_14[373]},
      {stage1_16[61],stage1_15[65],stage1_14[81],stage1_13[145],stage1_12[193]}
   );
   gpc615_5 gpc516 (
      {stage0_12[446], stage0_12[447], stage0_12[448], stage0_12[449], stage0_12[450]},
      {stage0_13[44]},
      {stage0_14[374], stage0_14[375], stage0_14[376], stage0_14[377], stage0_14[378], stage0_14[379]},
      {stage1_16[62],stage1_15[66],stage1_14[82],stage1_13[146],stage1_12[194]}
   );
   gpc615_5 gpc517 (
      {stage0_12[451], stage0_12[452], stage0_12[453], stage0_12[454], stage0_12[455]},
      {stage0_13[45]},
      {stage0_14[380], stage0_14[381], stage0_14[382], stage0_14[383], stage0_14[384], stage0_14[385]},
      {stage1_16[63],stage1_15[67],stage1_14[83],stage1_13[147],stage1_12[195]}
   );
   gpc615_5 gpc518 (
      {stage0_12[456], stage0_12[457], stage0_12[458], stage0_12[459], stage0_12[460]},
      {stage0_13[46]},
      {stage0_14[386], stage0_14[387], stage0_14[388], stage0_14[389], stage0_14[390], stage0_14[391]},
      {stage1_16[64],stage1_15[68],stage1_14[84],stage1_13[148],stage1_12[196]}
   );
   gpc615_5 gpc519 (
      {stage0_12[461], stage0_12[462], stage0_12[463], stage0_12[464], stage0_12[465]},
      {stage0_13[47]},
      {stage0_14[392], stage0_14[393], stage0_14[394], stage0_14[395], stage0_14[396], stage0_14[397]},
      {stage1_16[65],stage1_15[69],stage1_14[85],stage1_13[149],stage1_12[197]}
   );
   gpc615_5 gpc520 (
      {stage0_12[466], stage0_12[467], stage0_12[468], stage0_12[469], stage0_12[470]},
      {stage0_13[48]},
      {stage0_14[398], stage0_14[399], stage0_14[400], stage0_14[401], stage0_14[402], stage0_14[403]},
      {stage1_16[66],stage1_15[70],stage1_14[86],stage1_13[150],stage1_12[198]}
   );
   gpc615_5 gpc521 (
      {stage0_12[471], stage0_12[472], stage0_12[473], stage0_12[474], stage0_12[475]},
      {stage0_13[49]},
      {stage0_14[404], stage0_14[405], stage0_14[406], stage0_14[407], stage0_14[408], stage0_14[409]},
      {stage1_16[67],stage1_15[71],stage1_14[87],stage1_13[151],stage1_12[199]}
   );
   gpc615_5 gpc522 (
      {stage0_12[476], stage0_12[477], stage0_12[478], stage0_12[479], stage0_12[480]},
      {stage0_13[50]},
      {stage0_14[410], stage0_14[411], stage0_14[412], stage0_14[413], stage0_14[414], stage0_14[415]},
      {stage1_16[68],stage1_15[72],stage1_14[88],stage1_13[152],stage1_12[200]}
   );
   gpc615_5 gpc523 (
      {stage0_12[481], stage0_12[482], stage0_12[483], stage0_12[484], stage0_12[485]},
      {stage0_13[51]},
      {stage0_14[416], stage0_14[417], stage0_14[418], stage0_14[419], stage0_14[420], stage0_14[421]},
      {stage1_16[69],stage1_15[73],stage1_14[89],stage1_13[153],stage1_12[201]}
   );
   gpc606_5 gpc524 (
      {stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[70],stage1_15[74],stage1_14[90],stage1_13[154]}
   );
   gpc606_5 gpc525 (
      {stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[71],stage1_15[75],stage1_14[91],stage1_13[155]}
   );
   gpc606_5 gpc526 (
      {stage0_13[64], stage0_13[65], stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[72],stage1_15[76],stage1_14[92],stage1_13[156]}
   );
   gpc606_5 gpc527 (
      {stage0_13[70], stage0_13[71], stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[73],stage1_15[77],stage1_14[93],stage1_13[157]}
   );
   gpc606_5 gpc528 (
      {stage0_13[76], stage0_13[77], stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[74],stage1_15[78],stage1_14[94],stage1_13[158]}
   );
   gpc606_5 gpc529 (
      {stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[75],stage1_15[79],stage1_14[95],stage1_13[159]}
   );
   gpc606_5 gpc530 (
      {stage0_13[88], stage0_13[89], stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[76],stage1_15[80],stage1_14[96],stage1_13[160]}
   );
   gpc606_5 gpc531 (
      {stage0_13[94], stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[77],stage1_15[81],stage1_14[97],stage1_13[161]}
   );
   gpc606_5 gpc532 (
      {stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[78],stage1_15[82],stage1_14[98],stage1_13[162]}
   );
   gpc606_5 gpc533 (
      {stage0_13[106], stage0_13[107], stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[79],stage1_15[83],stage1_14[99],stage1_13[163]}
   );
   gpc606_5 gpc534 (
      {stage0_13[112], stage0_13[113], stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[80],stage1_15[84],stage1_14[100],stage1_13[164]}
   );
   gpc606_5 gpc535 (
      {stage0_13[118], stage0_13[119], stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[81],stage1_15[85],stage1_14[101],stage1_13[165]}
   );
   gpc606_5 gpc536 (
      {stage0_13[124], stage0_13[125], stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[82],stage1_15[86],stage1_14[102],stage1_13[166]}
   );
   gpc606_5 gpc537 (
      {stage0_13[130], stage0_13[131], stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[83],stage1_15[87],stage1_14[103],stage1_13[167]}
   );
   gpc606_5 gpc538 (
      {stage0_13[136], stage0_13[137], stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[84],stage1_15[88],stage1_14[104],stage1_13[168]}
   );
   gpc606_5 gpc539 (
      {stage0_13[142], stage0_13[143], stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[85],stage1_15[89],stage1_14[105],stage1_13[169]}
   );
   gpc606_5 gpc540 (
      {stage0_13[148], stage0_13[149], stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[86],stage1_15[90],stage1_14[106],stage1_13[170]}
   );
   gpc606_5 gpc541 (
      {stage0_13[154], stage0_13[155], stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[87],stage1_15[91],stage1_14[107],stage1_13[171]}
   );
   gpc606_5 gpc542 (
      {stage0_13[160], stage0_13[161], stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[88],stage1_15[92],stage1_14[108],stage1_13[172]}
   );
   gpc606_5 gpc543 (
      {stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169], stage0_13[170], stage0_13[171]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[89],stage1_15[93],stage1_14[109],stage1_13[173]}
   );
   gpc606_5 gpc544 (
      {stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175], stage0_13[176], stage0_13[177]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[90],stage1_15[94],stage1_14[110],stage1_13[174]}
   );
   gpc606_5 gpc545 (
      {stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181], stage0_13[182], stage0_13[183]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[91],stage1_15[95],stage1_14[111],stage1_13[175]}
   );
   gpc606_5 gpc546 (
      {stage0_13[184], stage0_13[185], stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[92],stage1_15[96],stage1_14[112],stage1_13[176]}
   );
   gpc606_5 gpc547 (
      {stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[93],stage1_15[97],stage1_14[113],stage1_13[177]}
   );
   gpc606_5 gpc548 (
      {stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200], stage0_13[201]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[94],stage1_15[98],stage1_14[114],stage1_13[178]}
   );
   gpc606_5 gpc549 (
      {stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205], stage0_13[206], stage0_13[207]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[95],stage1_15[99],stage1_14[115],stage1_13[179]}
   );
   gpc606_5 gpc550 (
      {stage0_13[208], stage0_13[209], stage0_13[210], stage0_13[211], stage0_13[212], stage0_13[213]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[96],stage1_15[100],stage1_14[116],stage1_13[180]}
   );
   gpc606_5 gpc551 (
      {stage0_13[214], stage0_13[215], stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[97],stage1_15[101],stage1_14[117],stage1_13[181]}
   );
   gpc606_5 gpc552 (
      {stage0_13[220], stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[98],stage1_15[102],stage1_14[118],stage1_13[182]}
   );
   gpc615_5 gpc553 (
      {stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230]},
      {stage0_14[422]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[99],stage1_15[103],stage1_14[119],stage1_13[183]}
   );
   gpc615_5 gpc554 (
      {stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235]},
      {stage0_14[423]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[100],stage1_15[104],stage1_14[120],stage1_13[184]}
   );
   gpc615_5 gpc555 (
      {stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240]},
      {stage0_14[424]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[101],stage1_15[105],stage1_14[121],stage1_13[185]}
   );
   gpc615_5 gpc556 (
      {stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245]},
      {stage0_14[425]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[102],stage1_15[106],stage1_14[122],stage1_13[186]}
   );
   gpc615_5 gpc557 (
      {stage0_13[246], stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250]},
      {stage0_14[426]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[103],stage1_15[107],stage1_14[123],stage1_13[187]}
   );
   gpc615_5 gpc558 (
      {stage0_13[251], stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255]},
      {stage0_14[427]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[104],stage1_15[108],stage1_14[124],stage1_13[188]}
   );
   gpc615_5 gpc559 (
      {stage0_13[256], stage0_13[257], stage0_13[258], stage0_13[259], stage0_13[260]},
      {stage0_14[428]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[105],stage1_15[109],stage1_14[125],stage1_13[189]}
   );
   gpc615_5 gpc560 (
      {stage0_13[261], stage0_13[262], stage0_13[263], stage0_13[264], stage0_13[265]},
      {stage0_14[429]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[106],stage1_15[110],stage1_14[126],stage1_13[190]}
   );
   gpc615_5 gpc561 (
      {stage0_13[266], stage0_13[267], stage0_13[268], stage0_13[269], stage0_13[270]},
      {stage0_14[430]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[107],stage1_15[111],stage1_14[127],stage1_13[191]}
   );
   gpc615_5 gpc562 (
      {stage0_13[271], stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275]},
      {stage0_14[431]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[108],stage1_15[112],stage1_14[128],stage1_13[192]}
   );
   gpc615_5 gpc563 (
      {stage0_13[276], stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280]},
      {stage0_14[432]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[109],stage1_15[113],stage1_14[129],stage1_13[193]}
   );
   gpc615_5 gpc564 (
      {stage0_13[281], stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285]},
      {stage0_14[433]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[110],stage1_15[114],stage1_14[130],stage1_13[194]}
   );
   gpc615_5 gpc565 (
      {stage0_13[286], stage0_13[287], stage0_13[288], stage0_13[289], stage0_13[290]},
      {stage0_14[434]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[111],stage1_15[115],stage1_14[131],stage1_13[195]}
   );
   gpc615_5 gpc566 (
      {stage0_13[291], stage0_13[292], stage0_13[293], stage0_13[294], stage0_13[295]},
      {stage0_14[435]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[112],stage1_15[116],stage1_14[132],stage1_13[196]}
   );
   gpc615_5 gpc567 (
      {stage0_13[296], stage0_13[297], stage0_13[298], stage0_13[299], stage0_13[300]},
      {stage0_14[436]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[113],stage1_15[117],stage1_14[133],stage1_13[197]}
   );
   gpc615_5 gpc568 (
      {stage0_13[301], stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305]},
      {stage0_14[437]},
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268], stage0_15[269]},
      {stage1_17[44],stage1_16[114],stage1_15[118],stage1_14[134],stage1_13[198]}
   );
   gpc615_5 gpc569 (
      {stage0_13[306], stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310]},
      {stage0_14[438]},
      {stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275]},
      {stage1_17[45],stage1_16[115],stage1_15[119],stage1_14[135],stage1_13[199]}
   );
   gpc615_5 gpc570 (
      {stage0_13[311], stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315]},
      {stage0_14[439]},
      {stage0_15[276], stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage1_17[46],stage1_16[116],stage1_15[120],stage1_14[136],stage1_13[200]}
   );
   gpc615_5 gpc571 (
      {stage0_13[316], stage0_13[317], stage0_13[318], stage0_13[319], stage0_13[320]},
      {stage0_14[440]},
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287]},
      {stage1_17[47],stage1_16[117],stage1_15[121],stage1_14[137],stage1_13[201]}
   );
   gpc615_5 gpc572 (
      {stage0_13[321], stage0_13[322], stage0_13[323], stage0_13[324], stage0_13[325]},
      {stage0_14[441]},
      {stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage1_17[48],stage1_16[118],stage1_15[122],stage1_14[138],stage1_13[202]}
   );
   gpc615_5 gpc573 (
      {stage0_13[326], stage0_13[327], stage0_13[328], stage0_13[329], stage0_13[330]},
      {stage0_14[442]},
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298], stage0_15[299]},
      {stage1_17[49],stage1_16[119],stage1_15[123],stage1_14[139],stage1_13[203]}
   );
   gpc615_5 gpc574 (
      {stage0_13[331], stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335]},
      {stage0_14[443]},
      {stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305]},
      {stage1_17[50],stage1_16[120],stage1_15[124],stage1_14[140],stage1_13[204]}
   );
   gpc615_5 gpc575 (
      {stage0_13[336], stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340]},
      {stage0_14[444]},
      {stage0_15[306], stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage1_17[51],stage1_16[121],stage1_15[125],stage1_14[141],stage1_13[205]}
   );
   gpc615_5 gpc576 (
      {stage0_13[341], stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345]},
      {stage0_14[445]},
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317]},
      {stage1_17[52],stage1_16[122],stage1_15[126],stage1_14[142],stage1_13[206]}
   );
   gpc615_5 gpc577 (
      {stage0_13[346], stage0_13[347], stage0_13[348], stage0_13[349], stage0_13[350]},
      {stage0_14[446]},
      {stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage1_17[53],stage1_16[123],stage1_15[127],stage1_14[143],stage1_13[207]}
   );
   gpc615_5 gpc578 (
      {stage0_13[351], stage0_13[352], stage0_13[353], stage0_13[354], stage0_13[355]},
      {stage0_14[447]},
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328], stage0_15[329]},
      {stage1_17[54],stage1_16[124],stage1_15[128],stage1_14[144],stage1_13[208]}
   );
   gpc615_5 gpc579 (
      {stage0_13[356], stage0_13[357], stage0_13[358], stage0_13[359], stage0_13[360]},
      {stage0_14[448]},
      {stage0_15[330], stage0_15[331], stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335]},
      {stage1_17[55],stage1_16[125],stage1_15[129],stage1_14[145],stage1_13[209]}
   );
   gpc615_5 gpc580 (
      {stage0_13[361], stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365]},
      {stage0_14[449]},
      {stage0_15[336], stage0_15[337], stage0_15[338], stage0_15[339], stage0_15[340], stage0_15[341]},
      {stage1_17[56],stage1_16[126],stage1_15[130],stage1_14[146],stage1_13[210]}
   );
   gpc615_5 gpc581 (
      {stage0_13[366], stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370]},
      {stage0_14[450]},
      {stage0_15[342], stage0_15[343], stage0_15[344], stage0_15[345], stage0_15[346], stage0_15[347]},
      {stage1_17[57],stage1_16[127],stage1_15[131],stage1_14[147],stage1_13[211]}
   );
   gpc615_5 gpc582 (
      {stage0_13[371], stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375]},
      {stage0_14[451]},
      {stage0_15[348], stage0_15[349], stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353]},
      {stage1_17[58],stage1_16[128],stage1_15[132],stage1_14[148],stage1_13[212]}
   );
   gpc615_5 gpc583 (
      {stage0_13[376], stage0_13[377], stage0_13[378], stage0_13[379], stage0_13[380]},
      {stage0_14[452]},
      {stage0_15[354], stage0_15[355], stage0_15[356], stage0_15[357], stage0_15[358], stage0_15[359]},
      {stage1_17[59],stage1_16[129],stage1_15[133],stage1_14[149],stage1_13[213]}
   );
   gpc615_5 gpc584 (
      {stage0_13[381], stage0_13[382], stage0_13[383], stage0_13[384], stage0_13[385]},
      {stage0_14[453]},
      {stage0_15[360], stage0_15[361], stage0_15[362], stage0_15[363], stage0_15[364], stage0_15[365]},
      {stage1_17[60],stage1_16[130],stage1_15[134],stage1_14[150],stage1_13[214]}
   );
   gpc615_5 gpc585 (
      {stage0_13[386], stage0_13[387], stage0_13[388], stage0_13[389], stage0_13[390]},
      {stage0_14[454]},
      {stage0_15[366], stage0_15[367], stage0_15[368], stage0_15[369], stage0_15[370], stage0_15[371]},
      {stage1_17[61],stage1_16[131],stage1_15[135],stage1_14[151],stage1_13[215]}
   );
   gpc615_5 gpc586 (
      {stage0_13[391], stage0_13[392], stage0_13[393], stage0_13[394], stage0_13[395]},
      {stage0_14[455]},
      {stage0_15[372], stage0_15[373], stage0_15[374], stage0_15[375], stage0_15[376], stage0_15[377]},
      {stage1_17[62],stage1_16[132],stage1_15[136],stage1_14[152],stage1_13[216]}
   );
   gpc615_5 gpc587 (
      {stage0_13[396], stage0_13[397], stage0_13[398], stage0_13[399], stage0_13[400]},
      {stage0_14[456]},
      {stage0_15[378], stage0_15[379], stage0_15[380], stage0_15[381], stage0_15[382], stage0_15[383]},
      {stage1_17[63],stage1_16[133],stage1_15[137],stage1_14[153],stage1_13[217]}
   );
   gpc615_5 gpc588 (
      {stage0_13[401], stage0_13[402], stage0_13[403], stage0_13[404], stage0_13[405]},
      {stage0_14[457]},
      {stage0_15[384], stage0_15[385], stage0_15[386], stage0_15[387], stage0_15[388], stage0_15[389]},
      {stage1_17[64],stage1_16[134],stage1_15[138],stage1_14[154],stage1_13[218]}
   );
   gpc615_5 gpc589 (
      {stage0_13[406], stage0_13[407], stage0_13[408], stage0_13[409], stage0_13[410]},
      {stage0_14[458]},
      {stage0_15[390], stage0_15[391], stage0_15[392], stage0_15[393], stage0_15[394], stage0_15[395]},
      {stage1_17[65],stage1_16[135],stage1_15[139],stage1_14[155],stage1_13[219]}
   );
   gpc615_5 gpc590 (
      {stage0_13[411], stage0_13[412], stage0_13[413], stage0_13[414], stage0_13[415]},
      {stage0_14[459]},
      {stage0_15[396], stage0_15[397], stage0_15[398], stage0_15[399], stage0_15[400], stage0_15[401]},
      {stage1_17[66],stage1_16[136],stage1_15[140],stage1_14[156],stage1_13[220]}
   );
   gpc615_5 gpc591 (
      {stage0_13[416], stage0_13[417], stage0_13[418], stage0_13[419], stage0_13[420]},
      {stage0_14[460]},
      {stage0_15[402], stage0_15[403], stage0_15[404], stage0_15[405], stage0_15[406], stage0_15[407]},
      {stage1_17[67],stage1_16[137],stage1_15[141],stage1_14[157],stage1_13[221]}
   );
   gpc615_5 gpc592 (
      {stage0_13[421], stage0_13[422], stage0_13[423], stage0_13[424], stage0_13[425]},
      {stage0_14[461]},
      {stage0_15[408], stage0_15[409], stage0_15[410], stage0_15[411], stage0_15[412], stage0_15[413]},
      {stage1_17[68],stage1_16[138],stage1_15[142],stage1_14[158],stage1_13[222]}
   );
   gpc615_5 gpc593 (
      {stage0_13[426], stage0_13[427], stage0_13[428], stage0_13[429], stage0_13[430]},
      {stage0_14[462]},
      {stage0_15[414], stage0_15[415], stage0_15[416], stage0_15[417], stage0_15[418], stage0_15[419]},
      {stage1_17[69],stage1_16[139],stage1_15[143],stage1_14[159],stage1_13[223]}
   );
   gpc615_5 gpc594 (
      {stage0_13[431], stage0_13[432], stage0_13[433], stage0_13[434], stage0_13[435]},
      {stage0_14[463]},
      {stage0_15[420], stage0_15[421], stage0_15[422], stage0_15[423], stage0_15[424], stage0_15[425]},
      {stage1_17[70],stage1_16[140],stage1_15[144],stage1_14[160],stage1_13[224]}
   );
   gpc615_5 gpc595 (
      {stage0_13[436], stage0_13[437], stage0_13[438], stage0_13[439], stage0_13[440]},
      {stage0_14[464]},
      {stage0_15[426], stage0_15[427], stage0_15[428], stage0_15[429], stage0_15[430], stage0_15[431]},
      {stage1_17[71],stage1_16[141],stage1_15[145],stage1_14[161],stage1_13[225]}
   );
   gpc615_5 gpc596 (
      {stage0_13[441], stage0_13[442], stage0_13[443], stage0_13[444], stage0_13[445]},
      {stage0_14[465]},
      {stage0_15[432], stage0_15[433], stage0_15[434], stage0_15[435], stage0_15[436], stage0_15[437]},
      {stage1_17[72],stage1_16[142],stage1_15[146],stage1_14[162],stage1_13[226]}
   );
   gpc615_5 gpc597 (
      {stage0_13[446], stage0_13[447], stage0_13[448], stage0_13[449], stage0_13[450]},
      {stage0_14[466]},
      {stage0_15[438], stage0_15[439], stage0_15[440], stage0_15[441], stage0_15[442], stage0_15[443]},
      {stage1_17[73],stage1_16[143],stage1_15[147],stage1_14[163],stage1_13[227]}
   );
   gpc615_5 gpc598 (
      {stage0_13[451], stage0_13[452], stage0_13[453], stage0_13[454], stage0_13[455]},
      {stage0_14[467]},
      {stage0_15[444], stage0_15[445], stage0_15[446], stage0_15[447], stage0_15[448], stage0_15[449]},
      {stage1_17[74],stage1_16[144],stage1_15[148],stage1_14[164],stage1_13[228]}
   );
   gpc615_5 gpc599 (
      {stage0_13[456], stage0_13[457], stage0_13[458], stage0_13[459], stage0_13[460]},
      {stage0_14[468]},
      {stage0_15[450], stage0_15[451], stage0_15[452], stage0_15[453], stage0_15[454], stage0_15[455]},
      {stage1_17[75],stage1_16[145],stage1_15[149],stage1_14[165],stage1_13[229]}
   );
   gpc615_5 gpc600 (
      {stage0_13[461], stage0_13[462], stage0_13[463], stage0_13[464], stage0_13[465]},
      {stage0_14[469]},
      {stage0_15[456], stage0_15[457], stage0_15[458], stage0_15[459], stage0_15[460], stage0_15[461]},
      {stage1_17[76],stage1_16[146],stage1_15[150],stage1_14[166],stage1_13[230]}
   );
   gpc615_5 gpc601 (
      {stage0_13[466], stage0_13[467], stage0_13[468], stage0_13[469], stage0_13[470]},
      {stage0_14[470]},
      {stage0_15[462], stage0_15[463], stage0_15[464], stage0_15[465], stage0_15[466], stage0_15[467]},
      {stage1_17[77],stage1_16[147],stage1_15[151],stage1_14[167],stage1_13[231]}
   );
   gpc615_5 gpc602 (
      {stage0_13[471], stage0_13[472], stage0_13[473], stage0_13[474], stage0_13[475]},
      {stage0_14[471]},
      {stage0_15[468], stage0_15[469], stage0_15[470], stage0_15[471], stage0_15[472], stage0_15[473]},
      {stage1_17[78],stage1_16[148],stage1_15[152],stage1_14[168],stage1_13[232]}
   );
   gpc615_5 gpc603 (
      {stage0_13[476], stage0_13[477], stage0_13[478], stage0_13[479], stage0_13[480]},
      {stage0_14[472]},
      {stage0_15[474], stage0_15[475], stage0_15[476], stage0_15[477], stage0_15[478], stage0_15[479]},
      {stage1_17[79],stage1_16[149],stage1_15[153],stage1_14[169],stage1_13[233]}
   );
   gpc615_5 gpc604 (
      {stage0_13[481], stage0_13[482], stage0_13[483], stage0_13[484], stage0_13[485]},
      {stage0_14[473]},
      {stage0_15[480], stage0_15[481], stage0_15[482], stage0_15[483], stage0_15[484], stage0_15[485]},
      {stage1_17[80],stage1_16[150],stage1_15[154],stage1_14[170],stage1_13[234]}
   );
   gpc1_1 gpc605 (
      {stage0_0[423]},
      {stage1_0[85]}
   );
   gpc1_1 gpc606 (
      {stage0_0[424]},
      {stage1_0[86]}
   );
   gpc1_1 gpc607 (
      {stage0_0[425]},
      {stage1_0[87]}
   );
   gpc1_1 gpc608 (
      {stage0_0[426]},
      {stage1_0[88]}
   );
   gpc1_1 gpc609 (
      {stage0_0[427]},
      {stage1_0[89]}
   );
   gpc1_1 gpc610 (
      {stage0_0[428]},
      {stage1_0[90]}
   );
   gpc1_1 gpc611 (
      {stage0_0[429]},
      {stage1_0[91]}
   );
   gpc1_1 gpc612 (
      {stage0_0[430]},
      {stage1_0[92]}
   );
   gpc1_1 gpc613 (
      {stage0_0[431]},
      {stage1_0[93]}
   );
   gpc1_1 gpc614 (
      {stage0_0[432]},
      {stage1_0[94]}
   );
   gpc1_1 gpc615 (
      {stage0_0[433]},
      {stage1_0[95]}
   );
   gpc1_1 gpc616 (
      {stage0_0[434]},
      {stage1_0[96]}
   );
   gpc1_1 gpc617 (
      {stage0_0[435]},
      {stage1_0[97]}
   );
   gpc1_1 gpc618 (
      {stage0_0[436]},
      {stage1_0[98]}
   );
   gpc1_1 gpc619 (
      {stage0_0[437]},
      {stage1_0[99]}
   );
   gpc1_1 gpc620 (
      {stage0_0[438]},
      {stage1_0[100]}
   );
   gpc1_1 gpc621 (
      {stage0_0[439]},
      {stage1_0[101]}
   );
   gpc1_1 gpc622 (
      {stage0_0[440]},
      {stage1_0[102]}
   );
   gpc1_1 gpc623 (
      {stage0_0[441]},
      {stage1_0[103]}
   );
   gpc1_1 gpc624 (
      {stage0_0[442]},
      {stage1_0[104]}
   );
   gpc1_1 gpc625 (
      {stage0_0[443]},
      {stage1_0[105]}
   );
   gpc1_1 gpc626 (
      {stage0_0[444]},
      {stage1_0[106]}
   );
   gpc1_1 gpc627 (
      {stage0_0[445]},
      {stage1_0[107]}
   );
   gpc1_1 gpc628 (
      {stage0_0[446]},
      {stage1_0[108]}
   );
   gpc1_1 gpc629 (
      {stage0_0[447]},
      {stage1_0[109]}
   );
   gpc1_1 gpc630 (
      {stage0_0[448]},
      {stage1_0[110]}
   );
   gpc1_1 gpc631 (
      {stage0_0[449]},
      {stage1_0[111]}
   );
   gpc1_1 gpc632 (
      {stage0_0[450]},
      {stage1_0[112]}
   );
   gpc1_1 gpc633 (
      {stage0_0[451]},
      {stage1_0[113]}
   );
   gpc1_1 gpc634 (
      {stage0_0[452]},
      {stage1_0[114]}
   );
   gpc1_1 gpc635 (
      {stage0_0[453]},
      {stage1_0[115]}
   );
   gpc1_1 gpc636 (
      {stage0_0[454]},
      {stage1_0[116]}
   );
   gpc1_1 gpc637 (
      {stage0_0[455]},
      {stage1_0[117]}
   );
   gpc1_1 gpc638 (
      {stage0_0[456]},
      {stage1_0[118]}
   );
   gpc1_1 gpc639 (
      {stage0_0[457]},
      {stage1_0[119]}
   );
   gpc1_1 gpc640 (
      {stage0_0[458]},
      {stage1_0[120]}
   );
   gpc1_1 gpc641 (
      {stage0_0[459]},
      {stage1_0[121]}
   );
   gpc1_1 gpc642 (
      {stage0_0[460]},
      {stage1_0[122]}
   );
   gpc1_1 gpc643 (
      {stage0_0[461]},
      {stage1_0[123]}
   );
   gpc1_1 gpc644 (
      {stage0_0[462]},
      {stage1_0[124]}
   );
   gpc1_1 gpc645 (
      {stage0_0[463]},
      {stage1_0[125]}
   );
   gpc1_1 gpc646 (
      {stage0_0[464]},
      {stage1_0[126]}
   );
   gpc1_1 gpc647 (
      {stage0_0[465]},
      {stage1_0[127]}
   );
   gpc1_1 gpc648 (
      {stage0_0[466]},
      {stage1_0[128]}
   );
   gpc1_1 gpc649 (
      {stage0_0[467]},
      {stage1_0[129]}
   );
   gpc1_1 gpc650 (
      {stage0_0[468]},
      {stage1_0[130]}
   );
   gpc1_1 gpc651 (
      {stage0_0[469]},
      {stage1_0[131]}
   );
   gpc1_1 gpc652 (
      {stage0_0[470]},
      {stage1_0[132]}
   );
   gpc1_1 gpc653 (
      {stage0_0[471]},
      {stage1_0[133]}
   );
   gpc1_1 gpc654 (
      {stage0_0[472]},
      {stage1_0[134]}
   );
   gpc1_1 gpc655 (
      {stage0_0[473]},
      {stage1_0[135]}
   );
   gpc1_1 gpc656 (
      {stage0_0[474]},
      {stage1_0[136]}
   );
   gpc1_1 gpc657 (
      {stage0_0[475]},
      {stage1_0[137]}
   );
   gpc1_1 gpc658 (
      {stage0_0[476]},
      {stage1_0[138]}
   );
   gpc1_1 gpc659 (
      {stage0_0[477]},
      {stage1_0[139]}
   );
   gpc1_1 gpc660 (
      {stage0_0[478]},
      {stage1_0[140]}
   );
   gpc1_1 gpc661 (
      {stage0_0[479]},
      {stage1_0[141]}
   );
   gpc1_1 gpc662 (
      {stage0_0[480]},
      {stage1_0[142]}
   );
   gpc1_1 gpc663 (
      {stage0_0[481]},
      {stage1_0[143]}
   );
   gpc1_1 gpc664 (
      {stage0_0[482]},
      {stage1_0[144]}
   );
   gpc1_1 gpc665 (
      {stage0_0[483]},
      {stage1_0[145]}
   );
   gpc1_1 gpc666 (
      {stage0_0[484]},
      {stage1_0[146]}
   );
   gpc1_1 gpc667 (
      {stage0_0[485]},
      {stage1_0[147]}
   );
   gpc1_1 gpc668 (
      {stage0_2[484]},
      {stage1_2[166]}
   );
   gpc1_1 gpc669 (
      {stage0_2[485]},
      {stage1_2[167]}
   );
   gpc1_1 gpc670 (
      {stage0_3[416]},
      {stage1_3[174]}
   );
   gpc1_1 gpc671 (
      {stage0_3[417]},
      {stage1_3[175]}
   );
   gpc1_1 gpc672 (
      {stage0_3[418]},
      {stage1_3[176]}
   );
   gpc1_1 gpc673 (
      {stage0_3[419]},
      {stage1_3[177]}
   );
   gpc1_1 gpc674 (
      {stage0_3[420]},
      {stage1_3[178]}
   );
   gpc1_1 gpc675 (
      {stage0_3[421]},
      {stage1_3[179]}
   );
   gpc1_1 gpc676 (
      {stage0_3[422]},
      {stage1_3[180]}
   );
   gpc1_1 gpc677 (
      {stage0_3[423]},
      {stage1_3[181]}
   );
   gpc1_1 gpc678 (
      {stage0_3[424]},
      {stage1_3[182]}
   );
   gpc1_1 gpc679 (
      {stage0_3[425]},
      {stage1_3[183]}
   );
   gpc1_1 gpc680 (
      {stage0_3[426]},
      {stage1_3[184]}
   );
   gpc1_1 gpc681 (
      {stage0_3[427]},
      {stage1_3[185]}
   );
   gpc1_1 gpc682 (
      {stage0_3[428]},
      {stage1_3[186]}
   );
   gpc1_1 gpc683 (
      {stage0_3[429]},
      {stage1_3[187]}
   );
   gpc1_1 gpc684 (
      {stage0_3[430]},
      {stage1_3[188]}
   );
   gpc1_1 gpc685 (
      {stage0_3[431]},
      {stage1_3[189]}
   );
   gpc1_1 gpc686 (
      {stage0_3[432]},
      {stage1_3[190]}
   );
   gpc1_1 gpc687 (
      {stage0_3[433]},
      {stage1_3[191]}
   );
   gpc1_1 gpc688 (
      {stage0_3[434]},
      {stage1_3[192]}
   );
   gpc1_1 gpc689 (
      {stage0_3[435]},
      {stage1_3[193]}
   );
   gpc1_1 gpc690 (
      {stage0_3[436]},
      {stage1_3[194]}
   );
   gpc1_1 gpc691 (
      {stage0_3[437]},
      {stage1_3[195]}
   );
   gpc1_1 gpc692 (
      {stage0_3[438]},
      {stage1_3[196]}
   );
   gpc1_1 gpc693 (
      {stage0_3[439]},
      {stage1_3[197]}
   );
   gpc1_1 gpc694 (
      {stage0_3[440]},
      {stage1_3[198]}
   );
   gpc1_1 gpc695 (
      {stage0_3[441]},
      {stage1_3[199]}
   );
   gpc1_1 gpc696 (
      {stage0_3[442]},
      {stage1_3[200]}
   );
   gpc1_1 gpc697 (
      {stage0_3[443]},
      {stage1_3[201]}
   );
   gpc1_1 gpc698 (
      {stage0_3[444]},
      {stage1_3[202]}
   );
   gpc1_1 gpc699 (
      {stage0_3[445]},
      {stage1_3[203]}
   );
   gpc1_1 gpc700 (
      {stage0_3[446]},
      {stage1_3[204]}
   );
   gpc1_1 gpc701 (
      {stage0_3[447]},
      {stage1_3[205]}
   );
   gpc1_1 gpc702 (
      {stage0_3[448]},
      {stage1_3[206]}
   );
   gpc1_1 gpc703 (
      {stage0_3[449]},
      {stage1_3[207]}
   );
   gpc1_1 gpc704 (
      {stage0_3[450]},
      {stage1_3[208]}
   );
   gpc1_1 gpc705 (
      {stage0_3[451]},
      {stage1_3[209]}
   );
   gpc1_1 gpc706 (
      {stage0_3[452]},
      {stage1_3[210]}
   );
   gpc1_1 gpc707 (
      {stage0_3[453]},
      {stage1_3[211]}
   );
   gpc1_1 gpc708 (
      {stage0_3[454]},
      {stage1_3[212]}
   );
   gpc1_1 gpc709 (
      {stage0_3[455]},
      {stage1_3[213]}
   );
   gpc1_1 gpc710 (
      {stage0_3[456]},
      {stage1_3[214]}
   );
   gpc1_1 gpc711 (
      {stage0_3[457]},
      {stage1_3[215]}
   );
   gpc1_1 gpc712 (
      {stage0_3[458]},
      {stage1_3[216]}
   );
   gpc1_1 gpc713 (
      {stage0_3[459]},
      {stage1_3[217]}
   );
   gpc1_1 gpc714 (
      {stage0_3[460]},
      {stage1_3[218]}
   );
   gpc1_1 gpc715 (
      {stage0_3[461]},
      {stage1_3[219]}
   );
   gpc1_1 gpc716 (
      {stage0_3[462]},
      {stage1_3[220]}
   );
   gpc1_1 gpc717 (
      {stage0_3[463]},
      {stage1_3[221]}
   );
   gpc1_1 gpc718 (
      {stage0_3[464]},
      {stage1_3[222]}
   );
   gpc1_1 gpc719 (
      {stage0_3[465]},
      {stage1_3[223]}
   );
   gpc1_1 gpc720 (
      {stage0_3[466]},
      {stage1_3[224]}
   );
   gpc1_1 gpc721 (
      {stage0_3[467]},
      {stage1_3[225]}
   );
   gpc1_1 gpc722 (
      {stage0_3[468]},
      {stage1_3[226]}
   );
   gpc1_1 gpc723 (
      {stage0_3[469]},
      {stage1_3[227]}
   );
   gpc1_1 gpc724 (
      {stage0_3[470]},
      {stage1_3[228]}
   );
   gpc1_1 gpc725 (
      {stage0_3[471]},
      {stage1_3[229]}
   );
   gpc1_1 gpc726 (
      {stage0_3[472]},
      {stage1_3[230]}
   );
   gpc1_1 gpc727 (
      {stage0_3[473]},
      {stage1_3[231]}
   );
   gpc1_1 gpc728 (
      {stage0_3[474]},
      {stage1_3[232]}
   );
   gpc1_1 gpc729 (
      {stage0_3[475]},
      {stage1_3[233]}
   );
   gpc1_1 gpc730 (
      {stage0_3[476]},
      {stage1_3[234]}
   );
   gpc1_1 gpc731 (
      {stage0_3[477]},
      {stage1_3[235]}
   );
   gpc1_1 gpc732 (
      {stage0_3[478]},
      {stage1_3[236]}
   );
   gpc1_1 gpc733 (
      {stage0_3[479]},
      {stage1_3[237]}
   );
   gpc1_1 gpc734 (
      {stage0_3[480]},
      {stage1_3[238]}
   );
   gpc1_1 gpc735 (
      {stage0_3[481]},
      {stage1_3[239]}
   );
   gpc1_1 gpc736 (
      {stage0_3[482]},
      {stage1_3[240]}
   );
   gpc1_1 gpc737 (
      {stage0_3[483]},
      {stage1_3[241]}
   );
   gpc1_1 gpc738 (
      {stage0_3[484]},
      {stage1_3[242]}
   );
   gpc1_1 gpc739 (
      {stage0_3[485]},
      {stage1_3[243]}
   );
   gpc1_1 gpc740 (
      {stage0_5[337]},
      {stage1_5[188]}
   );
   gpc1_1 gpc741 (
      {stage0_5[338]},
      {stage1_5[189]}
   );
   gpc1_1 gpc742 (
      {stage0_5[339]},
      {stage1_5[190]}
   );
   gpc1_1 gpc743 (
      {stage0_5[340]},
      {stage1_5[191]}
   );
   gpc1_1 gpc744 (
      {stage0_5[341]},
      {stage1_5[192]}
   );
   gpc1_1 gpc745 (
      {stage0_5[342]},
      {stage1_5[193]}
   );
   gpc1_1 gpc746 (
      {stage0_5[343]},
      {stage1_5[194]}
   );
   gpc1_1 gpc747 (
      {stage0_5[344]},
      {stage1_5[195]}
   );
   gpc1_1 gpc748 (
      {stage0_5[345]},
      {stage1_5[196]}
   );
   gpc1_1 gpc749 (
      {stage0_5[346]},
      {stage1_5[197]}
   );
   gpc1_1 gpc750 (
      {stage0_5[347]},
      {stage1_5[198]}
   );
   gpc1_1 gpc751 (
      {stage0_5[348]},
      {stage1_5[199]}
   );
   gpc1_1 gpc752 (
      {stage0_5[349]},
      {stage1_5[200]}
   );
   gpc1_1 gpc753 (
      {stage0_5[350]},
      {stage1_5[201]}
   );
   gpc1_1 gpc754 (
      {stage0_5[351]},
      {stage1_5[202]}
   );
   gpc1_1 gpc755 (
      {stage0_5[352]},
      {stage1_5[203]}
   );
   gpc1_1 gpc756 (
      {stage0_5[353]},
      {stage1_5[204]}
   );
   gpc1_1 gpc757 (
      {stage0_5[354]},
      {stage1_5[205]}
   );
   gpc1_1 gpc758 (
      {stage0_5[355]},
      {stage1_5[206]}
   );
   gpc1_1 gpc759 (
      {stage0_5[356]},
      {stage1_5[207]}
   );
   gpc1_1 gpc760 (
      {stage0_5[357]},
      {stage1_5[208]}
   );
   gpc1_1 gpc761 (
      {stage0_5[358]},
      {stage1_5[209]}
   );
   gpc1_1 gpc762 (
      {stage0_5[359]},
      {stage1_5[210]}
   );
   gpc1_1 gpc763 (
      {stage0_5[360]},
      {stage1_5[211]}
   );
   gpc1_1 gpc764 (
      {stage0_5[361]},
      {stage1_5[212]}
   );
   gpc1_1 gpc765 (
      {stage0_5[362]},
      {stage1_5[213]}
   );
   gpc1_1 gpc766 (
      {stage0_5[363]},
      {stage1_5[214]}
   );
   gpc1_1 gpc767 (
      {stage0_5[364]},
      {stage1_5[215]}
   );
   gpc1_1 gpc768 (
      {stage0_5[365]},
      {stage1_5[216]}
   );
   gpc1_1 gpc769 (
      {stage0_5[366]},
      {stage1_5[217]}
   );
   gpc1_1 gpc770 (
      {stage0_5[367]},
      {stage1_5[218]}
   );
   gpc1_1 gpc771 (
      {stage0_5[368]},
      {stage1_5[219]}
   );
   gpc1_1 gpc772 (
      {stage0_5[369]},
      {stage1_5[220]}
   );
   gpc1_1 gpc773 (
      {stage0_5[370]},
      {stage1_5[221]}
   );
   gpc1_1 gpc774 (
      {stage0_5[371]},
      {stage1_5[222]}
   );
   gpc1_1 gpc775 (
      {stage0_5[372]},
      {stage1_5[223]}
   );
   gpc1_1 gpc776 (
      {stage0_5[373]},
      {stage1_5[224]}
   );
   gpc1_1 gpc777 (
      {stage0_5[374]},
      {stage1_5[225]}
   );
   gpc1_1 gpc778 (
      {stage0_5[375]},
      {stage1_5[226]}
   );
   gpc1_1 gpc779 (
      {stage0_5[376]},
      {stage1_5[227]}
   );
   gpc1_1 gpc780 (
      {stage0_5[377]},
      {stage1_5[228]}
   );
   gpc1_1 gpc781 (
      {stage0_5[378]},
      {stage1_5[229]}
   );
   gpc1_1 gpc782 (
      {stage0_5[379]},
      {stage1_5[230]}
   );
   gpc1_1 gpc783 (
      {stage0_5[380]},
      {stage1_5[231]}
   );
   gpc1_1 gpc784 (
      {stage0_5[381]},
      {stage1_5[232]}
   );
   gpc1_1 gpc785 (
      {stage0_5[382]},
      {stage1_5[233]}
   );
   gpc1_1 gpc786 (
      {stage0_5[383]},
      {stage1_5[234]}
   );
   gpc1_1 gpc787 (
      {stage0_5[384]},
      {stage1_5[235]}
   );
   gpc1_1 gpc788 (
      {stage0_5[385]},
      {stage1_5[236]}
   );
   gpc1_1 gpc789 (
      {stage0_5[386]},
      {stage1_5[237]}
   );
   gpc1_1 gpc790 (
      {stage0_5[387]},
      {stage1_5[238]}
   );
   gpc1_1 gpc791 (
      {stage0_5[388]},
      {stage1_5[239]}
   );
   gpc1_1 gpc792 (
      {stage0_5[389]},
      {stage1_5[240]}
   );
   gpc1_1 gpc793 (
      {stage0_5[390]},
      {stage1_5[241]}
   );
   gpc1_1 gpc794 (
      {stage0_5[391]},
      {stage1_5[242]}
   );
   gpc1_1 gpc795 (
      {stage0_5[392]},
      {stage1_5[243]}
   );
   gpc1_1 gpc796 (
      {stage0_5[393]},
      {stage1_5[244]}
   );
   gpc1_1 gpc797 (
      {stage0_5[394]},
      {stage1_5[245]}
   );
   gpc1_1 gpc798 (
      {stage0_5[395]},
      {stage1_5[246]}
   );
   gpc1_1 gpc799 (
      {stage0_5[396]},
      {stage1_5[247]}
   );
   gpc1_1 gpc800 (
      {stage0_5[397]},
      {stage1_5[248]}
   );
   gpc1_1 gpc801 (
      {stage0_5[398]},
      {stage1_5[249]}
   );
   gpc1_1 gpc802 (
      {stage0_5[399]},
      {stage1_5[250]}
   );
   gpc1_1 gpc803 (
      {stage0_5[400]},
      {stage1_5[251]}
   );
   gpc1_1 gpc804 (
      {stage0_5[401]},
      {stage1_5[252]}
   );
   gpc1_1 gpc805 (
      {stage0_5[402]},
      {stage1_5[253]}
   );
   gpc1_1 gpc806 (
      {stage0_5[403]},
      {stage1_5[254]}
   );
   gpc1_1 gpc807 (
      {stage0_5[404]},
      {stage1_5[255]}
   );
   gpc1_1 gpc808 (
      {stage0_5[405]},
      {stage1_5[256]}
   );
   gpc1_1 gpc809 (
      {stage0_5[406]},
      {stage1_5[257]}
   );
   gpc1_1 gpc810 (
      {stage0_5[407]},
      {stage1_5[258]}
   );
   gpc1_1 gpc811 (
      {stage0_5[408]},
      {stage1_5[259]}
   );
   gpc1_1 gpc812 (
      {stage0_5[409]},
      {stage1_5[260]}
   );
   gpc1_1 gpc813 (
      {stage0_5[410]},
      {stage1_5[261]}
   );
   gpc1_1 gpc814 (
      {stage0_5[411]},
      {stage1_5[262]}
   );
   gpc1_1 gpc815 (
      {stage0_5[412]},
      {stage1_5[263]}
   );
   gpc1_1 gpc816 (
      {stage0_5[413]},
      {stage1_5[264]}
   );
   gpc1_1 gpc817 (
      {stage0_5[414]},
      {stage1_5[265]}
   );
   gpc1_1 gpc818 (
      {stage0_5[415]},
      {stage1_5[266]}
   );
   gpc1_1 gpc819 (
      {stage0_5[416]},
      {stage1_5[267]}
   );
   gpc1_1 gpc820 (
      {stage0_5[417]},
      {stage1_5[268]}
   );
   gpc1_1 gpc821 (
      {stage0_5[418]},
      {stage1_5[269]}
   );
   gpc1_1 gpc822 (
      {stage0_5[419]},
      {stage1_5[270]}
   );
   gpc1_1 gpc823 (
      {stage0_5[420]},
      {stage1_5[271]}
   );
   gpc1_1 gpc824 (
      {stage0_5[421]},
      {stage1_5[272]}
   );
   gpc1_1 gpc825 (
      {stage0_5[422]},
      {stage1_5[273]}
   );
   gpc1_1 gpc826 (
      {stage0_5[423]},
      {stage1_5[274]}
   );
   gpc1_1 gpc827 (
      {stage0_5[424]},
      {stage1_5[275]}
   );
   gpc1_1 gpc828 (
      {stage0_5[425]},
      {stage1_5[276]}
   );
   gpc1_1 gpc829 (
      {stage0_5[426]},
      {stage1_5[277]}
   );
   gpc1_1 gpc830 (
      {stage0_5[427]},
      {stage1_5[278]}
   );
   gpc1_1 gpc831 (
      {stage0_5[428]},
      {stage1_5[279]}
   );
   gpc1_1 gpc832 (
      {stage0_5[429]},
      {stage1_5[280]}
   );
   gpc1_1 gpc833 (
      {stage0_5[430]},
      {stage1_5[281]}
   );
   gpc1_1 gpc834 (
      {stage0_5[431]},
      {stage1_5[282]}
   );
   gpc1_1 gpc835 (
      {stage0_5[432]},
      {stage1_5[283]}
   );
   gpc1_1 gpc836 (
      {stage0_5[433]},
      {stage1_5[284]}
   );
   gpc1_1 gpc837 (
      {stage0_5[434]},
      {stage1_5[285]}
   );
   gpc1_1 gpc838 (
      {stage0_5[435]},
      {stage1_5[286]}
   );
   gpc1_1 gpc839 (
      {stage0_5[436]},
      {stage1_5[287]}
   );
   gpc1_1 gpc840 (
      {stage0_5[437]},
      {stage1_5[288]}
   );
   gpc1_1 gpc841 (
      {stage0_5[438]},
      {stage1_5[289]}
   );
   gpc1_1 gpc842 (
      {stage0_5[439]},
      {stage1_5[290]}
   );
   gpc1_1 gpc843 (
      {stage0_5[440]},
      {stage1_5[291]}
   );
   gpc1_1 gpc844 (
      {stage0_5[441]},
      {stage1_5[292]}
   );
   gpc1_1 gpc845 (
      {stage0_5[442]},
      {stage1_5[293]}
   );
   gpc1_1 gpc846 (
      {stage0_5[443]},
      {stage1_5[294]}
   );
   gpc1_1 gpc847 (
      {stage0_5[444]},
      {stage1_5[295]}
   );
   gpc1_1 gpc848 (
      {stage0_5[445]},
      {stage1_5[296]}
   );
   gpc1_1 gpc849 (
      {stage0_5[446]},
      {stage1_5[297]}
   );
   gpc1_1 gpc850 (
      {stage0_5[447]},
      {stage1_5[298]}
   );
   gpc1_1 gpc851 (
      {stage0_5[448]},
      {stage1_5[299]}
   );
   gpc1_1 gpc852 (
      {stage0_5[449]},
      {stage1_5[300]}
   );
   gpc1_1 gpc853 (
      {stage0_5[450]},
      {stage1_5[301]}
   );
   gpc1_1 gpc854 (
      {stage0_5[451]},
      {stage1_5[302]}
   );
   gpc1_1 gpc855 (
      {stage0_5[452]},
      {stage1_5[303]}
   );
   gpc1_1 gpc856 (
      {stage0_5[453]},
      {stage1_5[304]}
   );
   gpc1_1 gpc857 (
      {stage0_5[454]},
      {stage1_5[305]}
   );
   gpc1_1 gpc858 (
      {stage0_5[455]},
      {stage1_5[306]}
   );
   gpc1_1 gpc859 (
      {stage0_5[456]},
      {stage1_5[307]}
   );
   gpc1_1 gpc860 (
      {stage0_5[457]},
      {stage1_5[308]}
   );
   gpc1_1 gpc861 (
      {stage0_5[458]},
      {stage1_5[309]}
   );
   gpc1_1 gpc862 (
      {stage0_5[459]},
      {stage1_5[310]}
   );
   gpc1_1 gpc863 (
      {stage0_5[460]},
      {stage1_5[311]}
   );
   gpc1_1 gpc864 (
      {stage0_5[461]},
      {stage1_5[312]}
   );
   gpc1_1 gpc865 (
      {stage0_5[462]},
      {stage1_5[313]}
   );
   gpc1_1 gpc866 (
      {stage0_5[463]},
      {stage1_5[314]}
   );
   gpc1_1 gpc867 (
      {stage0_5[464]},
      {stage1_5[315]}
   );
   gpc1_1 gpc868 (
      {stage0_5[465]},
      {stage1_5[316]}
   );
   gpc1_1 gpc869 (
      {stage0_5[466]},
      {stage1_5[317]}
   );
   gpc1_1 gpc870 (
      {stage0_5[467]},
      {stage1_5[318]}
   );
   gpc1_1 gpc871 (
      {stage0_5[468]},
      {stage1_5[319]}
   );
   gpc1_1 gpc872 (
      {stage0_5[469]},
      {stage1_5[320]}
   );
   gpc1_1 gpc873 (
      {stage0_5[470]},
      {stage1_5[321]}
   );
   gpc1_1 gpc874 (
      {stage0_5[471]},
      {stage1_5[322]}
   );
   gpc1_1 gpc875 (
      {stage0_5[472]},
      {stage1_5[323]}
   );
   gpc1_1 gpc876 (
      {stage0_5[473]},
      {stage1_5[324]}
   );
   gpc1_1 gpc877 (
      {stage0_5[474]},
      {stage1_5[325]}
   );
   gpc1_1 gpc878 (
      {stage0_5[475]},
      {stage1_5[326]}
   );
   gpc1_1 gpc879 (
      {stage0_5[476]},
      {stage1_5[327]}
   );
   gpc1_1 gpc880 (
      {stage0_5[477]},
      {stage1_5[328]}
   );
   gpc1_1 gpc881 (
      {stage0_5[478]},
      {stage1_5[329]}
   );
   gpc1_1 gpc882 (
      {stage0_5[479]},
      {stage1_5[330]}
   );
   gpc1_1 gpc883 (
      {stage0_5[480]},
      {stage1_5[331]}
   );
   gpc1_1 gpc884 (
      {stage0_5[481]},
      {stage1_5[332]}
   );
   gpc1_1 gpc885 (
      {stage0_5[482]},
      {stage1_5[333]}
   );
   gpc1_1 gpc886 (
      {stage0_5[483]},
      {stage1_5[334]}
   );
   gpc1_1 gpc887 (
      {stage0_5[484]},
      {stage1_5[335]}
   );
   gpc1_1 gpc888 (
      {stage0_5[485]},
      {stage1_5[336]}
   );
   gpc1_1 gpc889 (
      {stage0_6[457]},
      {stage1_6[168]}
   );
   gpc1_1 gpc890 (
      {stage0_6[458]},
      {stage1_6[169]}
   );
   gpc1_1 gpc891 (
      {stage0_6[459]},
      {stage1_6[170]}
   );
   gpc1_1 gpc892 (
      {stage0_6[460]},
      {stage1_6[171]}
   );
   gpc1_1 gpc893 (
      {stage0_6[461]},
      {stage1_6[172]}
   );
   gpc1_1 gpc894 (
      {stage0_6[462]},
      {stage1_6[173]}
   );
   gpc1_1 gpc895 (
      {stage0_6[463]},
      {stage1_6[174]}
   );
   gpc1_1 gpc896 (
      {stage0_6[464]},
      {stage1_6[175]}
   );
   gpc1_1 gpc897 (
      {stage0_6[465]},
      {stage1_6[176]}
   );
   gpc1_1 gpc898 (
      {stage0_6[466]},
      {stage1_6[177]}
   );
   gpc1_1 gpc899 (
      {stage0_6[467]},
      {stage1_6[178]}
   );
   gpc1_1 gpc900 (
      {stage0_6[468]},
      {stage1_6[179]}
   );
   gpc1_1 gpc901 (
      {stage0_6[469]},
      {stage1_6[180]}
   );
   gpc1_1 gpc902 (
      {stage0_6[470]},
      {stage1_6[181]}
   );
   gpc1_1 gpc903 (
      {stage0_6[471]},
      {stage1_6[182]}
   );
   gpc1_1 gpc904 (
      {stage0_6[472]},
      {stage1_6[183]}
   );
   gpc1_1 gpc905 (
      {stage0_6[473]},
      {stage1_6[184]}
   );
   gpc1_1 gpc906 (
      {stage0_6[474]},
      {stage1_6[185]}
   );
   gpc1_1 gpc907 (
      {stage0_6[475]},
      {stage1_6[186]}
   );
   gpc1_1 gpc908 (
      {stage0_6[476]},
      {stage1_6[187]}
   );
   gpc1_1 gpc909 (
      {stage0_6[477]},
      {stage1_6[188]}
   );
   gpc1_1 gpc910 (
      {stage0_6[478]},
      {stage1_6[189]}
   );
   gpc1_1 gpc911 (
      {stage0_6[479]},
      {stage1_6[190]}
   );
   gpc1_1 gpc912 (
      {stage0_6[480]},
      {stage1_6[191]}
   );
   gpc1_1 gpc913 (
      {stage0_6[481]},
      {stage1_6[192]}
   );
   gpc1_1 gpc914 (
      {stage0_6[482]},
      {stage1_6[193]}
   );
   gpc1_1 gpc915 (
      {stage0_6[483]},
      {stage1_6[194]}
   );
   gpc1_1 gpc916 (
      {stage0_6[484]},
      {stage1_6[195]}
   );
   gpc1_1 gpc917 (
      {stage0_6[485]},
      {stage1_6[196]}
   );
   gpc1_1 gpc918 (
      {stage0_7[425]},
      {stage1_7[156]}
   );
   gpc1_1 gpc919 (
      {stage0_7[426]},
      {stage1_7[157]}
   );
   gpc1_1 gpc920 (
      {stage0_7[427]},
      {stage1_7[158]}
   );
   gpc1_1 gpc921 (
      {stage0_7[428]},
      {stage1_7[159]}
   );
   gpc1_1 gpc922 (
      {stage0_7[429]},
      {stage1_7[160]}
   );
   gpc1_1 gpc923 (
      {stage0_7[430]},
      {stage1_7[161]}
   );
   gpc1_1 gpc924 (
      {stage0_7[431]},
      {stage1_7[162]}
   );
   gpc1_1 gpc925 (
      {stage0_7[432]},
      {stage1_7[163]}
   );
   gpc1_1 gpc926 (
      {stage0_7[433]},
      {stage1_7[164]}
   );
   gpc1_1 gpc927 (
      {stage0_7[434]},
      {stage1_7[165]}
   );
   gpc1_1 gpc928 (
      {stage0_7[435]},
      {stage1_7[166]}
   );
   gpc1_1 gpc929 (
      {stage0_7[436]},
      {stage1_7[167]}
   );
   gpc1_1 gpc930 (
      {stage0_7[437]},
      {stage1_7[168]}
   );
   gpc1_1 gpc931 (
      {stage0_7[438]},
      {stage1_7[169]}
   );
   gpc1_1 gpc932 (
      {stage0_7[439]},
      {stage1_7[170]}
   );
   gpc1_1 gpc933 (
      {stage0_7[440]},
      {stage1_7[171]}
   );
   gpc1_1 gpc934 (
      {stage0_7[441]},
      {stage1_7[172]}
   );
   gpc1_1 gpc935 (
      {stage0_7[442]},
      {stage1_7[173]}
   );
   gpc1_1 gpc936 (
      {stage0_7[443]},
      {stage1_7[174]}
   );
   gpc1_1 gpc937 (
      {stage0_7[444]},
      {stage1_7[175]}
   );
   gpc1_1 gpc938 (
      {stage0_7[445]},
      {stage1_7[176]}
   );
   gpc1_1 gpc939 (
      {stage0_7[446]},
      {stage1_7[177]}
   );
   gpc1_1 gpc940 (
      {stage0_7[447]},
      {stage1_7[178]}
   );
   gpc1_1 gpc941 (
      {stage0_7[448]},
      {stage1_7[179]}
   );
   gpc1_1 gpc942 (
      {stage0_7[449]},
      {stage1_7[180]}
   );
   gpc1_1 gpc943 (
      {stage0_7[450]},
      {stage1_7[181]}
   );
   gpc1_1 gpc944 (
      {stage0_7[451]},
      {stage1_7[182]}
   );
   gpc1_1 gpc945 (
      {stage0_7[452]},
      {stage1_7[183]}
   );
   gpc1_1 gpc946 (
      {stage0_7[453]},
      {stage1_7[184]}
   );
   gpc1_1 gpc947 (
      {stage0_7[454]},
      {stage1_7[185]}
   );
   gpc1_1 gpc948 (
      {stage0_7[455]},
      {stage1_7[186]}
   );
   gpc1_1 gpc949 (
      {stage0_7[456]},
      {stage1_7[187]}
   );
   gpc1_1 gpc950 (
      {stage0_7[457]},
      {stage1_7[188]}
   );
   gpc1_1 gpc951 (
      {stage0_7[458]},
      {stage1_7[189]}
   );
   gpc1_1 gpc952 (
      {stage0_7[459]},
      {stage1_7[190]}
   );
   gpc1_1 gpc953 (
      {stage0_7[460]},
      {stage1_7[191]}
   );
   gpc1_1 gpc954 (
      {stage0_7[461]},
      {stage1_7[192]}
   );
   gpc1_1 gpc955 (
      {stage0_7[462]},
      {stage1_7[193]}
   );
   gpc1_1 gpc956 (
      {stage0_7[463]},
      {stage1_7[194]}
   );
   gpc1_1 gpc957 (
      {stage0_7[464]},
      {stage1_7[195]}
   );
   gpc1_1 gpc958 (
      {stage0_7[465]},
      {stage1_7[196]}
   );
   gpc1_1 gpc959 (
      {stage0_7[466]},
      {stage1_7[197]}
   );
   gpc1_1 gpc960 (
      {stage0_7[467]},
      {stage1_7[198]}
   );
   gpc1_1 gpc961 (
      {stage0_7[468]},
      {stage1_7[199]}
   );
   gpc1_1 gpc962 (
      {stage0_7[469]},
      {stage1_7[200]}
   );
   gpc1_1 gpc963 (
      {stage0_7[470]},
      {stage1_7[201]}
   );
   gpc1_1 gpc964 (
      {stage0_7[471]},
      {stage1_7[202]}
   );
   gpc1_1 gpc965 (
      {stage0_7[472]},
      {stage1_7[203]}
   );
   gpc1_1 gpc966 (
      {stage0_7[473]},
      {stage1_7[204]}
   );
   gpc1_1 gpc967 (
      {stage0_7[474]},
      {stage1_7[205]}
   );
   gpc1_1 gpc968 (
      {stage0_7[475]},
      {stage1_7[206]}
   );
   gpc1_1 gpc969 (
      {stage0_7[476]},
      {stage1_7[207]}
   );
   gpc1_1 gpc970 (
      {stage0_7[477]},
      {stage1_7[208]}
   );
   gpc1_1 gpc971 (
      {stage0_7[478]},
      {stage1_7[209]}
   );
   gpc1_1 gpc972 (
      {stage0_7[479]},
      {stage1_7[210]}
   );
   gpc1_1 gpc973 (
      {stage0_7[480]},
      {stage1_7[211]}
   );
   gpc1_1 gpc974 (
      {stage0_7[481]},
      {stage1_7[212]}
   );
   gpc1_1 gpc975 (
      {stage0_7[482]},
      {stage1_7[213]}
   );
   gpc1_1 gpc976 (
      {stage0_7[483]},
      {stage1_7[214]}
   );
   gpc1_1 gpc977 (
      {stage0_7[484]},
      {stage1_7[215]}
   );
   gpc1_1 gpc978 (
      {stage0_7[485]},
      {stage1_7[216]}
   );
   gpc1_1 gpc979 (
      {stage0_10[381]},
      {stage1_10[177]}
   );
   gpc1_1 gpc980 (
      {stage0_10[382]},
      {stage1_10[178]}
   );
   gpc1_1 gpc981 (
      {stage0_10[383]},
      {stage1_10[179]}
   );
   gpc1_1 gpc982 (
      {stage0_10[384]},
      {stage1_10[180]}
   );
   gpc1_1 gpc983 (
      {stage0_10[385]},
      {stage1_10[181]}
   );
   gpc1_1 gpc984 (
      {stage0_10[386]},
      {stage1_10[182]}
   );
   gpc1_1 gpc985 (
      {stage0_10[387]},
      {stage1_10[183]}
   );
   gpc1_1 gpc986 (
      {stage0_10[388]},
      {stage1_10[184]}
   );
   gpc1_1 gpc987 (
      {stage0_10[389]},
      {stage1_10[185]}
   );
   gpc1_1 gpc988 (
      {stage0_10[390]},
      {stage1_10[186]}
   );
   gpc1_1 gpc989 (
      {stage0_10[391]},
      {stage1_10[187]}
   );
   gpc1_1 gpc990 (
      {stage0_10[392]},
      {stage1_10[188]}
   );
   gpc1_1 gpc991 (
      {stage0_10[393]},
      {stage1_10[189]}
   );
   gpc1_1 gpc992 (
      {stage0_10[394]},
      {stage1_10[190]}
   );
   gpc1_1 gpc993 (
      {stage0_10[395]},
      {stage1_10[191]}
   );
   gpc1_1 gpc994 (
      {stage0_10[396]},
      {stage1_10[192]}
   );
   gpc1_1 gpc995 (
      {stage0_10[397]},
      {stage1_10[193]}
   );
   gpc1_1 gpc996 (
      {stage0_10[398]},
      {stage1_10[194]}
   );
   gpc1_1 gpc997 (
      {stage0_10[399]},
      {stage1_10[195]}
   );
   gpc1_1 gpc998 (
      {stage0_10[400]},
      {stage1_10[196]}
   );
   gpc1_1 gpc999 (
      {stage0_10[401]},
      {stage1_10[197]}
   );
   gpc1_1 gpc1000 (
      {stage0_10[402]},
      {stage1_10[198]}
   );
   gpc1_1 gpc1001 (
      {stage0_10[403]},
      {stage1_10[199]}
   );
   gpc1_1 gpc1002 (
      {stage0_10[404]},
      {stage1_10[200]}
   );
   gpc1_1 gpc1003 (
      {stage0_10[405]},
      {stage1_10[201]}
   );
   gpc1_1 gpc1004 (
      {stage0_10[406]},
      {stage1_10[202]}
   );
   gpc1_1 gpc1005 (
      {stage0_10[407]},
      {stage1_10[203]}
   );
   gpc1_1 gpc1006 (
      {stage0_10[408]},
      {stage1_10[204]}
   );
   gpc1_1 gpc1007 (
      {stage0_10[409]},
      {stage1_10[205]}
   );
   gpc1_1 gpc1008 (
      {stage0_10[410]},
      {stage1_10[206]}
   );
   gpc1_1 gpc1009 (
      {stage0_10[411]},
      {stage1_10[207]}
   );
   gpc1_1 gpc1010 (
      {stage0_10[412]},
      {stage1_10[208]}
   );
   gpc1_1 gpc1011 (
      {stage0_10[413]},
      {stage1_10[209]}
   );
   gpc1_1 gpc1012 (
      {stage0_10[414]},
      {stage1_10[210]}
   );
   gpc1_1 gpc1013 (
      {stage0_10[415]},
      {stage1_10[211]}
   );
   gpc1_1 gpc1014 (
      {stage0_10[416]},
      {stage1_10[212]}
   );
   gpc1_1 gpc1015 (
      {stage0_10[417]},
      {stage1_10[213]}
   );
   gpc1_1 gpc1016 (
      {stage0_10[418]},
      {stage1_10[214]}
   );
   gpc1_1 gpc1017 (
      {stage0_10[419]},
      {stage1_10[215]}
   );
   gpc1_1 gpc1018 (
      {stage0_10[420]},
      {stage1_10[216]}
   );
   gpc1_1 gpc1019 (
      {stage0_10[421]},
      {stage1_10[217]}
   );
   gpc1_1 gpc1020 (
      {stage0_10[422]},
      {stage1_10[218]}
   );
   gpc1_1 gpc1021 (
      {stage0_10[423]},
      {stage1_10[219]}
   );
   gpc1_1 gpc1022 (
      {stage0_10[424]},
      {stage1_10[220]}
   );
   gpc1_1 gpc1023 (
      {stage0_10[425]},
      {stage1_10[221]}
   );
   gpc1_1 gpc1024 (
      {stage0_10[426]},
      {stage1_10[222]}
   );
   gpc1_1 gpc1025 (
      {stage0_10[427]},
      {stage1_10[223]}
   );
   gpc1_1 gpc1026 (
      {stage0_10[428]},
      {stage1_10[224]}
   );
   gpc1_1 gpc1027 (
      {stage0_10[429]},
      {stage1_10[225]}
   );
   gpc1_1 gpc1028 (
      {stage0_10[430]},
      {stage1_10[226]}
   );
   gpc1_1 gpc1029 (
      {stage0_10[431]},
      {stage1_10[227]}
   );
   gpc1_1 gpc1030 (
      {stage0_10[432]},
      {stage1_10[228]}
   );
   gpc1_1 gpc1031 (
      {stage0_10[433]},
      {stage1_10[229]}
   );
   gpc1_1 gpc1032 (
      {stage0_10[434]},
      {stage1_10[230]}
   );
   gpc1_1 gpc1033 (
      {stage0_10[435]},
      {stage1_10[231]}
   );
   gpc1_1 gpc1034 (
      {stage0_10[436]},
      {stage1_10[232]}
   );
   gpc1_1 gpc1035 (
      {stage0_10[437]},
      {stage1_10[233]}
   );
   gpc1_1 gpc1036 (
      {stage0_10[438]},
      {stage1_10[234]}
   );
   gpc1_1 gpc1037 (
      {stage0_10[439]},
      {stage1_10[235]}
   );
   gpc1_1 gpc1038 (
      {stage0_10[440]},
      {stage1_10[236]}
   );
   gpc1_1 gpc1039 (
      {stage0_10[441]},
      {stage1_10[237]}
   );
   gpc1_1 gpc1040 (
      {stage0_10[442]},
      {stage1_10[238]}
   );
   gpc1_1 gpc1041 (
      {stage0_10[443]},
      {stage1_10[239]}
   );
   gpc1_1 gpc1042 (
      {stage0_10[444]},
      {stage1_10[240]}
   );
   gpc1_1 gpc1043 (
      {stage0_10[445]},
      {stage1_10[241]}
   );
   gpc1_1 gpc1044 (
      {stage0_10[446]},
      {stage1_10[242]}
   );
   gpc1_1 gpc1045 (
      {stage0_10[447]},
      {stage1_10[243]}
   );
   gpc1_1 gpc1046 (
      {stage0_10[448]},
      {stage1_10[244]}
   );
   gpc1_1 gpc1047 (
      {stage0_10[449]},
      {stage1_10[245]}
   );
   gpc1_1 gpc1048 (
      {stage0_10[450]},
      {stage1_10[246]}
   );
   gpc1_1 gpc1049 (
      {stage0_10[451]},
      {stage1_10[247]}
   );
   gpc1_1 gpc1050 (
      {stage0_10[452]},
      {stage1_10[248]}
   );
   gpc1_1 gpc1051 (
      {stage0_10[453]},
      {stage1_10[249]}
   );
   gpc1_1 gpc1052 (
      {stage0_10[454]},
      {stage1_10[250]}
   );
   gpc1_1 gpc1053 (
      {stage0_10[455]},
      {stage1_10[251]}
   );
   gpc1_1 gpc1054 (
      {stage0_10[456]},
      {stage1_10[252]}
   );
   gpc1_1 gpc1055 (
      {stage0_10[457]},
      {stage1_10[253]}
   );
   gpc1_1 gpc1056 (
      {stage0_10[458]},
      {stage1_10[254]}
   );
   gpc1_1 gpc1057 (
      {stage0_10[459]},
      {stage1_10[255]}
   );
   gpc1_1 gpc1058 (
      {stage0_10[460]},
      {stage1_10[256]}
   );
   gpc1_1 gpc1059 (
      {stage0_10[461]},
      {stage1_10[257]}
   );
   gpc1_1 gpc1060 (
      {stage0_10[462]},
      {stage1_10[258]}
   );
   gpc1_1 gpc1061 (
      {stage0_10[463]},
      {stage1_10[259]}
   );
   gpc1_1 gpc1062 (
      {stage0_10[464]},
      {stage1_10[260]}
   );
   gpc1_1 gpc1063 (
      {stage0_10[465]},
      {stage1_10[261]}
   );
   gpc1_1 gpc1064 (
      {stage0_10[466]},
      {stage1_10[262]}
   );
   gpc1_1 gpc1065 (
      {stage0_10[467]},
      {stage1_10[263]}
   );
   gpc1_1 gpc1066 (
      {stage0_10[468]},
      {stage1_10[264]}
   );
   gpc1_1 gpc1067 (
      {stage0_10[469]},
      {stage1_10[265]}
   );
   gpc1_1 gpc1068 (
      {stage0_10[470]},
      {stage1_10[266]}
   );
   gpc1_1 gpc1069 (
      {stage0_10[471]},
      {stage1_10[267]}
   );
   gpc1_1 gpc1070 (
      {stage0_10[472]},
      {stage1_10[268]}
   );
   gpc1_1 gpc1071 (
      {stage0_10[473]},
      {stage1_10[269]}
   );
   gpc1_1 gpc1072 (
      {stage0_10[474]},
      {stage1_10[270]}
   );
   gpc1_1 gpc1073 (
      {stage0_10[475]},
      {stage1_10[271]}
   );
   gpc1_1 gpc1074 (
      {stage0_10[476]},
      {stage1_10[272]}
   );
   gpc1_1 gpc1075 (
      {stage0_10[477]},
      {stage1_10[273]}
   );
   gpc1_1 gpc1076 (
      {stage0_10[478]},
      {stage1_10[274]}
   );
   gpc1_1 gpc1077 (
      {stage0_10[479]},
      {stage1_10[275]}
   );
   gpc1_1 gpc1078 (
      {stage0_10[480]},
      {stage1_10[276]}
   );
   gpc1_1 gpc1079 (
      {stage0_10[481]},
      {stage1_10[277]}
   );
   gpc1_1 gpc1080 (
      {stage0_10[482]},
      {stage1_10[278]}
   );
   gpc1_1 gpc1081 (
      {stage0_10[483]},
      {stage1_10[279]}
   );
   gpc1_1 gpc1082 (
      {stage0_10[484]},
      {stage1_10[280]}
   );
   gpc1_1 gpc1083 (
      {stage0_10[485]},
      {stage1_10[281]}
   );
   gpc1_1 gpc1084 (
      {stage0_11[423]},
      {stage1_11[151]}
   );
   gpc1_1 gpc1085 (
      {stage0_11[424]},
      {stage1_11[152]}
   );
   gpc1_1 gpc1086 (
      {stage0_11[425]},
      {stage1_11[153]}
   );
   gpc1_1 gpc1087 (
      {stage0_11[426]},
      {stage1_11[154]}
   );
   gpc1_1 gpc1088 (
      {stage0_11[427]},
      {stage1_11[155]}
   );
   gpc1_1 gpc1089 (
      {stage0_11[428]},
      {stage1_11[156]}
   );
   gpc1_1 gpc1090 (
      {stage0_11[429]},
      {stage1_11[157]}
   );
   gpc1_1 gpc1091 (
      {stage0_11[430]},
      {stage1_11[158]}
   );
   gpc1_1 gpc1092 (
      {stage0_11[431]},
      {stage1_11[159]}
   );
   gpc1_1 gpc1093 (
      {stage0_11[432]},
      {stage1_11[160]}
   );
   gpc1_1 gpc1094 (
      {stage0_11[433]},
      {stage1_11[161]}
   );
   gpc1_1 gpc1095 (
      {stage0_11[434]},
      {stage1_11[162]}
   );
   gpc1_1 gpc1096 (
      {stage0_11[435]},
      {stage1_11[163]}
   );
   gpc1_1 gpc1097 (
      {stage0_11[436]},
      {stage1_11[164]}
   );
   gpc1_1 gpc1098 (
      {stage0_11[437]},
      {stage1_11[165]}
   );
   gpc1_1 gpc1099 (
      {stage0_11[438]},
      {stage1_11[166]}
   );
   gpc1_1 gpc1100 (
      {stage0_11[439]},
      {stage1_11[167]}
   );
   gpc1_1 gpc1101 (
      {stage0_11[440]},
      {stage1_11[168]}
   );
   gpc1_1 gpc1102 (
      {stage0_11[441]},
      {stage1_11[169]}
   );
   gpc1_1 gpc1103 (
      {stage0_11[442]},
      {stage1_11[170]}
   );
   gpc1_1 gpc1104 (
      {stage0_11[443]},
      {stage1_11[171]}
   );
   gpc1_1 gpc1105 (
      {stage0_11[444]},
      {stage1_11[172]}
   );
   gpc1_1 gpc1106 (
      {stage0_11[445]},
      {stage1_11[173]}
   );
   gpc1_1 gpc1107 (
      {stage0_11[446]},
      {stage1_11[174]}
   );
   gpc1_1 gpc1108 (
      {stage0_11[447]},
      {stage1_11[175]}
   );
   gpc1_1 gpc1109 (
      {stage0_11[448]},
      {stage1_11[176]}
   );
   gpc1_1 gpc1110 (
      {stage0_11[449]},
      {stage1_11[177]}
   );
   gpc1_1 gpc1111 (
      {stage0_11[450]},
      {stage1_11[178]}
   );
   gpc1_1 gpc1112 (
      {stage0_11[451]},
      {stage1_11[179]}
   );
   gpc1_1 gpc1113 (
      {stage0_11[452]},
      {stage1_11[180]}
   );
   gpc1_1 gpc1114 (
      {stage0_11[453]},
      {stage1_11[181]}
   );
   gpc1_1 gpc1115 (
      {stage0_11[454]},
      {stage1_11[182]}
   );
   gpc1_1 gpc1116 (
      {stage0_11[455]},
      {stage1_11[183]}
   );
   gpc1_1 gpc1117 (
      {stage0_11[456]},
      {stage1_11[184]}
   );
   gpc1_1 gpc1118 (
      {stage0_11[457]},
      {stage1_11[185]}
   );
   gpc1_1 gpc1119 (
      {stage0_11[458]},
      {stage1_11[186]}
   );
   gpc1_1 gpc1120 (
      {stage0_11[459]},
      {stage1_11[187]}
   );
   gpc1_1 gpc1121 (
      {stage0_11[460]},
      {stage1_11[188]}
   );
   gpc1_1 gpc1122 (
      {stage0_11[461]},
      {stage1_11[189]}
   );
   gpc1_1 gpc1123 (
      {stage0_11[462]},
      {stage1_11[190]}
   );
   gpc1_1 gpc1124 (
      {stage0_11[463]},
      {stage1_11[191]}
   );
   gpc1_1 gpc1125 (
      {stage0_11[464]},
      {stage1_11[192]}
   );
   gpc1_1 gpc1126 (
      {stage0_11[465]},
      {stage1_11[193]}
   );
   gpc1_1 gpc1127 (
      {stage0_11[466]},
      {stage1_11[194]}
   );
   gpc1_1 gpc1128 (
      {stage0_11[467]},
      {stage1_11[195]}
   );
   gpc1_1 gpc1129 (
      {stage0_11[468]},
      {stage1_11[196]}
   );
   gpc1_1 gpc1130 (
      {stage0_11[469]},
      {stage1_11[197]}
   );
   gpc1_1 gpc1131 (
      {stage0_11[470]},
      {stage1_11[198]}
   );
   gpc1_1 gpc1132 (
      {stage0_11[471]},
      {stage1_11[199]}
   );
   gpc1_1 gpc1133 (
      {stage0_11[472]},
      {stage1_11[200]}
   );
   gpc1_1 gpc1134 (
      {stage0_11[473]},
      {stage1_11[201]}
   );
   gpc1_1 gpc1135 (
      {stage0_11[474]},
      {stage1_11[202]}
   );
   gpc1_1 gpc1136 (
      {stage0_11[475]},
      {stage1_11[203]}
   );
   gpc1_1 gpc1137 (
      {stage0_11[476]},
      {stage1_11[204]}
   );
   gpc1_1 gpc1138 (
      {stage0_11[477]},
      {stage1_11[205]}
   );
   gpc1_1 gpc1139 (
      {stage0_11[478]},
      {stage1_11[206]}
   );
   gpc1_1 gpc1140 (
      {stage0_11[479]},
      {stage1_11[207]}
   );
   gpc1_1 gpc1141 (
      {stage0_11[480]},
      {stage1_11[208]}
   );
   gpc1_1 gpc1142 (
      {stage0_11[481]},
      {stage1_11[209]}
   );
   gpc1_1 gpc1143 (
      {stage0_11[482]},
      {stage1_11[210]}
   );
   gpc1_1 gpc1144 (
      {stage0_11[483]},
      {stage1_11[211]}
   );
   gpc1_1 gpc1145 (
      {stage0_11[484]},
      {stage1_11[212]}
   );
   gpc1_1 gpc1146 (
      {stage0_11[485]},
      {stage1_11[213]}
   );
   gpc1_1 gpc1147 (
      {stage0_14[474]},
      {stage1_14[171]}
   );
   gpc1_1 gpc1148 (
      {stage0_14[475]},
      {stage1_14[172]}
   );
   gpc1_1 gpc1149 (
      {stage0_14[476]},
      {stage1_14[173]}
   );
   gpc1_1 gpc1150 (
      {stage0_14[477]},
      {stage1_14[174]}
   );
   gpc1_1 gpc1151 (
      {stage0_14[478]},
      {stage1_14[175]}
   );
   gpc1_1 gpc1152 (
      {stage0_14[479]},
      {stage1_14[176]}
   );
   gpc1_1 gpc1153 (
      {stage0_14[480]},
      {stage1_14[177]}
   );
   gpc1_1 gpc1154 (
      {stage0_14[481]},
      {stage1_14[178]}
   );
   gpc1_1 gpc1155 (
      {stage0_14[482]},
      {stage1_14[179]}
   );
   gpc1_1 gpc1156 (
      {stage0_14[483]},
      {stage1_14[180]}
   );
   gpc1_1 gpc1157 (
      {stage0_14[484]},
      {stage1_14[181]}
   );
   gpc1_1 gpc1158 (
      {stage0_14[485]},
      {stage1_14[182]}
   );
   gpc1163_5 gpc1159 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc1160 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc1161 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc1162 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc1163 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc1164 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc1165 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc1166 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc1167 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc1168 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc1169 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc606_5 gpc1170 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc1171 (
      {stage1_0[42], stage1_0[43], stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc1172 (
      {stage1_0[48], stage1_0[49], stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53]},
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc606_5 gpc1173 (
      {stage1_0[54], stage1_0[55], stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc606_5 gpc1174 (
      {stage1_0[60], stage1_0[61], stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65]},
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc606_5 gpc1175 (
      {stage1_0[66], stage1_0[67], stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71]},
      {stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc606_5 gpc1176 (
      {stage1_0[72], stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc606_5 gpc1177 (
      {stage1_0[78], stage1_0[79], stage1_0[80], stage1_0[81], stage1_0[82], stage1_0[83]},
      {stage1_2[58], stage1_2[59], stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc606_5 gpc1178 (
      {stage1_0[84], stage1_0[85], stage1_0[86], stage1_0[87], stage1_0[88], stage1_0[89]},
      {stage1_2[64], stage1_2[65], stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc606_5 gpc1179 (
      {stage1_0[90], stage1_0[91], stage1_0[92], stage1_0[93], stage1_0[94], stage1_0[95]},
      {stage1_2[70], stage1_2[71], stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc1180 (
      {stage1_0[96], stage1_0[97], stage1_0[98], stage1_0[99], stage1_0[100], stage1_0[101]},
      {stage1_2[76], stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc606_5 gpc1181 (
      {stage1_0[102], stage1_0[103], stage1_0[104], stage1_0[105], stage1_0[106], stage1_0[107]},
      {stage1_2[82], stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87]},
      {stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22],stage2_0[22]}
   );
   gpc606_5 gpc1182 (
      {stage1_0[108], stage1_0[109], stage1_0[110], stage1_0[111], stage1_0[112], stage1_0[113]},
      {stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91], stage1_2[92], stage1_2[93]},
      {stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23],stage2_0[23]}
   );
   gpc606_5 gpc1183 (
      {stage1_0[114], stage1_0[115], stage1_0[116], stage1_0[117], stage1_0[118], stage1_0[119]},
      {stage1_2[94], stage1_2[95], stage1_2[96], stage1_2[97], stage1_2[98], stage1_2[99]},
      {stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24],stage2_0[24]}
   );
   gpc606_5 gpc1184 (
      {stage1_0[120], stage1_0[121], stage1_0[122], stage1_0[123], stage1_0[124], stage1_0[125]},
      {stage1_2[100], stage1_2[101], stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105]},
      {stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25],stage2_0[25]}
   );
   gpc606_5 gpc1185 (
      {stage1_0[126], stage1_0[127], stage1_0[128], stage1_0[129], stage1_0[130], stage1_0[131]},
      {stage1_2[106], stage1_2[107], stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111]},
      {stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26],stage2_0[26]}
   );
   gpc606_5 gpc1186 (
      {stage1_0[132], stage1_0[133], stage1_0[134], stage1_0[135], stage1_0[136], stage1_0[137]},
      {stage1_2[112], stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117]},
      {stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27],stage2_0[27]}
   );
   gpc606_5 gpc1187 (
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15]},
      {stage2_5[0],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc1188 (
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage2_5[1],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc1189 (
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage2_5[2],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc1190 (
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage2_5[3],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc1191 (
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39]},
      {stage2_5[4],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc1192 (
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45]},
      {stage2_5[5],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc1193 (
      {stage1_1[96], stage1_1[97], stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101]},
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage2_5[6],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc1194 (
      {stage1_1[102], stage1_1[103], stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107]},
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57]},
      {stage2_5[7],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc615_5 gpc1195 (
      {stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121], stage1_2[122]},
      {stage1_3[58]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[8],stage2_4[36],stage2_3[36],stage2_2[36]}
   );
   gpc615_5 gpc1196 (
      {stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126], stage1_2[127]},
      {stage1_3[59]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[9],stage2_4[37],stage2_3[37],stage2_2[37]}
   );
   gpc615_5 gpc1197 (
      {stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131], stage1_2[132]},
      {stage1_3[60]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[10],stage2_4[38],stage2_3[38],stage2_2[38]}
   );
   gpc615_5 gpc1198 (
      {stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137]},
      {stage1_3[61]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[11],stage2_4[39],stage2_3[39],stage2_2[39]}
   );
   gpc615_5 gpc1199 (
      {stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142]},
      {stage1_3[62]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[12],stage2_4[40],stage2_3[40],stage2_2[40]}
   );
   gpc615_5 gpc1200 (
      {stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146], stage1_2[147]},
      {stage1_3[63]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[13],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc615_5 gpc1201 (
      {stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151], stage1_2[152]},
      {stage1_3[64]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[14],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc615_5 gpc1202 (
      {stage1_2[153], stage1_2[154], stage1_2[155], stage1_2[156], stage1_2[157]},
      {stage1_3[65]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[15],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc1203 (
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_4[48]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[8],stage2_5[16],stage2_4[44],stage2_3[44]}
   );
   gpc615_5 gpc1204 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage1_4[49]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[9],stage2_5[17],stage2_4[45],stage2_3[45]}
   );
   gpc615_5 gpc1205 (
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80]},
      {stage1_4[50]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[10],stage2_5[18],stage2_4[46],stage2_3[46]}
   );
   gpc615_5 gpc1206 (
      {stage1_3[81], stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85]},
      {stage1_4[51]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[11],stage2_5[19],stage2_4[47],stage2_3[47]}
   );
   gpc615_5 gpc1207 (
      {stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90]},
      {stage1_4[52]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[12],stage2_5[20],stage2_4[48],stage2_3[48]}
   );
   gpc615_5 gpc1208 (
      {stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage1_4[53]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[13],stage2_5[21],stage2_4[49],stage2_3[49]}
   );
   gpc615_5 gpc1209 (
      {stage1_3[96], stage1_3[97], stage1_3[98], stage1_3[99], stage1_3[100]},
      {stage1_4[54]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[14],stage2_5[22],stage2_4[50],stage2_3[50]}
   );
   gpc615_5 gpc1210 (
      {stage1_3[101], stage1_3[102], stage1_3[103], stage1_3[104], stage1_3[105]},
      {stage1_4[55]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[15],stage2_5[23],stage2_4[51],stage2_3[51]}
   );
   gpc615_5 gpc1211 (
      {stage1_3[106], stage1_3[107], stage1_3[108], stage1_3[109], stage1_3[110]},
      {stage1_4[56]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[16],stage2_5[24],stage2_4[52],stage2_3[52]}
   );
   gpc615_5 gpc1212 (
      {stage1_3[111], stage1_3[112], stage1_3[113], stage1_3[114], stage1_3[115]},
      {stage1_4[57]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[17],stage2_5[25],stage2_4[53],stage2_3[53]}
   );
   gpc615_5 gpc1213 (
      {stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119], stage1_3[120]},
      {stage1_4[58]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[18],stage2_5[26],stage2_4[54],stage2_3[54]}
   );
   gpc615_5 gpc1214 (
      {stage1_3[121], stage1_3[122], stage1_3[123], stage1_3[124], stage1_3[125]},
      {stage1_4[59]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[19],stage2_5[27],stage2_4[55],stage2_3[55]}
   );
   gpc615_5 gpc1215 (
      {stage1_3[126], stage1_3[127], stage1_3[128], stage1_3[129], stage1_3[130]},
      {stage1_4[60]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[20],stage2_5[28],stage2_4[56],stage2_3[56]}
   );
   gpc615_5 gpc1216 (
      {stage1_3[131], stage1_3[132], stage1_3[133], stage1_3[134], stage1_3[135]},
      {stage1_4[61]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[21],stage2_5[29],stage2_4[57],stage2_3[57]}
   );
   gpc615_5 gpc1217 (
      {stage1_3[136], stage1_3[137], stage1_3[138], stage1_3[139], stage1_3[140]},
      {stage1_4[62]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[22],stage2_5[30],stage2_4[58],stage2_3[58]}
   );
   gpc615_5 gpc1218 (
      {stage1_3[141], stage1_3[142], stage1_3[143], stage1_3[144], stage1_3[145]},
      {stage1_4[63]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[23],stage2_5[31],stage2_4[59],stage2_3[59]}
   );
   gpc615_5 gpc1219 (
      {stage1_3[146], stage1_3[147], stage1_3[148], stage1_3[149], stage1_3[150]},
      {stage1_4[64]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[24],stage2_5[32],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc1220 (
      {stage1_3[151], stage1_3[152], stage1_3[153], stage1_3[154], stage1_3[155]},
      {stage1_4[65]},
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage2_7[17],stage2_6[25],stage2_5[33],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc1221 (
      {stage1_3[156], stage1_3[157], stage1_3[158], stage1_3[159], stage1_3[160]},
      {stage1_4[66]},
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage2_7[18],stage2_6[26],stage2_5[34],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc1222 (
      {stage1_3[161], stage1_3[162], stage1_3[163], stage1_3[164], stage1_3[165]},
      {stage1_4[67]},
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage2_7[19],stage2_6[27],stage2_5[35],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc1223 (
      {stage1_3[166], stage1_3[167], stage1_3[168], stage1_3[169], stage1_3[170]},
      {stage1_4[68]},
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage2_7[20],stage2_6[28],stage2_5[36],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc1224 (
      {stage1_3[171], stage1_3[172], stage1_3[173], stage1_3[174], stage1_3[175]},
      {stage1_4[69]},
      {stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131]},
      {stage2_7[21],stage2_6[29],stage2_5[37],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc1225 (
      {stage1_3[176], stage1_3[177], stage1_3[178], stage1_3[179], stage1_3[180]},
      {stage1_4[70]},
      {stage1_5[132], stage1_5[133], stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137]},
      {stage2_7[22],stage2_6[30],stage2_5[38],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc1226 (
      {stage1_3[181], stage1_3[182], stage1_3[183], stage1_3[184], stage1_3[185]},
      {stage1_4[71]},
      {stage1_5[138], stage1_5[139], stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143]},
      {stage2_7[23],stage2_6[31],stage2_5[39],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc1227 (
      {stage1_3[186], stage1_3[187], stage1_3[188], stage1_3[189], stage1_3[190]},
      {stage1_4[72]},
      {stage1_5[144], stage1_5[145], stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149]},
      {stage2_7[24],stage2_6[32],stage2_5[40],stage2_4[68],stage2_3[68]}
   );
   gpc615_5 gpc1228 (
      {stage1_3[191], stage1_3[192], stage1_3[193], stage1_3[194], stage1_3[195]},
      {stage1_4[73]},
      {stage1_5[150], stage1_5[151], stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155]},
      {stage2_7[25],stage2_6[33],stage2_5[41],stage2_4[69],stage2_3[69]}
   );
   gpc615_5 gpc1229 (
      {stage1_3[196], stage1_3[197], stage1_3[198], stage1_3[199], stage1_3[200]},
      {stage1_4[74]},
      {stage1_5[156], stage1_5[157], stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161]},
      {stage2_7[26],stage2_6[34],stage2_5[42],stage2_4[70],stage2_3[70]}
   );
   gpc615_5 gpc1230 (
      {stage1_3[201], stage1_3[202], stage1_3[203], stage1_3[204], stage1_3[205]},
      {stage1_4[75]},
      {stage1_5[162], stage1_5[163], stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167]},
      {stage2_7[27],stage2_6[35],stage2_5[43],stage2_4[71],stage2_3[71]}
   );
   gpc615_5 gpc1231 (
      {stage1_3[206], stage1_3[207], stage1_3[208], stage1_3[209], stage1_3[210]},
      {stage1_4[76]},
      {stage1_5[168], stage1_5[169], stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173]},
      {stage2_7[28],stage2_6[36],stage2_5[44],stage2_4[72],stage2_3[72]}
   );
   gpc615_5 gpc1232 (
      {stage1_3[211], stage1_3[212], stage1_3[213], stage1_3[214], stage1_3[215]},
      {stage1_4[77]},
      {stage1_5[174], stage1_5[175], stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179]},
      {stage2_7[29],stage2_6[37],stage2_5[45],stage2_4[73],stage2_3[73]}
   );
   gpc615_5 gpc1233 (
      {stage1_3[216], stage1_3[217], stage1_3[218], stage1_3[219], stage1_3[220]},
      {stage1_4[78]},
      {stage1_5[180], stage1_5[181], stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185]},
      {stage2_7[30],stage2_6[38],stage2_5[46],stage2_4[74],stage2_3[74]}
   );
   gpc615_5 gpc1234 (
      {stage1_3[221], stage1_3[222], stage1_3[223], stage1_3[224], stage1_3[225]},
      {stage1_4[79]},
      {stage1_5[186], stage1_5[187], stage1_5[188], stage1_5[189], stage1_5[190], stage1_5[191]},
      {stage2_7[31],stage2_6[39],stage2_5[47],stage2_4[75],stage2_3[75]}
   );
   gpc615_5 gpc1235 (
      {stage1_3[226], stage1_3[227], stage1_3[228], stage1_3[229], stage1_3[230]},
      {stage1_4[80]},
      {stage1_5[192], stage1_5[193], stage1_5[194], stage1_5[195], stage1_5[196], stage1_5[197]},
      {stage2_7[32],stage2_6[40],stage2_5[48],stage2_4[76],stage2_3[76]}
   );
   gpc615_5 gpc1236 (
      {stage1_3[231], stage1_3[232], stage1_3[233], stage1_3[234], stage1_3[235]},
      {stage1_4[81]},
      {stage1_5[198], stage1_5[199], stage1_5[200], stage1_5[201], stage1_5[202], stage1_5[203]},
      {stage2_7[33],stage2_6[41],stage2_5[49],stage2_4[77],stage2_3[77]}
   );
   gpc615_5 gpc1237 (
      {stage1_4[82], stage1_4[83], stage1_4[84], stage1_4[85], stage1_4[86]},
      {stage1_5[204]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[34],stage2_6[42],stage2_5[50],stage2_4[78]}
   );
   gpc615_5 gpc1238 (
      {stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91]},
      {stage1_5[205]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[35],stage2_6[43],stage2_5[51],stage2_4[79]}
   );
   gpc615_5 gpc1239 (
      {stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96]},
      {stage1_5[206]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[36],stage2_6[44],stage2_5[52],stage2_4[80]}
   );
   gpc615_5 gpc1240 (
      {stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage1_5[207]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[37],stage2_6[45],stage2_5[53],stage2_4[81]}
   );
   gpc615_5 gpc1241 (
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106]},
      {stage1_5[208]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[38],stage2_6[46],stage2_5[54],stage2_4[82]}
   );
   gpc615_5 gpc1242 (
      {stage1_4[107], stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111]},
      {stage1_5[209]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[39],stage2_6[47],stage2_5[55],stage2_4[83]}
   );
   gpc615_5 gpc1243 (
      {stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116]},
      {stage1_5[210]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[40],stage2_6[48],stage2_5[56],stage2_4[84]}
   );
   gpc615_5 gpc1244 (
      {stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121]},
      {stage1_5[211]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[41],stage2_6[49],stage2_5[57],stage2_4[85]}
   );
   gpc615_5 gpc1245 (
      {stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125], stage1_4[126]},
      {stage1_5[212]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[42],stage2_6[50],stage2_5[58],stage2_4[86]}
   );
   gpc615_5 gpc1246 (
      {stage1_4[127], stage1_4[128], stage1_4[129], stage1_4[130], stage1_4[131]},
      {stage1_5[213]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[43],stage2_6[51],stage2_5[59],stage2_4[87]}
   );
   gpc615_5 gpc1247 (
      {stage1_4[132], stage1_4[133], stage1_4[134], stage1_4[135], stage1_4[136]},
      {stage1_5[214]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[44],stage2_6[52],stage2_5[60],stage2_4[88]}
   );
   gpc615_5 gpc1248 (
      {stage1_4[137], stage1_4[138], stage1_4[139], stage1_4[140], stage1_4[141]},
      {stage1_5[215]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[45],stage2_6[53],stage2_5[61],stage2_4[89]}
   );
   gpc615_5 gpc1249 (
      {stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145], stage1_4[146]},
      {stage1_5[216]},
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage2_8[12],stage2_7[46],stage2_6[54],stage2_5[62],stage2_4[90]}
   );
   gpc615_5 gpc1250 (
      {stage1_4[147], stage1_4[148], stage1_4[149], stage1_4[150], stage1_4[151]},
      {stage1_5[217]},
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage2_8[13],stage2_7[47],stage2_6[55],stage2_5[63],stage2_4[91]}
   );
   gpc615_5 gpc1251 (
      {stage1_4[152], stage1_4[153], stage1_4[154], stage1_4[155], stage1_4[156]},
      {stage1_5[218]},
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage2_8[14],stage2_7[48],stage2_6[56],stage2_5[64],stage2_4[92]}
   );
   gpc615_5 gpc1252 (
      {stage1_4[157], stage1_4[158], stage1_4[159], stage1_4[160], stage1_4[161]},
      {stage1_5[219]},
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage2_8[15],stage2_7[49],stage2_6[57],stage2_5[65],stage2_4[93]}
   );
   gpc615_5 gpc1253 (
      {stage1_4[162], stage1_4[163], stage1_4[164], stage1_4[165], stage1_4[166]},
      {stage1_5[220]},
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage2_8[16],stage2_7[50],stage2_6[58],stage2_5[66],stage2_4[94]}
   );
   gpc615_5 gpc1254 (
      {stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170], stage1_4[171]},
      {stage1_5[221]},
      {stage1_6[102], stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107]},
      {stage2_8[17],stage2_7[51],stage2_6[59],stage2_5[67],stage2_4[95]}
   );
   gpc615_5 gpc1255 (
      {stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175], stage1_4[176]},
      {stage1_5[222]},
      {stage1_6[108], stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113]},
      {stage2_8[18],stage2_7[52],stage2_6[60],stage2_5[68],stage2_4[96]}
   );
   gpc615_5 gpc1256 (
      {stage1_4[177], stage1_4[178], stage1_4[179], stage1_4[180], stage1_4[181]},
      {stage1_5[223]},
      {stage1_6[114], stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119]},
      {stage2_8[19],stage2_7[53],stage2_6[61],stage2_5[69],stage2_4[97]}
   );
   gpc615_5 gpc1257 (
      {stage1_4[182], stage1_4[183], stage1_4[184], stage1_4[185], stage1_4[186]},
      {stage1_5[224]},
      {stage1_6[120], stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125]},
      {stage2_8[20],stage2_7[54],stage2_6[62],stage2_5[70],stage2_4[98]}
   );
   gpc615_5 gpc1258 (
      {stage1_4[187], stage1_4[188], stage1_4[189], stage1_4[190], stage1_4[191]},
      {stage1_5[225]},
      {stage1_6[126], stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131]},
      {stage2_8[21],stage2_7[55],stage2_6[63],stage2_5[71],stage2_4[99]}
   );
   gpc615_5 gpc1259 (
      {stage1_4[192], stage1_4[193], stage1_4[194], stage1_4[195], stage1_4[196]},
      {stage1_5[226]},
      {stage1_6[132], stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137]},
      {stage2_8[22],stage2_7[56],stage2_6[64],stage2_5[72],stage2_4[100]}
   );
   gpc615_5 gpc1260 (
      {stage1_4[197], stage1_4[198], stage1_4[199], stage1_4[200], stage1_4[201]},
      {stage1_5[227]},
      {stage1_6[138], stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143]},
      {stage2_8[23],stage2_7[57],stage2_6[65],stage2_5[73],stage2_4[101]}
   );
   gpc615_5 gpc1261 (
      {stage1_4[202], stage1_4[203], stage1_4[204], stage1_4[205], stage1_4[206]},
      {stage1_5[228]},
      {stage1_6[144], stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149]},
      {stage2_8[24],stage2_7[58],stage2_6[66],stage2_5[74],stage2_4[102]}
   );
   gpc615_5 gpc1262 (
      {stage1_4[207], stage1_4[208], stage1_4[209], stage1_4[210], stage1_4[211]},
      {stage1_5[229]},
      {stage1_6[150], stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155]},
      {stage2_8[25],stage2_7[59],stage2_6[67],stage2_5[75],stage2_4[103]}
   );
   gpc615_5 gpc1263 (
      {stage1_4[212], stage1_4[213], stage1_4[214], stage1_4[215], stage1_4[216]},
      {stage1_5[230]},
      {stage1_6[156], stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161]},
      {stage2_8[26],stage2_7[60],stage2_6[68],stage2_5[76],stage2_4[104]}
   );
   gpc615_5 gpc1264 (
      {stage1_4[217], stage1_4[218], stage1_4[219], stage1_4[220], stage1_4[221]},
      {stage1_5[231]},
      {stage1_6[162], stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166], stage1_6[167]},
      {stage2_8[27],stage2_7[61],stage2_6[69],stage2_5[77],stage2_4[105]}
   );
   gpc606_5 gpc1265 (
      {stage1_5[232], stage1_5[233], stage1_5[234], stage1_5[235], stage1_5[236], stage1_5[237]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[28],stage2_7[62],stage2_6[70],stage2_5[78]}
   );
   gpc606_5 gpc1266 (
      {stage1_5[238], stage1_5[239], stage1_5[240], stage1_5[241], stage1_5[242], stage1_5[243]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[29],stage2_7[63],stage2_6[71],stage2_5[79]}
   );
   gpc606_5 gpc1267 (
      {stage1_5[244], stage1_5[245], stage1_5[246], stage1_5[247], stage1_5[248], stage1_5[249]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[30],stage2_7[64],stage2_6[72],stage2_5[80]}
   );
   gpc606_5 gpc1268 (
      {stage1_5[250], stage1_5[251], stage1_5[252], stage1_5[253], stage1_5[254], stage1_5[255]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[31],stage2_7[65],stage2_6[73],stage2_5[81]}
   );
   gpc606_5 gpc1269 (
      {stage1_5[256], stage1_5[257], stage1_5[258], stage1_5[259], stage1_5[260], stage1_5[261]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[32],stage2_7[66],stage2_6[74],stage2_5[82]}
   );
   gpc606_5 gpc1270 (
      {stage1_5[262], stage1_5[263], stage1_5[264], stage1_5[265], stage1_5[266], stage1_5[267]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[33],stage2_7[67],stage2_6[75],stage2_5[83]}
   );
   gpc606_5 gpc1271 (
      {stage1_5[268], stage1_5[269], stage1_5[270], stage1_5[271], stage1_5[272], stage1_5[273]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[34],stage2_7[68],stage2_6[76],stage2_5[84]}
   );
   gpc606_5 gpc1272 (
      {stage1_5[274], stage1_5[275], stage1_5[276], stage1_5[277], stage1_5[278], stage1_5[279]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[35],stage2_7[69],stage2_6[77],stage2_5[85]}
   );
   gpc606_5 gpc1273 (
      {stage1_5[280], stage1_5[281], stage1_5[282], stage1_5[283], stage1_5[284], stage1_5[285]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[36],stage2_7[70],stage2_6[78],stage2_5[86]}
   );
   gpc606_5 gpc1274 (
      {stage1_5[286], stage1_5[287], stage1_5[288], stage1_5[289], stage1_5[290], stage1_5[291]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[37],stage2_7[71],stage2_6[79],stage2_5[87]}
   );
   gpc606_5 gpc1275 (
      {stage1_5[292], stage1_5[293], stage1_5[294], stage1_5[295], stage1_5[296], stage1_5[297]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[38],stage2_7[72],stage2_6[80],stage2_5[88]}
   );
   gpc606_5 gpc1276 (
      {stage1_5[298], stage1_5[299], stage1_5[300], stage1_5[301], stage1_5[302], stage1_5[303]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[39],stage2_7[73],stage2_6[81],stage2_5[89]}
   );
   gpc606_5 gpc1277 (
      {stage1_5[304], stage1_5[305], stage1_5[306], stage1_5[307], stage1_5[308], stage1_5[309]},
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77]},
      {stage2_9[12],stage2_8[40],stage2_7[74],stage2_6[82],stage2_5[90]}
   );
   gpc606_5 gpc1278 (
      {stage1_5[310], stage1_5[311], stage1_5[312], stage1_5[313], stage1_5[314], stage1_5[315]},
      {stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83]},
      {stage2_9[13],stage2_8[41],stage2_7[75],stage2_6[83],stage2_5[91]}
   );
   gpc606_5 gpc1279 (
      {stage1_5[316], stage1_5[317], stage1_5[318], stage1_5[319], stage1_5[320], stage1_5[321]},
      {stage1_7[84], stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage2_9[14],stage2_8[42],stage2_7[76],stage2_6[84],stage2_5[92]}
   );
   gpc606_5 gpc1280 (
      {stage1_6[168], stage1_6[169], stage1_6[170], stage1_6[171], stage1_6[172], stage1_6[173]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[15],stage2_8[43],stage2_7[77],stage2_6[85]}
   );
   gpc606_5 gpc1281 (
      {stage1_6[174], stage1_6[175], stage1_6[176], stage1_6[177], stage1_6[178], stage1_6[179]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[16],stage2_8[44],stage2_7[78],stage2_6[86]}
   );
   gpc606_5 gpc1282 (
      {stage1_6[180], stage1_6[181], stage1_6[182], stage1_6[183], stage1_6[184], stage1_6[185]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[17],stage2_8[45],stage2_7[79],stage2_6[87]}
   );
   gpc606_5 gpc1283 (
      {stage1_6[186], stage1_6[187], stage1_6[188], stage1_6[189], stage1_6[190], stage1_6[191]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[18],stage2_8[46],stage2_7[80],stage2_6[88]}
   );
   gpc615_5 gpc1284 (
      {stage1_6[192], stage1_6[193], stage1_6[194], stage1_6[195], stage1_6[196]},
      {stage1_7[90]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[19],stage2_8[47],stage2_7[81],stage2_6[89]}
   );
   gpc606_5 gpc1285 (
      {stage1_7[91], stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95], stage1_7[96]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[5],stage2_9[20],stage2_8[48],stage2_7[82]}
   );
   gpc606_5 gpc1286 (
      {stage1_7[97], stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101], stage1_7[102]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[6],stage2_9[21],stage2_8[49],stage2_7[83]}
   );
   gpc606_5 gpc1287 (
      {stage1_7[103], stage1_7[104], stage1_7[105], stage1_7[106], stage1_7[107], stage1_7[108]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[7],stage2_9[22],stage2_8[50],stage2_7[84]}
   );
   gpc606_5 gpc1288 (
      {stage1_7[109], stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113], stage1_7[114]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[8],stage2_9[23],stage2_8[51],stage2_7[85]}
   );
   gpc606_5 gpc1289 (
      {stage1_7[115], stage1_7[116], stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[9],stage2_9[24],stage2_8[52],stage2_7[86]}
   );
   gpc606_5 gpc1290 (
      {stage1_7[121], stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125], stage1_7[126]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[10],stage2_9[25],stage2_8[53],stage2_7[87]}
   );
   gpc606_5 gpc1291 (
      {stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130], stage1_7[131], stage1_7[132]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[11],stage2_9[26],stage2_8[54],stage2_7[88]}
   );
   gpc606_5 gpc1292 (
      {stage1_7[133], stage1_7[134], stage1_7[135], stage1_7[136], stage1_7[137], stage1_7[138]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[12],stage2_9[27],stage2_8[55],stage2_7[89]}
   );
   gpc606_5 gpc1293 (
      {stage1_7[139], stage1_7[140], stage1_7[141], stage1_7[142], stage1_7[143], stage1_7[144]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[13],stage2_9[28],stage2_8[56],stage2_7[90]}
   );
   gpc606_5 gpc1294 (
      {stage1_7[145], stage1_7[146], stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[14],stage2_9[29],stage2_8[57],stage2_7[91]}
   );
   gpc606_5 gpc1295 (
      {stage1_7[151], stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155], stage1_7[156]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[15],stage2_9[30],stage2_8[58],stage2_7[92]}
   );
   gpc606_5 gpc1296 (
      {stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160], stage1_7[161], stage1_7[162]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[16],stage2_9[31],stage2_8[59],stage2_7[93]}
   );
   gpc606_5 gpc1297 (
      {stage1_7[163], stage1_7[164], stage1_7[165], stage1_7[166], stage1_7[167], stage1_7[168]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[17],stage2_9[32],stage2_8[60],stage2_7[94]}
   );
   gpc606_5 gpc1298 (
      {stage1_7[169], stage1_7[170], stage1_7[171], stage1_7[172], stage1_7[173], stage1_7[174]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[18],stage2_9[33],stage2_8[61],stage2_7[95]}
   );
   gpc606_5 gpc1299 (
      {stage1_7[175], stage1_7[176], stage1_7[177], stage1_7[178], stage1_7[179], stage1_7[180]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[19],stage2_9[34],stage2_8[62],stage2_7[96]}
   );
   gpc606_5 gpc1300 (
      {stage1_7[181], stage1_7[182], stage1_7[183], stage1_7[184], stage1_7[185], stage1_7[186]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[20],stage2_9[35],stage2_8[63],stage2_7[97]}
   );
   gpc606_5 gpc1301 (
      {stage1_7[187], stage1_7[188], stage1_7[189], stage1_7[190], stage1_7[191], stage1_7[192]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[21],stage2_9[36],stage2_8[64],stage2_7[98]}
   );
   gpc606_5 gpc1302 (
      {stage1_7[193], stage1_7[194], stage1_7[195], stage1_7[196], stage1_7[197], stage1_7[198]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[22],stage2_9[37],stage2_8[65],stage2_7[99]}
   );
   gpc606_5 gpc1303 (
      {stage1_7[199], stage1_7[200], stage1_7[201], stage1_7[202], stage1_7[203], stage1_7[204]},
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage2_11[18],stage2_10[23],stage2_9[38],stage2_8[66],stage2_7[100]}
   );
   gpc606_5 gpc1304 (
      {stage1_7[205], stage1_7[206], stage1_7[207], stage1_7[208], stage1_7[209], stage1_7[210]},
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage2_11[19],stage2_10[24],stage2_9[39],stage2_8[67],stage2_7[101]}
   );
   gpc606_5 gpc1305 (
      {stage1_7[211], stage1_7[212], stage1_7[213], stage1_7[214], stage1_7[215], stage1_7[216]},
      {stage1_9[120], stage1_9[121], stage1_9[122], stage1_9[123], stage1_9[124], stage1_9[125]},
      {stage2_11[20],stage2_10[25],stage2_9[40],stage2_8[68],stage2_7[102]}
   );
   gpc606_5 gpc1306 (
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[21],stage2_10[26],stage2_9[41],stage2_8[69]}
   );
   gpc606_5 gpc1307 (
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[22],stage2_10[27],stage2_9[42],stage2_8[70]}
   );
   gpc606_5 gpc1308 (
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[23],stage2_10[28],stage2_9[43],stage2_8[71]}
   );
   gpc606_5 gpc1309 (
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[24],stage2_10[29],stage2_9[44],stage2_8[72]}
   );
   gpc606_5 gpc1310 (
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[25],stage2_10[30],stage2_9[45],stage2_8[73]}
   );
   gpc606_5 gpc1311 (
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[26],stage2_10[31],stage2_9[46],stage2_8[74]}
   );
   gpc606_5 gpc1312 (
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[27],stage2_10[32],stage2_9[47],stage2_8[75]}
   );
   gpc606_5 gpc1313 (
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[28],stage2_10[33],stage2_9[48],stage2_8[76]}
   );
   gpc606_5 gpc1314 (
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[29],stage2_10[34],stage2_9[49],stage2_8[77]}
   );
   gpc606_5 gpc1315 (
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[30],stage2_10[35],stage2_9[50],stage2_8[78]}
   );
   gpc606_5 gpc1316 (
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[31],stage2_10[36],stage2_9[51],stage2_8[79]}
   );
   gpc606_5 gpc1317 (
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[32],stage2_10[37],stage2_9[52],stage2_8[80]}
   );
   gpc606_5 gpc1318 (
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[33],stage2_10[38],stage2_9[53],stage2_8[81]}
   );
   gpc606_5 gpc1319 (
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[34],stage2_10[39],stage2_9[54],stage2_8[82]}
   );
   gpc606_5 gpc1320 (
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[35],stage2_10[40],stage2_9[55],stage2_8[83]}
   );
   gpc606_5 gpc1321 (
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[36],stage2_10[41],stage2_9[56],stage2_8[84]}
   );
   gpc606_5 gpc1322 (
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage2_12[16],stage2_11[37],stage2_10[42],stage2_9[57],stage2_8[85]}
   );
   gpc606_5 gpc1323 (
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106], stage1_10[107]},
      {stage2_12[17],stage2_11[38],stage2_10[43],stage2_9[58],stage2_8[86]}
   );
   gpc606_5 gpc1324 (
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142], stage1_8[143]},
      {stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage2_12[18],stage2_11[39],stage2_10[44],stage2_9[59],stage2_8[87]}
   );
   gpc606_5 gpc1325 (
      {stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147], stage1_8[148], stage1_8[149]},
      {stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119]},
      {stage2_12[19],stage2_11[40],stage2_10[45],stage2_9[60],stage2_8[88]}
   );
   gpc606_5 gpc1326 (
      {stage1_8[150], stage1_8[151], stage1_8[152], stage1_8[153], stage1_8[154], stage1_8[155]},
      {stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124], stage1_10[125]},
      {stage2_12[20],stage2_11[41],stage2_10[46],stage2_9[61],stage2_8[89]}
   );
   gpc606_5 gpc1327 (
      {stage1_8[156], stage1_8[157], stage1_8[158], stage1_8[159], stage1_8[160], stage1_8[161]},
      {stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130], stage1_10[131]},
      {stage2_12[21],stage2_11[42],stage2_10[47],stage2_9[62],stage2_8[90]}
   );
   gpc606_5 gpc1328 (
      {stage1_8[162], stage1_8[163], stage1_8[164], stage1_8[165], stage1_8[166], stage1_8[167]},
      {stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136], stage1_10[137]},
      {stage2_12[22],stage2_11[43],stage2_10[48],stage2_9[63],stage2_8[91]}
   );
   gpc606_5 gpc1329 (
      {stage1_8[168], stage1_8[169], stage1_8[170], stage1_8[171], stage1_8[172], stage1_8[173]},
      {stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141], stage1_10[142], stage1_10[143]},
      {stage2_12[23],stage2_11[44],stage2_10[49],stage2_9[64],stage2_8[92]}
   );
   gpc606_5 gpc1330 (
      {stage1_8[174], stage1_8[175], stage1_8[176], stage1_8[177], stage1_8[178], stage1_8[179]},
      {stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148], stage1_10[149]},
      {stage2_12[24],stage2_11[45],stage2_10[50],stage2_9[65],stage2_8[93]}
   );
   gpc615_5 gpc1331 (
      {stage1_8[180], stage1_8[181], stage1_8[182], stage1_8[183], stage1_8[184]},
      {stage1_9[126]},
      {stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154], stage1_10[155]},
      {stage2_12[25],stage2_11[46],stage2_10[51],stage2_9[66],stage2_8[94]}
   );
   gpc606_5 gpc1332 (
      {stage1_9[127], stage1_9[128], stage1_9[129], stage1_9[130], stage1_9[131], stage1_9[132]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[26],stage2_11[47],stage2_10[52],stage2_9[67]}
   );
   gpc606_5 gpc1333 (
      {stage1_9[133], stage1_9[134], stage1_9[135], stage1_9[136], stage1_9[137], stage1_9[138]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[27],stage2_11[48],stage2_10[53],stage2_9[68]}
   );
   gpc606_5 gpc1334 (
      {stage1_9[139], stage1_9[140], stage1_9[141], stage1_9[142], stage1_9[143], stage1_9[144]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[28],stage2_11[49],stage2_10[54],stage2_9[69]}
   );
   gpc606_5 gpc1335 (
      {stage1_9[145], stage1_9[146], stage1_9[147], stage1_9[148], stage1_9[149], stage1_9[150]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[29],stage2_11[50],stage2_10[55],stage2_9[70]}
   );
   gpc606_5 gpc1336 (
      {stage1_9[151], stage1_9[152], stage1_9[153], stage1_9[154], stage1_9[155], stage1_9[156]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[30],stage2_11[51],stage2_10[56],stage2_9[71]}
   );
   gpc606_5 gpc1337 (
      {stage1_9[157], stage1_9[158], stage1_9[159], stage1_9[160], stage1_9[161], stage1_9[162]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[31],stage2_11[52],stage2_10[57],stage2_9[72]}
   );
   gpc606_5 gpc1338 (
      {stage1_9[163], stage1_9[164], stage1_9[165], stage1_9[166], stage1_9[167], stage1_9[168]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[32],stage2_11[53],stage2_10[58],stage2_9[73]}
   );
   gpc606_5 gpc1339 (
      {stage1_9[169], stage1_9[170], stage1_9[171], stage1_9[172], stage1_9[173], stage1_9[174]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[33],stage2_11[54],stage2_10[59],stage2_9[74]}
   );
   gpc606_5 gpc1340 (
      {stage1_9[175], stage1_9[176], stage1_9[177], stage1_9[178], stage1_9[179], stage1_9[180]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[34],stage2_11[55],stage2_10[60],stage2_9[75]}
   );
   gpc606_5 gpc1341 (
      {stage1_9[181], stage1_9[182], stage1_9[183], stage1_9[184], stage1_9[185], stage1_9[186]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[35],stage2_11[56],stage2_10[61],stage2_9[76]}
   );
   gpc606_5 gpc1342 (
      {stage1_9[187], stage1_9[188], stage1_9[189], stage1_9[190], stage1_9[191], stage1_9[192]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[36],stage2_11[57],stage2_10[62],stage2_9[77]}
   );
   gpc606_5 gpc1343 (
      {stage1_9[193], stage1_9[194], stage1_9[195], stage1_9[196], stage1_9[197], stage1_9[198]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[37],stage2_11[58],stage2_10[63],stage2_9[78]}
   );
   gpc606_5 gpc1344 (
      {stage1_9[199], stage1_9[200], stage1_9[201], stage1_9[202], stage1_9[203], stage1_9[204]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[38],stage2_11[59],stage2_10[64],stage2_9[79]}
   );
   gpc606_5 gpc1345 (
      {stage1_9[205], stage1_9[206], stage1_9[207], stage1_9[208], stage1_9[209], stage1_9[210]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[39],stage2_11[60],stage2_10[65],stage2_9[80]}
   );
   gpc606_5 gpc1346 (
      {stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160], stage1_10[161]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[14],stage2_12[40],stage2_11[61],stage2_10[66]}
   );
   gpc606_5 gpc1347 (
      {stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166], stage1_10[167]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[15],stage2_12[41],stage2_11[62],stage2_10[67]}
   );
   gpc606_5 gpc1348 (
      {stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171], stage1_10[172], stage1_10[173]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[16],stage2_12[42],stage2_11[63],stage2_10[68]}
   );
   gpc606_5 gpc1349 (
      {stage1_10[174], stage1_10[175], stage1_10[176], stage1_10[177], stage1_10[178], stage1_10[179]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[17],stage2_12[43],stage2_11[64],stage2_10[69]}
   );
   gpc606_5 gpc1350 (
      {stage1_10[180], stage1_10[181], stage1_10[182], stage1_10[183], stage1_10[184], stage1_10[185]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[18],stage2_12[44],stage2_11[65],stage2_10[70]}
   );
   gpc606_5 gpc1351 (
      {stage1_10[186], stage1_10[187], stage1_10[188], stage1_10[189], stage1_10[190], stage1_10[191]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[19],stage2_12[45],stage2_11[66],stage2_10[71]}
   );
   gpc606_5 gpc1352 (
      {stage1_10[192], stage1_10[193], stage1_10[194], stage1_10[195], stage1_10[196], stage1_10[197]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[20],stage2_12[46],stage2_11[67],stage2_10[72]}
   );
   gpc606_5 gpc1353 (
      {stage1_10[198], stage1_10[199], stage1_10[200], stage1_10[201], stage1_10[202], stage1_10[203]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[21],stage2_12[47],stage2_11[68],stage2_10[73]}
   );
   gpc606_5 gpc1354 (
      {stage1_10[204], stage1_10[205], stage1_10[206], stage1_10[207], stage1_10[208], stage1_10[209]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[22],stage2_12[48],stage2_11[69],stage2_10[74]}
   );
   gpc606_5 gpc1355 (
      {stage1_10[210], stage1_10[211], stage1_10[212], stage1_10[213], stage1_10[214], stage1_10[215]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[23],stage2_12[49],stage2_11[70],stage2_10[75]}
   );
   gpc615_5 gpc1356 (
      {stage1_10[216], stage1_10[217], stage1_10[218], stage1_10[219], stage1_10[220]},
      {stage1_11[84]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[24],stage2_12[50],stage2_11[71],stage2_10[76]}
   );
   gpc615_5 gpc1357 (
      {stage1_10[221], stage1_10[222], stage1_10[223], stage1_10[224], stage1_10[225]},
      {stage1_11[85]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[25],stage2_12[51],stage2_11[72],stage2_10[77]}
   );
   gpc615_5 gpc1358 (
      {stage1_10[226], stage1_10[227], stage1_10[228], stage1_10[229], stage1_10[230]},
      {stage1_11[86]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[26],stage2_12[52],stage2_11[73],stage2_10[78]}
   );
   gpc615_5 gpc1359 (
      {stage1_10[231], stage1_10[232], stage1_10[233], stage1_10[234], stage1_10[235]},
      {stage1_11[87]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[27],stage2_12[53],stage2_11[74],stage2_10[79]}
   );
   gpc615_5 gpc1360 (
      {stage1_10[236], stage1_10[237], stage1_10[238], stage1_10[239], stage1_10[240]},
      {stage1_11[88]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[28],stage2_12[54],stage2_11[75],stage2_10[80]}
   );
   gpc615_5 gpc1361 (
      {stage1_10[241], stage1_10[242], stage1_10[243], stage1_10[244], stage1_10[245]},
      {stage1_11[89]},
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage2_14[15],stage2_13[29],stage2_12[55],stage2_11[76],stage2_10[81]}
   );
   gpc615_5 gpc1362 (
      {stage1_10[246], stage1_10[247], stage1_10[248], stage1_10[249], stage1_10[250]},
      {stage1_11[90]},
      {stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage2_14[16],stage2_13[30],stage2_12[56],stage2_11[77],stage2_10[82]}
   );
   gpc615_5 gpc1363 (
      {stage1_10[251], stage1_10[252], stage1_10[253], stage1_10[254], stage1_10[255]},
      {stage1_11[91]},
      {stage1_12[102], stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107]},
      {stage2_14[17],stage2_13[31],stage2_12[57],stage2_11[78],stage2_10[83]}
   );
   gpc615_5 gpc1364 (
      {stage1_10[256], stage1_10[257], stage1_10[258], stage1_10[259], stage1_10[260]},
      {stage1_11[92]},
      {stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113]},
      {stage2_14[18],stage2_13[32],stage2_12[58],stage2_11[79],stage2_10[84]}
   );
   gpc615_5 gpc1365 (
      {stage1_10[261], stage1_10[262], stage1_10[263], stage1_10[264], stage1_10[265]},
      {stage1_11[93]},
      {stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage2_14[19],stage2_13[33],stage2_12[59],stage2_11[80],stage2_10[85]}
   );
   gpc615_5 gpc1366 (
      {stage1_10[266], stage1_10[267], stage1_10[268], stage1_10[269], stage1_10[270]},
      {stage1_11[94]},
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125]},
      {stage2_14[20],stage2_13[34],stage2_12[60],stage2_11[81],stage2_10[86]}
   );
   gpc615_5 gpc1367 (
      {stage1_10[271], stage1_10[272], stage1_10[273], stage1_10[274], stage1_10[275]},
      {stage1_11[95]},
      {stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131]},
      {stage2_14[21],stage2_13[35],stage2_12[61],stage2_11[82],stage2_10[87]}
   );
   gpc615_5 gpc1368 (
      {stage1_10[276], stage1_10[277], stage1_10[278], stage1_10[279], stage1_10[280]},
      {stage1_11[96]},
      {stage1_12[132], stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136], stage1_12[137]},
      {stage2_14[22],stage2_13[36],stage2_12[62],stage2_11[83],stage2_10[88]}
   );
   gpc606_5 gpc1369 (
      {stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101], stage1_11[102]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[23],stage2_13[37],stage2_12[63],stage2_11[84]}
   );
   gpc606_5 gpc1370 (
      {stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[24],stage2_13[38],stage2_12[64],stage2_11[85]}
   );
   gpc615_5 gpc1371 (
      {stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113]},
      {stage1_12[138]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[25],stage2_13[39],stage2_12[65],stage2_11[86]}
   );
   gpc615_5 gpc1372 (
      {stage1_11[114], stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118]},
      {stage1_12[139]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[26],stage2_13[40],stage2_12[66],stage2_11[87]}
   );
   gpc615_5 gpc1373 (
      {stage1_11[119], stage1_11[120], stage1_11[121], stage1_11[122], stage1_11[123]},
      {stage1_12[140]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[27],stage2_13[41],stage2_12[67],stage2_11[88]}
   );
   gpc615_5 gpc1374 (
      {stage1_11[124], stage1_11[125], stage1_11[126], stage1_11[127], stage1_11[128]},
      {stage1_12[141]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[28],stage2_13[42],stage2_12[68],stage2_11[89]}
   );
   gpc615_5 gpc1375 (
      {stage1_11[129], stage1_11[130], stage1_11[131], stage1_11[132], stage1_11[133]},
      {stage1_12[142]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[29],stage2_13[43],stage2_12[69],stage2_11[90]}
   );
   gpc615_5 gpc1376 (
      {stage1_11[134], stage1_11[135], stage1_11[136], stage1_11[137], stage1_11[138]},
      {stage1_12[143]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[30],stage2_13[44],stage2_12[70],stage2_11[91]}
   );
   gpc615_5 gpc1377 (
      {stage1_11[139], stage1_11[140], stage1_11[141], stage1_11[142], stage1_11[143]},
      {stage1_12[144]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[31],stage2_13[45],stage2_12[71],stage2_11[92]}
   );
   gpc615_5 gpc1378 (
      {stage1_11[144], stage1_11[145], stage1_11[146], stage1_11[147], stage1_11[148]},
      {stage1_12[145]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[32],stage2_13[46],stage2_12[72],stage2_11[93]}
   );
   gpc615_5 gpc1379 (
      {stage1_11[149], stage1_11[150], stage1_11[151], stage1_11[152], stage1_11[153]},
      {stage1_12[146]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[33],stage2_13[47],stage2_12[73],stage2_11[94]}
   );
   gpc615_5 gpc1380 (
      {stage1_11[154], stage1_11[155], stage1_11[156], stage1_11[157], stage1_11[158]},
      {stage1_12[147]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[34],stage2_13[48],stage2_12[74],stage2_11[95]}
   );
   gpc615_5 gpc1381 (
      {stage1_11[159], stage1_11[160], stage1_11[161], stage1_11[162], stage1_11[163]},
      {stage1_12[148]},
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage2_15[12],stage2_14[35],stage2_13[49],stage2_12[75],stage2_11[96]}
   );
   gpc615_5 gpc1382 (
      {stage1_11[164], stage1_11[165], stage1_11[166], stage1_11[167], stage1_11[168]},
      {stage1_12[149]},
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage2_15[13],stage2_14[36],stage2_13[50],stage2_12[76],stage2_11[97]}
   );
   gpc615_5 gpc1383 (
      {stage1_11[169], stage1_11[170], stage1_11[171], stage1_11[172], stage1_11[173]},
      {stage1_12[150]},
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage2_15[14],stage2_14[37],stage2_13[51],stage2_12[77],stage2_11[98]}
   );
   gpc615_5 gpc1384 (
      {stage1_11[174], stage1_11[175], stage1_11[176], stage1_11[177], stage1_11[178]},
      {stage1_12[151]},
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage2_15[15],stage2_14[38],stage2_13[52],stage2_12[78],stage2_11[99]}
   );
   gpc615_5 gpc1385 (
      {stage1_11[179], stage1_11[180], stage1_11[181], stage1_11[182], stage1_11[183]},
      {stage1_12[152]},
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage2_15[16],stage2_14[39],stage2_13[53],stage2_12[79],stage2_11[100]}
   );
   gpc615_5 gpc1386 (
      {stage1_11[184], stage1_11[185], stage1_11[186], stage1_11[187], stage1_11[188]},
      {stage1_12[153]},
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage2_15[17],stage2_14[40],stage2_13[54],stage2_12[80],stage2_11[101]}
   );
   gpc615_5 gpc1387 (
      {stage1_11[189], stage1_11[190], stage1_11[191], stage1_11[192], stage1_11[193]},
      {stage1_12[154]},
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage2_15[18],stage2_14[41],stage2_13[55],stage2_12[81],stage2_11[102]}
   );
   gpc615_5 gpc1388 (
      {stage1_11[194], stage1_11[195], stage1_11[196], stage1_11[197], stage1_11[198]},
      {stage1_12[155]},
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage2_15[19],stage2_14[42],stage2_13[56],stage2_12[82],stage2_11[103]}
   );
   gpc615_5 gpc1389 (
      {stage1_11[199], stage1_11[200], stage1_11[201], stage1_11[202], stage1_11[203]},
      {stage1_12[156]},
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage2_15[20],stage2_14[43],stage2_13[57],stage2_12[83],stage2_11[104]}
   );
   gpc615_5 gpc1390 (
      {stage1_11[204], stage1_11[205], stage1_11[206], stage1_11[207], stage1_11[208]},
      {stage1_12[157]},
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage2_15[21],stage2_14[44],stage2_13[58],stage2_12[84],stage2_11[105]}
   );
   gpc615_5 gpc1391 (
      {stage1_11[209], stage1_11[210], stage1_11[211], stage1_11[212], stage1_11[213]},
      {stage1_12[158]},
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136], stage1_13[137]},
      {stage2_15[22],stage2_14[45],stage2_13[59],stage2_12[85],stage2_11[106]}
   );
   gpc606_5 gpc1392 (
      {stage1_12[159], stage1_12[160], stage1_12[161], stage1_12[162], stage1_12[163], stage1_12[164]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[23],stage2_14[46],stage2_13[60],stage2_12[86]}
   );
   gpc606_5 gpc1393 (
      {stage1_12[165], stage1_12[166], stage1_12[167], stage1_12[168], stage1_12[169], stage1_12[170]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[24],stage2_14[47],stage2_13[61],stage2_12[87]}
   );
   gpc606_5 gpc1394 (
      {stage1_12[171], stage1_12[172], stage1_12[173], stage1_12[174], stage1_12[175], stage1_12[176]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[25],stage2_14[48],stage2_13[62],stage2_12[88]}
   );
   gpc606_5 gpc1395 (
      {stage1_12[177], stage1_12[178], stage1_12[179], stage1_12[180], stage1_12[181], stage1_12[182]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[26],stage2_14[49],stage2_13[63],stage2_12[89]}
   );
   gpc606_5 gpc1396 (
      {stage1_12[183], stage1_12[184], stage1_12[185], stage1_12[186], stage1_12[187], stage1_12[188]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[27],stage2_14[50],stage2_13[64],stage2_12[90]}
   );
   gpc606_5 gpc1397 (
      {stage1_12[189], stage1_12[190], stage1_12[191], stage1_12[192], stage1_12[193], stage1_12[194]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[28],stage2_14[51],stage2_13[65],stage2_12[91]}
   );
   gpc606_5 gpc1398 (
      {stage1_12[195], stage1_12[196], stage1_12[197], stage1_12[198], stage1_12[199], stage1_12[200]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[29],stage2_14[52],stage2_13[66],stage2_12[92]}
   );
   gpc606_5 gpc1399 (
      {stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141], stage1_13[142], stage1_13[143]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[7],stage2_15[30],stage2_14[53],stage2_13[67]}
   );
   gpc606_5 gpc1400 (
      {stage1_13[144], stage1_13[145], stage1_13[146], stage1_13[147], stage1_13[148], stage1_13[149]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[8],stage2_15[31],stage2_14[54],stage2_13[68]}
   );
   gpc615_5 gpc1401 (
      {stage1_13[150], stage1_13[151], stage1_13[152], stage1_13[153], stage1_13[154]},
      {stage1_14[42]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[9],stage2_15[32],stage2_14[55],stage2_13[69]}
   );
   gpc615_5 gpc1402 (
      {stage1_13[155], stage1_13[156], stage1_13[157], stage1_13[158], stage1_13[159]},
      {stage1_14[43]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[10],stage2_15[33],stage2_14[56],stage2_13[70]}
   );
   gpc615_5 gpc1403 (
      {stage1_13[160], stage1_13[161], stage1_13[162], stage1_13[163], stage1_13[164]},
      {stage1_14[44]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[11],stage2_15[34],stage2_14[57],stage2_13[71]}
   );
   gpc615_5 gpc1404 (
      {stage1_13[165], stage1_13[166], stage1_13[167], stage1_13[168], stage1_13[169]},
      {stage1_14[45]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[12],stage2_15[35],stage2_14[58],stage2_13[72]}
   );
   gpc615_5 gpc1405 (
      {stage1_13[170], stage1_13[171], stage1_13[172], stage1_13[173], stage1_13[174]},
      {stage1_14[46]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[13],stage2_15[36],stage2_14[59],stage2_13[73]}
   );
   gpc615_5 gpc1406 (
      {stage1_13[175], stage1_13[176], stage1_13[177], stage1_13[178], stage1_13[179]},
      {stage1_14[47]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[14],stage2_15[37],stage2_14[60],stage2_13[74]}
   );
   gpc615_5 gpc1407 (
      {stage1_13[180], stage1_13[181], stage1_13[182], stage1_13[183], stage1_13[184]},
      {stage1_14[48]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage2_17[8],stage2_16[15],stage2_15[38],stage2_14[61],stage2_13[75]}
   );
   gpc615_5 gpc1408 (
      {stage1_13[185], stage1_13[186], stage1_13[187], stage1_13[188], stage1_13[189]},
      {stage1_14[49]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage2_17[9],stage2_16[16],stage2_15[39],stage2_14[62],stage2_13[76]}
   );
   gpc615_5 gpc1409 (
      {stage1_13[190], stage1_13[191], stage1_13[192], stage1_13[193], stage1_13[194]},
      {stage1_14[50]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage2_17[10],stage2_16[17],stage2_15[40],stage2_14[63],stage2_13[77]}
   );
   gpc615_5 gpc1410 (
      {stage1_13[195], stage1_13[196], stage1_13[197], stage1_13[198], stage1_13[199]},
      {stage1_14[51]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage2_17[11],stage2_16[18],stage2_15[41],stage2_14[64],stage2_13[78]}
   );
   gpc615_5 gpc1411 (
      {stage1_13[200], stage1_13[201], stage1_13[202], stage1_13[203], stage1_13[204]},
      {stage1_14[52]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage2_17[12],stage2_16[19],stage2_15[42],stage2_14[65],stage2_13[79]}
   );
   gpc615_5 gpc1412 (
      {stage1_13[205], stage1_13[206], stage1_13[207], stage1_13[208], stage1_13[209]},
      {stage1_14[53]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage2_17[13],stage2_16[20],stage2_15[43],stage2_14[66],stage2_13[80]}
   );
   gpc615_5 gpc1413 (
      {stage1_13[210], stage1_13[211], stage1_13[212], stage1_13[213], stage1_13[214]},
      {stage1_14[54]},
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89]},
      {stage2_17[14],stage2_16[21],stage2_15[44],stage2_14[67],stage2_13[81]}
   );
   gpc615_5 gpc1414 (
      {stage1_13[215], stage1_13[216], stage1_13[217], stage1_13[218], stage1_13[219]},
      {stage1_14[55]},
      {stage1_15[90], stage1_15[91], stage1_15[92], stage1_15[93], stage1_15[94], stage1_15[95]},
      {stage2_17[15],stage2_16[22],stage2_15[45],stage2_14[68],stage2_13[82]}
   );
   gpc615_5 gpc1415 (
      {stage1_13[220], stage1_13[221], stage1_13[222], stage1_13[223], stage1_13[224]},
      {stage1_14[56]},
      {stage1_15[96], stage1_15[97], stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101]},
      {stage2_17[16],stage2_16[23],stage2_15[46],stage2_14[69],stage2_13[83]}
   );
   gpc615_5 gpc1416 (
      {stage1_13[225], stage1_13[226], stage1_13[227], stage1_13[228], stage1_13[229]},
      {stage1_14[57]},
      {stage1_15[102], stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage2_17[17],stage2_16[24],stage2_15[47],stage2_14[70],stage2_13[84]}
   );
   gpc615_5 gpc1417 (
      {stage1_13[230], stage1_13[231], stage1_13[232], stage1_13[233], stage1_13[234]},
      {stage1_14[58]},
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112], stage1_15[113]},
      {stage2_17[18],stage2_16[25],stage2_15[48],stage2_14[71],stage2_13[85]}
   );
   gpc606_5 gpc1418 (
      {stage1_14[59], stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[19],stage2_16[26],stage2_15[49],stage2_14[72]}
   );
   gpc606_5 gpc1419 (
      {stage1_14[65], stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[20],stage2_16[27],stage2_15[50],stage2_14[73]}
   );
   gpc606_5 gpc1420 (
      {stage1_14[71], stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[21],stage2_16[28],stage2_15[51],stage2_14[74]}
   );
   gpc606_5 gpc1421 (
      {stage1_14[77], stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[22],stage2_16[29],stage2_15[52],stage2_14[75]}
   );
   gpc606_5 gpc1422 (
      {stage1_14[83], stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[23],stage2_16[30],stage2_15[53],stage2_14[76]}
   );
   gpc606_5 gpc1423 (
      {stage1_14[89], stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[24],stage2_16[31],stage2_15[54],stage2_14[77]}
   );
   gpc606_5 gpc1424 (
      {stage1_14[95], stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[25],stage2_16[32],stage2_15[55],stage2_14[78]}
   );
   gpc606_5 gpc1425 (
      {stage1_14[101], stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[26],stage2_16[33],stage2_15[56],stage2_14[79]}
   );
   gpc606_5 gpc1426 (
      {stage1_14[107], stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111], stage1_14[112]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[27],stage2_16[34],stage2_15[57],stage2_14[80]}
   );
   gpc606_5 gpc1427 (
      {stage1_14[113], stage1_14[114], stage1_14[115], stage1_14[116], stage1_14[117], stage1_14[118]},
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage2_18[9],stage2_17[28],stage2_16[35],stage2_15[58],stage2_14[81]}
   );
   gpc615_5 gpc1428 (
      {stage1_14[119], stage1_14[120], stage1_14[121], stage1_14[122], stage1_14[123]},
      {stage1_15[114]},
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65]},
      {stage2_18[10],stage2_17[29],stage2_16[36],stage2_15[59],stage2_14[82]}
   );
   gpc615_5 gpc1429 (
      {stage1_14[124], stage1_14[125], stage1_14[126], stage1_14[127], stage1_14[128]},
      {stage1_15[115]},
      {stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71]},
      {stage2_18[11],stage2_17[30],stage2_16[37],stage2_15[60],stage2_14[83]}
   );
   gpc615_5 gpc1430 (
      {stage1_14[129], stage1_14[130], stage1_14[131], stage1_14[132], stage1_14[133]},
      {stage1_15[116]},
      {stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77]},
      {stage2_18[12],stage2_17[31],stage2_16[38],stage2_15[61],stage2_14[84]}
   );
   gpc615_5 gpc1431 (
      {stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137], stage1_14[138]},
      {stage1_15[117]},
      {stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83]},
      {stage2_18[13],stage2_17[32],stage2_16[39],stage2_15[62],stage2_14[85]}
   );
   gpc615_5 gpc1432 (
      {stage1_14[139], stage1_14[140], stage1_14[141], stage1_14[142], stage1_14[143]},
      {stage1_15[118]},
      {stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage2_18[14],stage2_17[33],stage2_16[40],stage2_15[63],stage2_14[86]}
   );
   gpc615_5 gpc1433 (
      {stage1_14[144], stage1_14[145], stage1_14[146], stage1_14[147], stage1_14[148]},
      {stage1_15[119]},
      {stage1_16[90], stage1_16[91], stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95]},
      {stage2_18[15],stage2_17[34],stage2_16[41],stage2_15[64],stage2_14[87]}
   );
   gpc615_5 gpc1434 (
      {stage1_14[149], stage1_14[150], stage1_14[151], stage1_14[152], stage1_14[153]},
      {stage1_15[120]},
      {stage1_16[96], stage1_16[97], stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101]},
      {stage2_18[16],stage2_17[35],stage2_16[42],stage2_15[65],stage2_14[88]}
   );
   gpc615_5 gpc1435 (
      {stage1_14[154], stage1_14[155], stage1_14[156], stage1_14[157], stage1_14[158]},
      {stage1_15[121]},
      {stage1_16[102], stage1_16[103], stage1_16[104], stage1_16[105], stage1_16[106], stage1_16[107]},
      {stage2_18[17],stage2_17[36],stage2_16[43],stage2_15[66],stage2_14[89]}
   );
   gpc615_5 gpc1436 (
      {stage1_14[159], stage1_14[160], stage1_14[161], stage1_14[162], stage1_14[163]},
      {stage1_15[122]},
      {stage1_16[108], stage1_16[109], stage1_16[110], stage1_16[111], stage1_16[112], stage1_16[113]},
      {stage2_18[18],stage2_17[37],stage2_16[44],stage2_15[67],stage2_14[90]}
   );
   gpc615_5 gpc1437 (
      {stage1_14[164], stage1_14[165], stage1_14[166], stage1_14[167], stage1_14[168]},
      {stage1_15[123]},
      {stage1_16[114], stage1_16[115], stage1_16[116], stage1_16[117], stage1_16[118], stage1_16[119]},
      {stage2_18[19],stage2_17[38],stage2_16[45],stage2_15[68],stage2_14[91]}
   );
   gpc615_5 gpc1438 (
      {stage1_14[169], stage1_14[170], stage1_14[171], stage1_14[172], stage1_14[173]},
      {stage1_15[124]},
      {stage1_16[120], stage1_16[121], stage1_16[122], stage1_16[123], stage1_16[124], stage1_16[125]},
      {stage2_18[20],stage2_17[39],stage2_16[46],stage2_15[69],stage2_14[92]}
   );
   gpc606_5 gpc1439 (
      {stage1_15[125], stage1_15[126], stage1_15[127], stage1_15[128], stage1_15[129], stage1_15[130]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[21],stage2_17[40],stage2_16[47],stage2_15[70]}
   );
   gpc606_5 gpc1440 (
      {stage1_15[131], stage1_15[132], stage1_15[133], stage1_15[134], stage1_15[135], stage1_15[136]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[22],stage2_17[41],stage2_16[48],stage2_15[71]}
   );
   gpc606_5 gpc1441 (
      {stage1_15[137], stage1_15[138], stage1_15[139], stage1_15[140], stage1_15[141], stage1_15[142]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[23],stage2_17[42],stage2_16[49],stage2_15[72]}
   );
   gpc606_5 gpc1442 (
      {stage1_15[143], stage1_15[144], stage1_15[145], stage1_15[146], stage1_15[147], stage1_15[148]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[24],stage2_17[43],stage2_16[50],stage2_15[73]}
   );
   gpc606_5 gpc1443 (
      {stage1_15[149], stage1_15[150], stage1_15[151], stage1_15[152], stage1_15[153], stage1_15[154]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[25],stage2_17[44],stage2_16[51],stage2_15[74]}
   );
   gpc1_1 gpc1444 (
      {stage1_0[138]},
      {stage2_0[28]}
   );
   gpc1_1 gpc1445 (
      {stage1_0[139]},
      {stage2_0[29]}
   );
   gpc1_1 gpc1446 (
      {stage1_0[140]},
      {stage2_0[30]}
   );
   gpc1_1 gpc1447 (
      {stage1_0[141]},
      {stage2_0[31]}
   );
   gpc1_1 gpc1448 (
      {stage1_0[142]},
      {stage2_0[32]}
   );
   gpc1_1 gpc1449 (
      {stage1_0[143]},
      {stage2_0[33]}
   );
   gpc1_1 gpc1450 (
      {stage1_0[144]},
      {stage2_0[34]}
   );
   gpc1_1 gpc1451 (
      {stage1_0[145]},
      {stage2_0[35]}
   );
   gpc1_1 gpc1452 (
      {stage1_0[146]},
      {stage2_0[36]}
   );
   gpc1_1 gpc1453 (
      {stage1_0[147]},
      {stage2_0[37]}
   );
   gpc1_1 gpc1454 (
      {stage1_1[108]},
      {stage2_1[36]}
   );
   gpc1_1 gpc1455 (
      {stage1_1[109]},
      {stage2_1[37]}
   );
   gpc1_1 gpc1456 (
      {stage1_1[110]},
      {stage2_1[38]}
   );
   gpc1_1 gpc1457 (
      {stage1_1[111]},
      {stage2_1[39]}
   );
   gpc1_1 gpc1458 (
      {stage1_1[112]},
      {stage2_1[40]}
   );
   gpc1_1 gpc1459 (
      {stage1_1[113]},
      {stage2_1[41]}
   );
   gpc1_1 gpc1460 (
      {stage1_1[114]},
      {stage2_1[42]}
   );
   gpc1_1 gpc1461 (
      {stage1_1[115]},
      {stage2_1[43]}
   );
   gpc1_1 gpc1462 (
      {stage1_1[116]},
      {stage2_1[44]}
   );
   gpc1_1 gpc1463 (
      {stage1_1[117]},
      {stage2_1[45]}
   );
   gpc1_1 gpc1464 (
      {stage1_1[118]},
      {stage2_1[46]}
   );
   gpc1_1 gpc1465 (
      {stage1_1[119]},
      {stage2_1[47]}
   );
   gpc1_1 gpc1466 (
      {stage1_1[120]},
      {stage2_1[48]}
   );
   gpc1_1 gpc1467 (
      {stage1_1[121]},
      {stage2_1[49]}
   );
   gpc1_1 gpc1468 (
      {stage1_1[122]},
      {stage2_1[50]}
   );
   gpc1_1 gpc1469 (
      {stage1_1[123]},
      {stage2_1[51]}
   );
   gpc1_1 gpc1470 (
      {stage1_1[124]},
      {stage2_1[52]}
   );
   gpc1_1 gpc1471 (
      {stage1_1[125]},
      {stage2_1[53]}
   );
   gpc1_1 gpc1472 (
      {stage1_1[126]},
      {stage2_1[54]}
   );
   gpc1_1 gpc1473 (
      {stage1_1[127]},
      {stage2_1[55]}
   );
   gpc1_1 gpc1474 (
      {stage1_1[128]},
      {stage2_1[56]}
   );
   gpc1_1 gpc1475 (
      {stage1_1[129]},
      {stage2_1[57]}
   );
   gpc1_1 gpc1476 (
      {stage1_1[130]},
      {stage2_1[58]}
   );
   gpc1_1 gpc1477 (
      {stage1_1[131]},
      {stage2_1[59]}
   );
   gpc1_1 gpc1478 (
      {stage1_1[132]},
      {stage2_1[60]}
   );
   gpc1_1 gpc1479 (
      {stage1_1[133]},
      {stage2_1[61]}
   );
   gpc1_1 gpc1480 (
      {stage1_1[134]},
      {stage2_1[62]}
   );
   gpc1_1 gpc1481 (
      {stage1_2[158]},
      {stage2_2[44]}
   );
   gpc1_1 gpc1482 (
      {stage1_2[159]},
      {stage2_2[45]}
   );
   gpc1_1 gpc1483 (
      {stage1_2[160]},
      {stage2_2[46]}
   );
   gpc1_1 gpc1484 (
      {stage1_2[161]},
      {stage2_2[47]}
   );
   gpc1_1 gpc1485 (
      {stage1_2[162]},
      {stage2_2[48]}
   );
   gpc1_1 gpc1486 (
      {stage1_2[163]},
      {stage2_2[49]}
   );
   gpc1_1 gpc1487 (
      {stage1_2[164]},
      {stage2_2[50]}
   );
   gpc1_1 gpc1488 (
      {stage1_2[165]},
      {stage2_2[51]}
   );
   gpc1_1 gpc1489 (
      {stage1_2[166]},
      {stage2_2[52]}
   );
   gpc1_1 gpc1490 (
      {stage1_2[167]},
      {stage2_2[53]}
   );
   gpc1_1 gpc1491 (
      {stage1_3[236]},
      {stage2_3[78]}
   );
   gpc1_1 gpc1492 (
      {stage1_3[237]},
      {stage2_3[79]}
   );
   gpc1_1 gpc1493 (
      {stage1_3[238]},
      {stage2_3[80]}
   );
   gpc1_1 gpc1494 (
      {stage1_3[239]},
      {stage2_3[81]}
   );
   gpc1_1 gpc1495 (
      {stage1_3[240]},
      {stage2_3[82]}
   );
   gpc1_1 gpc1496 (
      {stage1_3[241]},
      {stage2_3[83]}
   );
   gpc1_1 gpc1497 (
      {stage1_3[242]},
      {stage2_3[84]}
   );
   gpc1_1 gpc1498 (
      {stage1_3[243]},
      {stage2_3[85]}
   );
   gpc1_1 gpc1499 (
      {stage1_4[222]},
      {stage2_4[106]}
   );
   gpc1_1 gpc1500 (
      {stage1_5[322]},
      {stage2_5[93]}
   );
   gpc1_1 gpc1501 (
      {stage1_5[323]},
      {stage2_5[94]}
   );
   gpc1_1 gpc1502 (
      {stage1_5[324]},
      {stage2_5[95]}
   );
   gpc1_1 gpc1503 (
      {stage1_5[325]},
      {stage2_5[96]}
   );
   gpc1_1 gpc1504 (
      {stage1_5[326]},
      {stage2_5[97]}
   );
   gpc1_1 gpc1505 (
      {stage1_5[327]},
      {stage2_5[98]}
   );
   gpc1_1 gpc1506 (
      {stage1_5[328]},
      {stage2_5[99]}
   );
   gpc1_1 gpc1507 (
      {stage1_5[329]},
      {stage2_5[100]}
   );
   gpc1_1 gpc1508 (
      {stage1_5[330]},
      {stage2_5[101]}
   );
   gpc1_1 gpc1509 (
      {stage1_5[331]},
      {stage2_5[102]}
   );
   gpc1_1 gpc1510 (
      {stage1_5[332]},
      {stage2_5[103]}
   );
   gpc1_1 gpc1511 (
      {stage1_5[333]},
      {stage2_5[104]}
   );
   gpc1_1 gpc1512 (
      {stage1_5[334]},
      {stage2_5[105]}
   );
   gpc1_1 gpc1513 (
      {stage1_5[335]},
      {stage2_5[106]}
   );
   gpc1_1 gpc1514 (
      {stage1_5[336]},
      {stage2_5[107]}
   );
   gpc1_1 gpc1515 (
      {stage1_8[185]},
      {stage2_8[95]}
   );
   gpc1_1 gpc1516 (
      {stage1_8[186]},
      {stage2_8[96]}
   );
   gpc1_1 gpc1517 (
      {stage1_8[187]},
      {stage2_8[97]}
   );
   gpc1_1 gpc1518 (
      {stage1_8[188]},
      {stage2_8[98]}
   );
   gpc1_1 gpc1519 (
      {stage1_8[189]},
      {stage2_8[99]}
   );
   gpc1_1 gpc1520 (
      {stage1_8[190]},
      {stage2_8[100]}
   );
   gpc1_1 gpc1521 (
      {stage1_8[191]},
      {stage2_8[101]}
   );
   gpc1_1 gpc1522 (
      {stage1_8[192]},
      {stage2_8[102]}
   );
   gpc1_1 gpc1523 (
      {stage1_8[193]},
      {stage2_8[103]}
   );
   gpc1_1 gpc1524 (
      {stage1_8[194]},
      {stage2_8[104]}
   );
   gpc1_1 gpc1525 (
      {stage1_8[195]},
      {stage2_8[105]}
   );
   gpc1_1 gpc1526 (
      {stage1_10[281]},
      {stage2_10[89]}
   );
   gpc1_1 gpc1527 (
      {stage1_12[201]},
      {stage2_12[93]}
   );
   gpc1_1 gpc1528 (
      {stage1_14[174]},
      {stage2_14[93]}
   );
   gpc1_1 gpc1529 (
      {stage1_14[175]},
      {stage2_14[94]}
   );
   gpc1_1 gpc1530 (
      {stage1_14[176]},
      {stage2_14[95]}
   );
   gpc1_1 gpc1531 (
      {stage1_14[177]},
      {stage2_14[96]}
   );
   gpc1_1 gpc1532 (
      {stage1_14[178]},
      {stage2_14[97]}
   );
   gpc1_1 gpc1533 (
      {stage1_14[179]},
      {stage2_14[98]}
   );
   gpc1_1 gpc1534 (
      {stage1_14[180]},
      {stage2_14[99]}
   );
   gpc1_1 gpc1535 (
      {stage1_14[181]},
      {stage2_14[100]}
   );
   gpc1_1 gpc1536 (
      {stage1_14[182]},
      {stage2_14[101]}
   );
   gpc1_1 gpc1537 (
      {stage1_16[126]},
      {stage2_16[52]}
   );
   gpc1_1 gpc1538 (
      {stage1_16[127]},
      {stage2_16[53]}
   );
   gpc1_1 gpc1539 (
      {stage1_16[128]},
      {stage2_16[54]}
   );
   gpc1_1 gpc1540 (
      {stage1_16[129]},
      {stage2_16[55]}
   );
   gpc1_1 gpc1541 (
      {stage1_16[130]},
      {stage2_16[56]}
   );
   gpc1_1 gpc1542 (
      {stage1_16[131]},
      {stage2_16[57]}
   );
   gpc1_1 gpc1543 (
      {stage1_16[132]},
      {stage2_16[58]}
   );
   gpc1_1 gpc1544 (
      {stage1_16[133]},
      {stage2_16[59]}
   );
   gpc1_1 gpc1545 (
      {stage1_16[134]},
      {stage2_16[60]}
   );
   gpc1_1 gpc1546 (
      {stage1_16[135]},
      {stage2_16[61]}
   );
   gpc1_1 gpc1547 (
      {stage1_16[136]},
      {stage2_16[62]}
   );
   gpc1_1 gpc1548 (
      {stage1_16[137]},
      {stage2_16[63]}
   );
   gpc1_1 gpc1549 (
      {stage1_16[138]},
      {stage2_16[64]}
   );
   gpc1_1 gpc1550 (
      {stage1_16[139]},
      {stage2_16[65]}
   );
   gpc1_1 gpc1551 (
      {stage1_16[140]},
      {stage2_16[66]}
   );
   gpc1_1 gpc1552 (
      {stage1_16[141]},
      {stage2_16[67]}
   );
   gpc1_1 gpc1553 (
      {stage1_16[142]},
      {stage2_16[68]}
   );
   gpc1_1 gpc1554 (
      {stage1_16[143]},
      {stage2_16[69]}
   );
   gpc1_1 gpc1555 (
      {stage1_16[144]},
      {stage2_16[70]}
   );
   gpc1_1 gpc1556 (
      {stage1_16[145]},
      {stage2_16[71]}
   );
   gpc1_1 gpc1557 (
      {stage1_16[146]},
      {stage2_16[72]}
   );
   gpc1_1 gpc1558 (
      {stage1_16[147]},
      {stage2_16[73]}
   );
   gpc1_1 gpc1559 (
      {stage1_16[148]},
      {stage2_16[74]}
   );
   gpc1_1 gpc1560 (
      {stage1_16[149]},
      {stage2_16[75]}
   );
   gpc1_1 gpc1561 (
      {stage1_16[150]},
      {stage2_16[76]}
   );
   gpc1_1 gpc1562 (
      {stage1_17[30]},
      {stage2_17[45]}
   );
   gpc1_1 gpc1563 (
      {stage1_17[31]},
      {stage2_17[46]}
   );
   gpc1_1 gpc1564 (
      {stage1_17[32]},
      {stage2_17[47]}
   );
   gpc1_1 gpc1565 (
      {stage1_17[33]},
      {stage2_17[48]}
   );
   gpc1_1 gpc1566 (
      {stage1_17[34]},
      {stage2_17[49]}
   );
   gpc1_1 gpc1567 (
      {stage1_17[35]},
      {stage2_17[50]}
   );
   gpc1_1 gpc1568 (
      {stage1_17[36]},
      {stage2_17[51]}
   );
   gpc1_1 gpc1569 (
      {stage1_17[37]},
      {stage2_17[52]}
   );
   gpc1_1 gpc1570 (
      {stage1_17[38]},
      {stage2_17[53]}
   );
   gpc1_1 gpc1571 (
      {stage1_17[39]},
      {stage2_17[54]}
   );
   gpc1_1 gpc1572 (
      {stage1_17[40]},
      {stage2_17[55]}
   );
   gpc1_1 gpc1573 (
      {stage1_17[41]},
      {stage2_17[56]}
   );
   gpc1_1 gpc1574 (
      {stage1_17[42]},
      {stage2_17[57]}
   );
   gpc1_1 gpc1575 (
      {stage1_17[43]},
      {stage2_17[58]}
   );
   gpc1_1 gpc1576 (
      {stage1_17[44]},
      {stage2_17[59]}
   );
   gpc1_1 gpc1577 (
      {stage1_17[45]},
      {stage2_17[60]}
   );
   gpc1_1 gpc1578 (
      {stage1_17[46]},
      {stage2_17[61]}
   );
   gpc1_1 gpc1579 (
      {stage1_17[47]},
      {stage2_17[62]}
   );
   gpc1_1 gpc1580 (
      {stage1_17[48]},
      {stage2_17[63]}
   );
   gpc1_1 gpc1581 (
      {stage1_17[49]},
      {stage2_17[64]}
   );
   gpc1_1 gpc1582 (
      {stage1_17[50]},
      {stage2_17[65]}
   );
   gpc1_1 gpc1583 (
      {stage1_17[51]},
      {stage2_17[66]}
   );
   gpc1_1 gpc1584 (
      {stage1_17[52]},
      {stage2_17[67]}
   );
   gpc1_1 gpc1585 (
      {stage1_17[53]},
      {stage2_17[68]}
   );
   gpc1_1 gpc1586 (
      {stage1_17[54]},
      {stage2_17[69]}
   );
   gpc1_1 gpc1587 (
      {stage1_17[55]},
      {stage2_17[70]}
   );
   gpc1_1 gpc1588 (
      {stage1_17[56]},
      {stage2_17[71]}
   );
   gpc1_1 gpc1589 (
      {stage1_17[57]},
      {stage2_17[72]}
   );
   gpc1_1 gpc1590 (
      {stage1_17[58]},
      {stage2_17[73]}
   );
   gpc1_1 gpc1591 (
      {stage1_17[59]},
      {stage2_17[74]}
   );
   gpc1_1 gpc1592 (
      {stage1_17[60]},
      {stage2_17[75]}
   );
   gpc1_1 gpc1593 (
      {stage1_17[61]},
      {stage2_17[76]}
   );
   gpc1_1 gpc1594 (
      {stage1_17[62]},
      {stage2_17[77]}
   );
   gpc1_1 gpc1595 (
      {stage1_17[63]},
      {stage2_17[78]}
   );
   gpc1_1 gpc1596 (
      {stage1_17[64]},
      {stage2_17[79]}
   );
   gpc1_1 gpc1597 (
      {stage1_17[65]},
      {stage2_17[80]}
   );
   gpc1_1 gpc1598 (
      {stage1_17[66]},
      {stage2_17[81]}
   );
   gpc1_1 gpc1599 (
      {stage1_17[67]},
      {stage2_17[82]}
   );
   gpc1_1 gpc1600 (
      {stage1_17[68]},
      {stage2_17[83]}
   );
   gpc1_1 gpc1601 (
      {stage1_17[69]},
      {stage2_17[84]}
   );
   gpc1_1 gpc1602 (
      {stage1_17[70]},
      {stage2_17[85]}
   );
   gpc1_1 gpc1603 (
      {stage1_17[71]},
      {stage2_17[86]}
   );
   gpc1_1 gpc1604 (
      {stage1_17[72]},
      {stage2_17[87]}
   );
   gpc1_1 gpc1605 (
      {stage1_17[73]},
      {stage2_17[88]}
   );
   gpc1_1 gpc1606 (
      {stage1_17[74]},
      {stage2_17[89]}
   );
   gpc1_1 gpc1607 (
      {stage1_17[75]},
      {stage2_17[90]}
   );
   gpc1_1 gpc1608 (
      {stage1_17[76]},
      {stage2_17[91]}
   );
   gpc1_1 gpc1609 (
      {stage1_17[77]},
      {stage2_17[92]}
   );
   gpc1_1 gpc1610 (
      {stage1_17[78]},
      {stage2_17[93]}
   );
   gpc1_1 gpc1611 (
      {stage1_17[79]},
      {stage2_17[94]}
   );
   gpc1_1 gpc1612 (
      {stage1_17[80]},
      {stage2_17[95]}
   );
   gpc1163_5 gpc1613 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc1614 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1163_5 gpc1615 (
      {stage2_0[6], stage2_0[7], stage2_0[8]},
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_2[2]},
      {stage2_3[2]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc1163_5 gpc1616 (
      {stage2_0[9], stage2_0[10], stage2_0[11]},
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_2[3]},
      {stage2_3[3]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc1617 (
      {stage2_0[12], stage2_0[13], stage2_0[14], stage2_0[15], stage2_0[16], stage2_0[17]},
      {stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc606_5 gpc1618 (
      {stage2_0[18], stage2_0[19], stage2_0[20], stage2_0[21], stage2_0[22], stage2_0[23]},
      {stage2_2[10], stage2_2[11], stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc606_5 gpc1619 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9]},
      {stage3_5[0],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc1620 (
      {stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34], stage2_1[35]},
      {stage2_3[10], stage2_3[11], stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15]},
      {stage3_5[1],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc1621 (
      {stage2_1[36], stage2_1[37], stage2_1[38], stage2_1[39], stage2_1[40], stage2_1[41]},
      {stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21]},
      {stage3_5[2],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc1622 (
      {stage2_1[42], stage2_1[43], stage2_1[44], stage2_1[45], stage2_1[46], stage2_1[47]},
      {stage2_3[22], stage2_3[23], stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27]},
      {stage3_5[3],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc606_5 gpc1623 (
      {stage2_1[48], stage2_1[49], stage2_1[50], stage2_1[51], stage2_1[52], stage2_1[53]},
      {stage2_3[28], stage2_3[29], stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33]},
      {stage3_5[4],stage3_4[10],stage3_3[10],stage3_2[10],stage3_1[10]}
   );
   gpc606_5 gpc1624 (
      {stage2_1[54], stage2_1[55], stage2_1[56], stage2_1[57], stage2_1[58], stage2_1[59]},
      {stage2_3[34], stage2_3[35], stage2_3[36], stage2_3[37], stage2_3[38], stage2_3[39]},
      {stage3_5[5],stage3_4[11],stage3_3[11],stage3_2[11],stage3_1[11]}
   );
   gpc606_5 gpc1625 (
      {stage2_2[16], stage2_2[17], stage2_2[18], stage2_2[19], stage2_2[20], stage2_2[21]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[6],stage3_4[12],stage3_3[12],stage3_2[12]}
   );
   gpc606_5 gpc1626 (
      {stage2_2[22], stage2_2[23], stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[7],stage3_4[13],stage3_3[13],stage3_2[13]}
   );
   gpc606_5 gpc1627 (
      {stage2_2[28], stage2_2[29], stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[8],stage3_4[14],stage3_3[14],stage3_2[14]}
   );
   gpc615_5 gpc1628 (
      {stage2_2[34], stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38]},
      {stage2_3[40]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[9],stage3_4[15],stage3_3[15],stage3_2[15]}
   );
   gpc615_5 gpc1629 (
      {stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43]},
      {stage2_3[41]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[10],stage3_4[16],stage3_3[16],stage3_2[16]}
   );
   gpc615_5 gpc1630 (
      {stage2_2[44], stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48]},
      {stage2_3[42]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[11],stage3_4[17],stage3_3[17],stage3_2[17]}
   );
   gpc615_5 gpc1631 (
      {stage2_2[49], stage2_2[50], stage2_2[51], stage2_2[52], stage2_2[53]},
      {stage2_3[43]},
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage3_6[6],stage3_5[12],stage3_4[18],stage3_3[18],stage3_2[18]}
   );
   gpc615_5 gpc1632 (
      {stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48]},
      {stage2_4[42]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[7],stage3_5[13],stage3_4[19],stage3_3[19]}
   );
   gpc615_5 gpc1633 (
      {stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52], stage2_3[53]},
      {stage2_4[43]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[8],stage3_5[14],stage3_4[20],stage3_3[20]}
   );
   gpc615_5 gpc1634 (
      {stage2_3[54], stage2_3[55], stage2_3[56], stage2_3[57], stage2_3[58]},
      {stage2_4[44]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[9],stage3_5[15],stage3_4[21],stage3_3[21]}
   );
   gpc615_5 gpc1635 (
      {stage2_3[59], stage2_3[60], stage2_3[61], stage2_3[62], stage2_3[63]},
      {stage2_4[45]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[10],stage3_5[16],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc1636 (
      {stage2_3[64], stage2_3[65], stage2_3[66], stage2_3[67], stage2_3[68]},
      {stage2_4[46]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[11],stage3_5[17],stage3_4[23],stage3_3[23]}
   );
   gpc606_5 gpc1637 (
      {stage2_4[47], stage2_4[48], stage2_4[49], stage2_4[50], stage2_4[51], stage2_4[52]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[5],stage3_6[12],stage3_5[18],stage3_4[24]}
   );
   gpc606_5 gpc1638 (
      {stage2_4[53], stage2_4[54], stage2_4[55], stage2_4[56], stage2_4[57], stage2_4[58]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[6],stage3_6[13],stage3_5[19],stage3_4[25]}
   );
   gpc606_5 gpc1639 (
      {stage2_4[59], stage2_4[60], stage2_4[61], stage2_4[62], stage2_4[63], stage2_4[64]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[7],stage3_6[14],stage3_5[20],stage3_4[26]}
   );
   gpc606_5 gpc1640 (
      {stage2_4[65], stage2_4[66], stage2_4[67], stage2_4[68], stage2_4[69], stage2_4[70]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[8],stage3_6[15],stage3_5[21],stage3_4[27]}
   );
   gpc606_5 gpc1641 (
      {stage2_4[71], stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75], stage2_4[76]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[9],stage3_6[16],stage3_5[22],stage3_4[28]}
   );
   gpc606_5 gpc1642 (
      {stage2_4[77], stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81], stage2_4[82]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[10],stage3_6[17],stage3_5[23],stage3_4[29]}
   );
   gpc606_5 gpc1643 (
      {stage2_4[83], stage2_4[84], stage2_4[85], stage2_4[86], stage2_4[87], stage2_4[88]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[11],stage3_6[18],stage3_5[24],stage3_4[30]}
   );
   gpc606_5 gpc1644 (
      {stage2_4[89], stage2_4[90], stage2_4[91], stage2_4[92], stage2_4[93], stage2_4[94]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[12],stage3_6[19],stage3_5[25],stage3_4[31]}
   );
   gpc606_5 gpc1645 (
      {stage2_4[95], stage2_4[96], stage2_4[97], stage2_4[98], stage2_4[99], stage2_4[100]},
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52], stage2_6[53]},
      {stage3_8[8],stage3_7[13],stage3_6[20],stage3_5[26],stage3_4[32]}
   );
   gpc606_5 gpc1646 (
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[9],stage3_7[14],stage3_6[21],stage3_5[27]}
   );
   gpc606_5 gpc1647 (
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[10],stage3_7[15],stage3_6[22],stage3_5[28]}
   );
   gpc606_5 gpc1648 (
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[11],stage3_7[16],stage3_6[23],stage3_5[29]}
   );
   gpc606_5 gpc1649 (
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[12],stage3_7[17],stage3_6[24],stage3_5[30]}
   );
   gpc606_5 gpc1650 (
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage3_9[4],stage3_8[13],stage3_7[18],stage3_6[25],stage3_5[31]}
   );
   gpc606_5 gpc1651 (
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64], stage2_5[65]},
      {stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35]},
      {stage3_9[5],stage3_8[14],stage3_7[19],stage3_6[26],stage3_5[32]}
   );
   gpc606_5 gpc1652 (
      {stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70], stage2_5[71]},
      {stage2_7[36], stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage3_9[6],stage3_8[15],stage3_7[20],stage3_6[27],stage3_5[33]}
   );
   gpc606_5 gpc1653 (
      {stage2_5[72], stage2_5[73], stage2_5[74], stage2_5[75], stage2_5[76], stage2_5[77]},
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46], stage2_7[47]},
      {stage3_9[7],stage3_8[16],stage3_7[21],stage3_6[28],stage3_5[34]}
   );
   gpc606_5 gpc1654 (
      {stage2_5[78], stage2_5[79], stage2_5[80], stage2_5[81], stage2_5[82], stage2_5[83]},
      {stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51], stage2_7[52], stage2_7[53]},
      {stage3_9[8],stage3_8[17],stage3_7[22],stage3_6[29],stage3_5[35]}
   );
   gpc606_5 gpc1655 (
      {stage2_5[84], stage2_5[85], stage2_5[86], stage2_5[87], stage2_5[88], stage2_5[89]},
      {stage2_7[54], stage2_7[55], stage2_7[56], stage2_7[57], stage2_7[58], stage2_7[59]},
      {stage3_9[9],stage3_8[18],stage3_7[23],stage3_6[30],stage3_5[36]}
   );
   gpc606_5 gpc1656 (
      {stage2_5[90], stage2_5[91], stage2_5[92], stage2_5[93], stage2_5[94], stage2_5[95]},
      {stage2_7[60], stage2_7[61], stage2_7[62], stage2_7[63], stage2_7[64], stage2_7[65]},
      {stage3_9[10],stage3_8[19],stage3_7[24],stage3_6[31],stage3_5[37]}
   );
   gpc606_5 gpc1657 (
      {stage2_5[96], stage2_5[97], stage2_5[98], stage2_5[99], stage2_5[100], stage2_5[101]},
      {stage2_7[66], stage2_7[67], stage2_7[68], stage2_7[69], stage2_7[70], stage2_7[71]},
      {stage3_9[11],stage3_8[20],stage3_7[25],stage3_6[32],stage3_5[38]}
   );
   gpc606_5 gpc1658 (
      {stage2_5[102], stage2_5[103], stage2_5[104], stage2_5[105], stage2_5[106], stage2_5[107]},
      {stage2_7[72], stage2_7[73], stage2_7[74], stage2_7[75], stage2_7[76], stage2_7[77]},
      {stage3_9[12],stage3_8[21],stage3_7[26],stage3_6[33],stage3_5[39]}
   );
   gpc615_5 gpc1659 (
      {stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57], stage2_6[58]},
      {stage2_7[78]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[13],stage3_8[22],stage3_7[27],stage3_6[34]}
   );
   gpc615_5 gpc1660 (
      {stage2_6[59], stage2_6[60], stage2_6[61], stage2_6[62], stage2_6[63]},
      {stage2_7[79]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[14],stage3_8[23],stage3_7[28],stage3_6[35]}
   );
   gpc615_5 gpc1661 (
      {stage2_6[64], stage2_6[65], stage2_6[66], stage2_6[67], stage2_6[68]},
      {stage2_7[80]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[15],stage3_8[24],stage3_7[29],stage3_6[36]}
   );
   gpc615_5 gpc1662 (
      {stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72], stage2_6[73]},
      {stage2_7[81]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[16],stage3_8[25],stage3_7[30],stage3_6[37]}
   );
   gpc615_5 gpc1663 (
      {stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77], stage2_6[78]},
      {stage2_7[82]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[17],stage3_8[26],stage3_7[31],stage3_6[38]}
   );
   gpc615_5 gpc1664 (
      {stage2_7[83], stage2_7[84], stage2_7[85], stage2_7[86], stage2_7[87]},
      {stage2_8[30]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[5],stage3_9[18],stage3_8[27],stage3_7[32]}
   );
   gpc615_5 gpc1665 (
      {stage2_7[88], stage2_7[89], stage2_7[90], stage2_7[91], stage2_7[92]},
      {stage2_8[31]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[6],stage3_9[19],stage3_8[28],stage3_7[33]}
   );
   gpc615_5 gpc1666 (
      {stage2_7[93], stage2_7[94], stage2_7[95], stage2_7[96], stage2_7[97]},
      {stage2_8[32]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[7],stage3_9[20],stage3_8[29],stage3_7[34]}
   );
   gpc615_5 gpc1667 (
      {stage2_7[98], stage2_7[99], stage2_7[100], stage2_7[101], stage2_7[102]},
      {stage2_8[33]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[8],stage3_9[21],stage3_8[30],stage3_7[35]}
   );
   gpc606_5 gpc1668 (
      {stage2_8[34], stage2_8[35], stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[9],stage3_9[22],stage3_8[31]}
   );
   gpc606_5 gpc1669 (
      {stage2_8[40], stage2_8[41], stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[10],stage3_9[23],stage3_8[32]}
   );
   gpc606_5 gpc1670 (
      {stage2_8[46], stage2_8[47], stage2_8[48], stage2_8[49], stage2_8[50], stage2_8[51]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[11],stage3_9[24],stage3_8[33]}
   );
   gpc606_5 gpc1671 (
      {stage2_8[52], stage2_8[53], stage2_8[54], stage2_8[55], stage2_8[56], stage2_8[57]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[7],stage3_10[12],stage3_9[25],stage3_8[34]}
   );
   gpc606_5 gpc1672 (
      {stage2_8[58], stage2_8[59], stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[8],stage3_10[13],stage3_9[26],stage3_8[35]}
   );
   gpc606_5 gpc1673 (
      {stage2_8[64], stage2_8[65], stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[9],stage3_10[14],stage3_9[27],stage3_8[36]}
   );
   gpc606_5 gpc1674 (
      {stage2_8[70], stage2_8[71], stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[6],stage3_11[10],stage3_10[15],stage3_9[28],stage3_8[37]}
   );
   gpc606_5 gpc1675 (
      {stage2_8[76], stage2_8[77], stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81]},
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage3_12[7],stage3_11[11],stage3_10[16],stage3_9[29],stage3_8[38]}
   );
   gpc606_5 gpc1676 (
      {stage2_8[82], stage2_8[83], stage2_8[84], stage2_8[85], stage2_8[86], stage2_8[87]},
      {stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53]},
      {stage3_12[8],stage3_11[12],stage3_10[17],stage3_9[30],stage3_8[39]}
   );
   gpc606_5 gpc1677 (
      {stage2_8[88], stage2_8[89], stage2_8[90], stage2_8[91], stage2_8[92], stage2_8[93]},
      {stage2_10[54], stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59]},
      {stage3_12[9],stage3_11[13],stage3_10[18],stage3_9[31],stage3_8[40]}
   );
   gpc606_5 gpc1678 (
      {stage2_8[94], stage2_8[95], stage2_8[96], stage2_8[97], stage2_8[98], stage2_8[99]},
      {stage2_10[60], stage2_10[61], stage2_10[62], stage2_10[63], stage2_10[64], stage2_10[65]},
      {stage3_12[10],stage3_11[14],stage3_10[19],stage3_9[32],stage3_8[41]}
   );
   gpc207_4 gpc1679 (
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29], stage2_9[30]},
      {stage2_11[0], stage2_11[1]},
      {stage3_12[11],stage3_11[15],stage3_10[20],stage3_9[33]}
   );
   gpc207_4 gpc1680 (
      {stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35], stage2_9[36], stage2_9[37]},
      {stage2_11[2], stage2_11[3]},
      {stage3_12[12],stage3_11[16],stage3_10[21],stage3_9[34]}
   );
   gpc606_5 gpc1681 (
      {stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41], stage2_9[42], stage2_9[43]},
      {stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9]},
      {stage3_13[0],stage3_12[13],stage3_11[17],stage3_10[22],stage3_9[35]}
   );
   gpc606_5 gpc1682 (
      {stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47], stage2_9[48], stage2_9[49]},
      {stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15]},
      {stage3_13[1],stage3_12[14],stage3_11[18],stage3_10[23],stage3_9[36]}
   );
   gpc606_5 gpc1683 (
      {stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53], stage2_9[54], stage2_9[55]},
      {stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21]},
      {stage3_13[2],stage3_12[15],stage3_11[19],stage3_10[24],stage3_9[37]}
   );
   gpc606_5 gpc1684 (
      {stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59], stage2_9[60], stage2_9[61]},
      {stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27]},
      {stage3_13[3],stage3_12[16],stage3_11[20],stage3_10[25],stage3_9[38]}
   );
   gpc606_5 gpc1685 (
      {stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65], stage2_9[66], stage2_9[67]},
      {stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33]},
      {stage3_13[4],stage3_12[17],stage3_11[21],stage3_10[26],stage3_9[39]}
   );
   gpc606_5 gpc1686 (
      {stage2_9[68], stage2_9[69], stage2_9[70], stage2_9[71], stage2_9[72], stage2_9[73]},
      {stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39]},
      {stage3_13[5],stage3_12[18],stage3_11[22],stage3_10[27],stage3_9[40]}
   );
   gpc606_5 gpc1687 (
      {stage2_9[74], stage2_9[75], stage2_9[76], stage2_9[77], stage2_9[78], stage2_9[79]},
      {stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45]},
      {stage3_13[6],stage3_12[19],stage3_11[23],stage3_10[28],stage3_9[41]}
   );
   gpc606_5 gpc1688 (
      {stage2_10[66], stage2_10[67], stage2_10[68], stage2_10[69], stage2_10[70], stage2_10[71]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[7],stage3_12[20],stage3_11[24],stage3_10[29]}
   );
   gpc615_5 gpc1689 (
      {stage2_10[72], stage2_10[73], stage2_10[74], stage2_10[75], stage2_10[76]},
      {stage2_11[46]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[8],stage3_12[21],stage3_11[25],stage3_10[30]}
   );
   gpc615_5 gpc1690 (
      {stage2_11[47], stage2_11[48], stage2_11[49], stage2_11[50], stage2_11[51]},
      {stage2_12[12]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[2],stage3_13[9],stage3_12[22],stage3_11[26]}
   );
   gpc615_5 gpc1691 (
      {stage2_11[52], stage2_11[53], stage2_11[54], stage2_11[55], stage2_11[56]},
      {stage2_12[13]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[3],stage3_13[10],stage3_12[23],stage3_11[27]}
   );
   gpc615_5 gpc1692 (
      {stage2_11[57], stage2_11[58], stage2_11[59], stage2_11[60], stage2_11[61]},
      {stage2_12[14]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[4],stage3_13[11],stage3_12[24],stage3_11[28]}
   );
   gpc615_5 gpc1693 (
      {stage2_11[62], stage2_11[63], stage2_11[64], stage2_11[65], stage2_11[66]},
      {stage2_12[15]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[5],stage3_13[12],stage3_12[25],stage3_11[29]}
   );
   gpc615_5 gpc1694 (
      {stage2_11[67], stage2_11[68], stage2_11[69], stage2_11[70], stage2_11[71]},
      {stage2_12[16]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[6],stage3_13[13],stage3_12[26],stage3_11[30]}
   );
   gpc615_5 gpc1695 (
      {stage2_11[72], stage2_11[73], stage2_11[74], stage2_11[75], stage2_11[76]},
      {stage2_12[17]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[7],stage3_13[14],stage3_12[27],stage3_11[31]}
   );
   gpc615_5 gpc1696 (
      {stage2_11[77], stage2_11[78], stage2_11[79], stage2_11[80], stage2_11[81]},
      {stage2_12[18]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[8],stage3_13[15],stage3_12[28],stage3_11[32]}
   );
   gpc615_5 gpc1697 (
      {stage2_11[82], stage2_11[83], stage2_11[84], stage2_11[85], stage2_11[86]},
      {stage2_12[19]},
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage3_15[7],stage3_14[9],stage3_13[16],stage3_12[29],stage3_11[33]}
   );
   gpc615_5 gpc1698 (
      {stage2_11[87], stage2_11[88], stage2_11[89], stage2_11[90], stage2_11[91]},
      {stage2_12[20]},
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage3_15[8],stage3_14[10],stage3_13[17],stage3_12[30],stage3_11[34]}
   );
   gpc615_5 gpc1699 (
      {stage2_11[92], stage2_11[93], stage2_11[94], stage2_11[95], stage2_11[96]},
      {stage2_12[21]},
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage3_15[9],stage3_14[11],stage3_13[18],stage3_12[31],stage3_11[35]}
   );
   gpc615_5 gpc1700 (
      {stage2_11[97], stage2_11[98], stage2_11[99], stage2_11[100], stage2_11[101]},
      {stage2_12[22]},
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage3_15[10],stage3_14[12],stage3_13[19],stage3_12[32],stage3_11[36]}
   );
   gpc615_5 gpc1701 (
      {stage2_11[102], stage2_11[103], stage2_11[104], stage2_11[105], stage2_11[106]},
      {stage2_12[23]},
      {stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69], stage2_13[70], stage2_13[71]},
      {stage3_15[11],stage3_14[13],stage3_13[20],stage3_12[33],stage3_11[37]}
   );
   gpc606_5 gpc1702 (
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[12],stage3_14[14],stage3_13[21],stage3_12[34]}
   );
   gpc606_5 gpc1703 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[13],stage3_14[15],stage3_13[22],stage3_12[35]}
   );
   gpc606_5 gpc1704 (
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[14],stage3_14[16],stage3_13[23],stage3_12[36]}
   );
   gpc606_5 gpc1705 (
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[15],stage3_14[17],stage3_13[24],stage3_12[37]}
   );
   gpc606_5 gpc1706 (
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[16],stage3_14[18],stage3_13[25],stage3_12[38]}
   );
   gpc615_5 gpc1707 (
      {stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58]},
      {stage2_13[72]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[17],stage3_14[19],stage3_13[26],stage3_12[39]}
   );
   gpc615_5 gpc1708 (
      {stage2_12[59], stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63]},
      {stage2_13[73]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[18],stage3_14[20],stage3_13[27],stage3_12[40]}
   );
   gpc615_5 gpc1709 (
      {stage2_12[64], stage2_12[65], stage2_12[66], stage2_12[67], stage2_12[68]},
      {stage2_13[74]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[19],stage3_14[21],stage3_13[28],stage3_12[41]}
   );
   gpc615_5 gpc1710 (
      {stage2_12[69], stage2_12[70], stage2_12[71], stage2_12[72], stage2_12[73]},
      {stage2_13[75]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[20],stage3_14[22],stage3_13[29],stage3_12[42]}
   );
   gpc615_5 gpc1711 (
      {stage2_12[74], stage2_12[75], stage2_12[76], stage2_12[77], stage2_12[78]},
      {stage2_13[76]},
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage3_16[9],stage3_15[21],stage3_14[23],stage3_13[30],stage3_12[43]}
   );
   gpc615_5 gpc1712 (
      {stage2_12[79], stage2_12[80], stage2_12[81], stage2_12[82], stage2_12[83]},
      {stage2_13[77]},
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage3_16[10],stage3_15[22],stage3_14[24],stage3_13[31],stage3_12[44]}
   );
   gpc615_5 gpc1713 (
      {stage2_12[84], stage2_12[85], stage2_12[86], stage2_12[87], stage2_12[88]},
      {stage2_13[78]},
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage3_16[11],stage3_15[23],stage3_14[25],stage3_13[32],stage3_12[45]}
   );
   gpc615_5 gpc1714 (
      {stage2_12[89], stage2_12[90], stage2_12[91], stage2_12[92], stage2_12[93]},
      {stage2_13[79]},
      {stage2_14[72], stage2_14[73], stage2_14[74], stage2_14[75], stage2_14[76], stage2_14[77]},
      {stage3_16[12],stage3_15[24],stage3_14[26],stage3_13[33],stage3_12[46]}
   );
   gpc615_5 gpc1715 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82]},
      {stage2_15[0]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[13],stage3_15[25],stage3_14[27]}
   );
   gpc615_5 gpc1716 (
      {stage2_14[83], stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87]},
      {stage2_15[1]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[14],stage3_15[26],stage3_14[28]}
   );
   gpc615_5 gpc1717 (
      {stage2_14[88], stage2_14[89], stage2_14[90], stage2_14[91], stage2_14[92]},
      {stage2_15[2]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[2],stage3_16[15],stage3_15[27],stage3_14[29]}
   );
   gpc615_5 gpc1718 (
      {stage2_14[93], stage2_14[94], stage2_14[95], stage2_14[96], stage2_14[97]},
      {stage2_15[3]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[3],stage3_16[16],stage3_15[28],stage3_14[30]}
   );
   gpc615_5 gpc1719 (
      {stage2_14[98], stage2_14[99], stage2_14[100], stage2_14[101], 1'b0},
      {stage2_15[4]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[4],stage3_16[17],stage3_15[29],stage3_14[31]}
   );
   gpc615_5 gpc1720 (
      {stage2_15[5], stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9]},
      {stage2_16[30]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[5],stage3_17[5],stage3_16[18],stage3_15[30]}
   );
   gpc615_5 gpc1721 (
      {stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13], stage2_15[14]},
      {stage2_16[31]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[6],stage3_17[6],stage3_16[19],stage3_15[31]}
   );
   gpc615_5 gpc1722 (
      {stage2_15[15], stage2_15[16], stage2_15[17], stage2_15[18], stage2_15[19]},
      {stage2_16[32]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[7],stage3_17[7],stage3_16[20],stage3_15[32]}
   );
   gpc615_5 gpc1723 (
      {stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23], stage2_15[24]},
      {stage2_16[33]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[8],stage3_17[8],stage3_16[21],stage3_15[33]}
   );
   gpc615_5 gpc1724 (
      {stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage2_16[34]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[9],stage3_17[9],stage3_16[22],stage3_15[34]}
   );
   gpc615_5 gpc1725 (
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34]},
      {stage2_16[35]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage3_19[5],stage3_18[10],stage3_17[10],stage3_16[23],stage3_15[35]}
   );
   gpc615_5 gpc1726 (
      {stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39]},
      {stage2_16[36]},
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage3_19[6],stage3_18[11],stage3_17[11],stage3_16[24],stage3_15[36]}
   );
   gpc615_5 gpc1727 (
      {stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44]},
      {stage2_16[37]},
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage3_19[7],stage3_18[12],stage3_17[12],stage3_16[25],stage3_15[37]}
   );
   gpc615_5 gpc1728 (
      {stage2_15[45], stage2_15[46], stage2_15[47], stage2_15[48], stage2_15[49]},
      {stage2_16[38]},
      {stage2_17[48], stage2_17[49], stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53]},
      {stage3_19[8],stage3_18[13],stage3_17[13],stage3_16[26],stage3_15[38]}
   );
   gpc615_5 gpc1729 (
      {stage2_15[50], stage2_15[51], stage2_15[52], stage2_15[53], stage2_15[54]},
      {stage2_16[39]},
      {stage2_17[54], stage2_17[55], stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59]},
      {stage3_19[9],stage3_18[14],stage3_17[14],stage3_16[27],stage3_15[39]}
   );
   gpc615_5 gpc1730 (
      {stage2_15[55], stage2_15[56], stage2_15[57], stage2_15[58], stage2_15[59]},
      {stage2_16[40]},
      {stage2_17[60], stage2_17[61], stage2_17[62], stage2_17[63], stage2_17[64], stage2_17[65]},
      {stage3_19[10],stage3_18[15],stage3_17[15],stage3_16[28],stage3_15[40]}
   );
   gpc615_5 gpc1731 (
      {stage2_15[60], stage2_15[61], stage2_15[62], stage2_15[63], stage2_15[64]},
      {stage2_16[41]},
      {stage2_17[66], stage2_17[67], stage2_17[68], stage2_17[69], stage2_17[70], stage2_17[71]},
      {stage3_19[11],stage3_18[16],stage3_17[16],stage3_16[29],stage3_15[41]}
   );
   gpc615_5 gpc1732 (
      {stage2_15[65], stage2_15[66], stage2_15[67], stage2_15[68], stage2_15[69]},
      {stage2_16[42]},
      {stage2_17[72], stage2_17[73], stage2_17[74], stage2_17[75], stage2_17[76], stage2_17[77]},
      {stage3_19[12],stage3_18[17],stage3_17[17],stage3_16[30],stage3_15[42]}
   );
   gpc615_5 gpc1733 (
      {stage2_15[70], stage2_15[71], stage2_15[72], stage2_15[73], stage2_15[74]},
      {stage2_16[43]},
      {stage2_17[78], stage2_17[79], stage2_17[80], stage2_17[81], stage2_17[82], stage2_17[83]},
      {stage3_19[13],stage3_18[18],stage3_17[18],stage3_16[31],stage3_15[43]}
   );
   gpc606_5 gpc1734 (
      {stage2_16[44], stage2_16[45], stage2_16[46], stage2_16[47], stage2_16[48], stage2_16[49]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[14],stage3_18[19],stage3_17[19],stage3_16[32]}
   );
   gpc606_5 gpc1735 (
      {stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53], stage2_16[54], stage2_16[55]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[15],stage3_18[20],stage3_17[20],stage3_16[33]}
   );
   gpc606_5 gpc1736 (
      {stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59], stage2_16[60], stage2_16[61]},
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage3_20[2],stage3_19[16],stage3_18[21],stage3_17[21],stage3_16[34]}
   );
   gpc606_5 gpc1737 (
      {stage2_16[62], stage2_16[63], stage2_16[64], stage2_16[65], stage2_16[66], stage2_16[67]},
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage3_20[3],stage3_19[17],stage3_18[22],stage3_17[22],stage3_16[35]}
   );
   gpc606_5 gpc1738 (
      {stage2_17[84], stage2_17[85], stage2_17[86], stage2_17[87], stage2_17[88], stage2_17[89]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], 1'b0},
      {stage3_21[0],stage3_20[4],stage3_19[18],stage3_18[23],stage3_17[23]}
   );
   gpc1_1 gpc1739 (
      {stage2_0[24]},
      {stage3_0[6]}
   );
   gpc1_1 gpc1740 (
      {stage2_0[25]},
      {stage3_0[7]}
   );
   gpc1_1 gpc1741 (
      {stage2_0[26]},
      {stage3_0[8]}
   );
   gpc1_1 gpc1742 (
      {stage2_0[27]},
      {stage3_0[9]}
   );
   gpc1_1 gpc1743 (
      {stage2_0[28]},
      {stage3_0[10]}
   );
   gpc1_1 gpc1744 (
      {stage2_0[29]},
      {stage3_0[11]}
   );
   gpc1_1 gpc1745 (
      {stage2_0[30]},
      {stage3_0[12]}
   );
   gpc1_1 gpc1746 (
      {stage2_0[31]},
      {stage3_0[13]}
   );
   gpc1_1 gpc1747 (
      {stage2_0[32]},
      {stage3_0[14]}
   );
   gpc1_1 gpc1748 (
      {stage2_0[33]},
      {stage3_0[15]}
   );
   gpc1_1 gpc1749 (
      {stage2_0[34]},
      {stage3_0[16]}
   );
   gpc1_1 gpc1750 (
      {stage2_0[35]},
      {stage3_0[17]}
   );
   gpc1_1 gpc1751 (
      {stage2_0[36]},
      {stage3_0[18]}
   );
   gpc1_1 gpc1752 (
      {stage2_0[37]},
      {stage3_0[19]}
   );
   gpc1_1 gpc1753 (
      {stage2_1[60]},
      {stage3_1[12]}
   );
   gpc1_1 gpc1754 (
      {stage2_1[61]},
      {stage3_1[13]}
   );
   gpc1_1 gpc1755 (
      {stage2_1[62]},
      {stage3_1[14]}
   );
   gpc1_1 gpc1756 (
      {stage2_3[69]},
      {stage3_3[24]}
   );
   gpc1_1 gpc1757 (
      {stage2_3[70]},
      {stage3_3[25]}
   );
   gpc1_1 gpc1758 (
      {stage2_3[71]},
      {stage3_3[26]}
   );
   gpc1_1 gpc1759 (
      {stage2_3[72]},
      {stage3_3[27]}
   );
   gpc1_1 gpc1760 (
      {stage2_3[73]},
      {stage3_3[28]}
   );
   gpc1_1 gpc1761 (
      {stage2_3[74]},
      {stage3_3[29]}
   );
   gpc1_1 gpc1762 (
      {stage2_3[75]},
      {stage3_3[30]}
   );
   gpc1_1 gpc1763 (
      {stage2_3[76]},
      {stage3_3[31]}
   );
   gpc1_1 gpc1764 (
      {stage2_3[77]},
      {stage3_3[32]}
   );
   gpc1_1 gpc1765 (
      {stage2_3[78]},
      {stage3_3[33]}
   );
   gpc1_1 gpc1766 (
      {stage2_3[79]},
      {stage3_3[34]}
   );
   gpc1_1 gpc1767 (
      {stage2_3[80]},
      {stage3_3[35]}
   );
   gpc1_1 gpc1768 (
      {stage2_3[81]},
      {stage3_3[36]}
   );
   gpc1_1 gpc1769 (
      {stage2_3[82]},
      {stage3_3[37]}
   );
   gpc1_1 gpc1770 (
      {stage2_3[83]},
      {stage3_3[38]}
   );
   gpc1_1 gpc1771 (
      {stage2_3[84]},
      {stage3_3[39]}
   );
   gpc1_1 gpc1772 (
      {stage2_3[85]},
      {stage3_3[40]}
   );
   gpc1_1 gpc1773 (
      {stage2_4[101]},
      {stage3_4[33]}
   );
   gpc1_1 gpc1774 (
      {stage2_4[102]},
      {stage3_4[34]}
   );
   gpc1_1 gpc1775 (
      {stage2_4[103]},
      {stage3_4[35]}
   );
   gpc1_1 gpc1776 (
      {stage2_4[104]},
      {stage3_4[36]}
   );
   gpc1_1 gpc1777 (
      {stage2_4[105]},
      {stage3_4[37]}
   );
   gpc1_1 gpc1778 (
      {stage2_4[106]},
      {stage3_4[38]}
   );
   gpc1_1 gpc1779 (
      {stage2_6[79]},
      {stage3_6[39]}
   );
   gpc1_1 gpc1780 (
      {stage2_6[80]},
      {stage3_6[40]}
   );
   gpc1_1 gpc1781 (
      {stage2_6[81]},
      {stage3_6[41]}
   );
   gpc1_1 gpc1782 (
      {stage2_6[82]},
      {stage3_6[42]}
   );
   gpc1_1 gpc1783 (
      {stage2_6[83]},
      {stage3_6[43]}
   );
   gpc1_1 gpc1784 (
      {stage2_6[84]},
      {stage3_6[44]}
   );
   gpc1_1 gpc1785 (
      {stage2_6[85]},
      {stage3_6[45]}
   );
   gpc1_1 gpc1786 (
      {stage2_6[86]},
      {stage3_6[46]}
   );
   gpc1_1 gpc1787 (
      {stage2_6[87]},
      {stage3_6[47]}
   );
   gpc1_1 gpc1788 (
      {stage2_6[88]},
      {stage3_6[48]}
   );
   gpc1_1 gpc1789 (
      {stage2_6[89]},
      {stage3_6[49]}
   );
   gpc1_1 gpc1790 (
      {stage2_8[100]},
      {stage3_8[42]}
   );
   gpc1_1 gpc1791 (
      {stage2_8[101]},
      {stage3_8[43]}
   );
   gpc1_1 gpc1792 (
      {stage2_8[102]},
      {stage3_8[44]}
   );
   gpc1_1 gpc1793 (
      {stage2_8[103]},
      {stage3_8[45]}
   );
   gpc1_1 gpc1794 (
      {stage2_8[104]},
      {stage3_8[46]}
   );
   gpc1_1 gpc1795 (
      {stage2_8[105]},
      {stage3_8[47]}
   );
   gpc1_1 gpc1796 (
      {stage2_9[80]},
      {stage3_9[42]}
   );
   gpc1_1 gpc1797 (
      {stage2_10[77]},
      {stage3_10[31]}
   );
   gpc1_1 gpc1798 (
      {stage2_10[78]},
      {stage3_10[32]}
   );
   gpc1_1 gpc1799 (
      {stage2_10[79]},
      {stage3_10[33]}
   );
   gpc1_1 gpc1800 (
      {stage2_10[80]},
      {stage3_10[34]}
   );
   gpc1_1 gpc1801 (
      {stage2_10[81]},
      {stage3_10[35]}
   );
   gpc1_1 gpc1802 (
      {stage2_10[82]},
      {stage3_10[36]}
   );
   gpc1_1 gpc1803 (
      {stage2_10[83]},
      {stage3_10[37]}
   );
   gpc1_1 gpc1804 (
      {stage2_10[84]},
      {stage3_10[38]}
   );
   gpc1_1 gpc1805 (
      {stage2_10[85]},
      {stage3_10[39]}
   );
   gpc1_1 gpc1806 (
      {stage2_10[86]},
      {stage3_10[40]}
   );
   gpc1_1 gpc1807 (
      {stage2_10[87]},
      {stage3_10[41]}
   );
   gpc1_1 gpc1808 (
      {stage2_10[88]},
      {stage3_10[42]}
   );
   gpc1_1 gpc1809 (
      {stage2_10[89]},
      {stage3_10[43]}
   );
   gpc1_1 gpc1810 (
      {stage2_13[80]},
      {stage3_13[34]}
   );
   gpc1_1 gpc1811 (
      {stage2_13[81]},
      {stage3_13[35]}
   );
   gpc1_1 gpc1812 (
      {stage2_13[82]},
      {stage3_13[36]}
   );
   gpc1_1 gpc1813 (
      {stage2_13[83]},
      {stage3_13[37]}
   );
   gpc1_1 gpc1814 (
      {stage2_13[84]},
      {stage3_13[38]}
   );
   gpc1_1 gpc1815 (
      {stage2_13[85]},
      {stage3_13[39]}
   );
   gpc1_1 gpc1816 (
      {stage2_16[68]},
      {stage3_16[36]}
   );
   gpc1_1 gpc1817 (
      {stage2_16[69]},
      {stage3_16[37]}
   );
   gpc1_1 gpc1818 (
      {stage2_16[70]},
      {stage3_16[38]}
   );
   gpc1_1 gpc1819 (
      {stage2_16[71]},
      {stage3_16[39]}
   );
   gpc1_1 gpc1820 (
      {stage2_16[72]},
      {stage3_16[40]}
   );
   gpc1_1 gpc1821 (
      {stage2_16[73]},
      {stage3_16[41]}
   );
   gpc1_1 gpc1822 (
      {stage2_16[74]},
      {stage3_16[42]}
   );
   gpc1_1 gpc1823 (
      {stage2_16[75]},
      {stage3_16[43]}
   );
   gpc1_1 gpc1824 (
      {stage2_16[76]},
      {stage3_16[44]}
   );
   gpc1_1 gpc1825 (
      {stage2_17[90]},
      {stage3_17[24]}
   );
   gpc1_1 gpc1826 (
      {stage2_17[91]},
      {stage3_17[25]}
   );
   gpc1_1 gpc1827 (
      {stage2_17[92]},
      {stage3_17[26]}
   );
   gpc1_1 gpc1828 (
      {stage2_17[93]},
      {stage3_17[27]}
   );
   gpc1_1 gpc1829 (
      {stage2_17[94]},
      {stage3_17[28]}
   );
   gpc1_1 gpc1830 (
      {stage2_17[95]},
      {stage3_17[29]}
   );
   gpc1_1 gpc1831 (
      {stage2_18[24]},
      {stage3_18[24]}
   );
   gpc1_1 gpc1832 (
      {stage2_18[25]},
      {stage3_18[25]}
   );
   gpc1406_5 gpc1833 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc1834 (
      {stage3_0[6], stage3_0[7], stage3_0[8], stage3_0[9], stage3_0[10], stage3_0[11]},
      {stage3_2[4], stage3_2[5], stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc1343_5 gpc1835 (
      {stage3_1[0], stage3_1[1], stage3_1[2]},
      {stage3_2[10], stage3_2[11], stage3_2[12], stage3_2[13]},
      {stage3_3[1], stage3_3[2], stage3_3[3]},
      {stage3_4[0]},
      {stage4_5[0],stage4_4[2],stage4_3[2],stage4_2[2],stage4_1[2]}
   );
   gpc606_5 gpc1836 (
      {stage3_1[3], stage3_1[4], stage3_1[5], stage3_1[6], stage3_1[7], stage3_1[8]},
      {stage3_3[4], stage3_3[5], stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9]},
      {stage4_5[1],stage4_4[3],stage4_3[3],stage4_2[3],stage4_1[3]}
   );
   gpc615_5 gpc1837 (
      {stage3_1[9], stage3_1[10], stage3_1[11], stage3_1[12], stage3_1[13]},
      {stage3_2[14]},
      {stage3_3[10], stage3_3[11], stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15]},
      {stage4_5[2],stage4_4[4],stage4_3[4],stage4_2[4],stage4_1[4]}
   );
   gpc615_5 gpc1838 (
      {stage3_3[16], stage3_3[17], stage3_3[18], stage3_3[19], stage3_3[20]},
      {stage3_4[1]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[0],stage4_5[3],stage4_4[5],stage4_3[5]}
   );
   gpc615_5 gpc1839 (
      {stage3_3[21], stage3_3[22], stage3_3[23], stage3_3[24], stage3_3[25]},
      {stage3_4[2]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[1],stage4_5[4],stage4_4[6],stage4_3[6]}
   );
   gpc615_5 gpc1840 (
      {stage3_3[26], stage3_3[27], stage3_3[28], stage3_3[29], stage3_3[30]},
      {stage3_4[3]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage4_7[2],stage4_6[2],stage4_5[5],stage4_4[7],stage4_3[7]}
   );
   gpc615_5 gpc1841 (
      {stage3_3[31], stage3_3[32], stage3_3[33], stage3_3[34], stage3_3[35]},
      {stage3_4[4]},
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage4_7[3],stage4_6[3],stage4_5[6],stage4_4[8],stage4_3[8]}
   );
   gpc615_5 gpc1842 (
      {stage3_3[36], stage3_3[37], stage3_3[38], stage3_3[39], stage3_3[40]},
      {stage3_4[5]},
      {stage3_5[24], stage3_5[25], stage3_5[26], stage3_5[27], stage3_5[28], stage3_5[29]},
      {stage4_7[4],stage4_6[4],stage4_5[7],stage4_4[9],stage4_3[9]}
   );
   gpc1415_5 gpc1843 (
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10]},
      {stage3_5[30]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[0]},
      {stage4_8[0],stage4_7[5],stage4_6[5],stage4_5[8],stage4_4[10]}
   );
   gpc606_5 gpc1844 (
      {stage3_4[11], stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16]},
      {stage3_6[4], stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage4_8[1],stage4_7[6],stage4_6[6],stage4_5[9],stage4_4[11]}
   );
   gpc606_5 gpc1845 (
      {stage3_4[17], stage3_4[18], stage3_4[19], stage3_4[20], stage3_4[21], stage3_4[22]},
      {stage3_6[10], stage3_6[11], stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15]},
      {stage4_8[2],stage4_7[7],stage4_6[7],stage4_5[10],stage4_4[12]}
   );
   gpc615_5 gpc1846 (
      {stage3_4[23], stage3_4[24], stage3_4[25], stage3_4[26], stage3_4[27]},
      {stage3_5[31]},
      {stage3_6[16], stage3_6[17], stage3_6[18], stage3_6[19], stage3_6[20], stage3_6[21]},
      {stage4_8[3],stage4_7[8],stage4_6[8],stage4_5[11],stage4_4[13]}
   );
   gpc615_5 gpc1847 (
      {stage3_4[28], stage3_4[29], stage3_4[30], stage3_4[31], stage3_4[32]},
      {stage3_5[32]},
      {stage3_6[22], stage3_6[23], stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27]},
      {stage4_8[4],stage4_7[9],stage4_6[9],stage4_5[12],stage4_4[14]}
   );
   gpc615_5 gpc1848 (
      {stage3_4[33], stage3_4[34], stage3_4[35], stage3_4[36], stage3_4[37]},
      {stage3_5[33]},
      {stage3_6[28], stage3_6[29], stage3_6[30], stage3_6[31], stage3_6[32], stage3_6[33]},
      {stage4_8[5],stage4_7[10],stage4_6[10],stage4_5[13],stage4_4[15]}
   );
   gpc606_5 gpc1849 (
      {stage3_5[34], stage3_5[35], stage3_5[36], stage3_5[37], stage3_5[38], stage3_5[39]},
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6]},
      {stage4_9[0],stage4_8[6],stage4_7[11],stage4_6[11],stage4_5[14]}
   );
   gpc615_5 gpc1850 (
      {stage3_6[34], stage3_6[35], stage3_6[36], stage3_6[37], stage3_6[38]},
      {stage3_7[7]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[1],stage4_8[7],stage4_7[12],stage4_6[12]}
   );
   gpc615_5 gpc1851 (
      {stage3_6[39], stage3_6[40], stage3_6[41], stage3_6[42], stage3_6[43]},
      {stage3_7[8]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[2],stage4_8[8],stage4_7[13],stage4_6[13]}
   );
   gpc615_5 gpc1852 (
      {stage3_6[44], stage3_6[45], stage3_6[46], stage3_6[47], stage3_6[48]},
      {stage3_7[9]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[3],stage4_8[9],stage4_7[14],stage4_6[14]}
   );
   gpc615_5 gpc1853 (
      {stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13], stage3_7[14]},
      {stage3_8[18]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[3],stage4_9[4],stage4_8[10],stage4_7[15]}
   );
   gpc615_5 gpc1854 (
      {stage3_7[15], stage3_7[16], stage3_7[17], stage3_7[18], stage3_7[19]},
      {stage3_8[19]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[4],stage4_9[5],stage4_8[11],stage4_7[16]}
   );
   gpc615_5 gpc1855 (
      {stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23], stage3_7[24]},
      {stage3_8[20]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[5],stage4_9[6],stage4_8[12],stage4_7[17]}
   );
   gpc615_5 gpc1856 (
      {stage3_7[25], stage3_7[26], stage3_7[27], stage3_7[28], stage3_7[29]},
      {stage3_8[21]},
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22], stage3_9[23]},
      {stage4_11[3],stage4_10[6],stage4_9[7],stage4_8[13],stage4_7[18]}
   );
   gpc615_5 gpc1857 (
      {stage3_7[30], stage3_7[31], stage3_7[32], stage3_7[33], stage3_7[34]},
      {stage3_8[22]},
      {stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27], stage3_9[28], stage3_9[29]},
      {stage4_11[4],stage4_10[7],stage4_9[8],stage4_8[14],stage4_7[19]}
   );
   gpc606_5 gpc1858 (
      {stage3_8[23], stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27], stage3_8[28]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[5],stage4_10[8],stage4_9[9],stage4_8[15]}
   );
   gpc606_5 gpc1859 (
      {stage3_8[29], stage3_8[30], stage3_8[31], stage3_8[32], stage3_8[33], stage3_8[34]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[6],stage4_10[9],stage4_9[10],stage4_8[16]}
   );
   gpc606_5 gpc1860 (
      {stage3_8[35], stage3_8[36], stage3_8[37], stage3_8[38], stage3_8[39], stage3_8[40]},
      {stage3_10[12], stage3_10[13], stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17]},
      {stage4_12[2],stage4_11[7],stage4_10[10],stage4_9[11],stage4_8[17]}
   );
   gpc606_5 gpc1861 (
      {stage3_8[41], stage3_8[42], stage3_8[43], stage3_8[44], stage3_8[45], stage3_8[46]},
      {stage3_10[18], stage3_10[19], stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23]},
      {stage4_12[3],stage4_11[8],stage4_10[11],stage4_9[12],stage4_8[18]}
   );
   gpc606_5 gpc1862 (
      {stage3_9[30], stage3_9[31], stage3_9[32], stage3_9[33], stage3_9[34], stage3_9[35]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[4],stage4_11[9],stage4_10[12],stage4_9[13]}
   );
   gpc606_5 gpc1863 (
      {stage3_9[36], stage3_9[37], stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[5],stage4_11[10],stage4_10[13],stage4_9[14]}
   );
   gpc615_5 gpc1864 (
      {stage3_10[24], stage3_10[25], stage3_10[26], stage3_10[27], stage3_10[28]},
      {stage3_11[12]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[2],stage4_12[6],stage4_11[11],stage4_10[14]}
   );
   gpc615_5 gpc1865 (
      {stage3_10[29], stage3_10[30], stage3_10[31], stage3_10[32], stage3_10[33]},
      {stage3_11[13]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[3],stage4_12[7],stage4_11[12],stage4_10[15]}
   );
   gpc615_5 gpc1866 (
      {stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37], stage3_10[38]},
      {stage3_11[14]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[4],stage4_12[8],stage4_11[13],stage4_10[16]}
   );
   gpc615_5 gpc1867 (
      {stage3_10[39], stage3_10[40], stage3_10[41], stage3_10[42], stage3_10[43]},
      {stage3_11[15]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage4_14[3],stage4_13[5],stage4_12[9],stage4_11[14],stage4_10[17]}
   );
   gpc606_5 gpc1868 (
      {stage3_11[16], stage3_11[17], stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[4],stage4_13[6],stage4_12[10],stage4_11[15]}
   );
   gpc606_5 gpc1869 (
      {stage3_11[22], stage3_11[23], stage3_11[24], stage3_11[25], stage3_11[26], stage3_11[27]},
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage4_15[1],stage4_14[5],stage4_13[7],stage4_12[11],stage4_11[16]}
   );
   gpc615_5 gpc1870 (
      {stage3_11[28], stage3_11[29], stage3_11[30], stage3_11[31], stage3_11[32]},
      {stage3_12[24]},
      {stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage4_15[2],stage4_14[6],stage4_13[8],stage4_12[12],stage4_11[17]}
   );
   gpc615_5 gpc1871 (
      {stage3_11[33], stage3_11[34], stage3_11[35], stage3_11[36], stage3_11[37]},
      {stage3_12[25]},
      {stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23]},
      {stage4_15[3],stage4_14[7],stage4_13[9],stage4_12[13],stage4_11[18]}
   );
   gpc117_4 gpc1872 (
      {stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29], stage3_12[30], stage3_12[31], stage3_12[32]},
      {stage3_13[24]},
      {stage3_14[0]},
      {stage4_15[4],stage4_14[8],stage4_13[10],stage4_12[14]}
   );
   gpc606_5 gpc1873 (
      {stage3_12[33], stage3_12[34], stage3_12[35], stage3_12[36], stage3_12[37], stage3_12[38]},
      {stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6]},
      {stage4_16[0],stage4_15[5],stage4_14[9],stage4_13[11],stage4_12[15]}
   );
   gpc606_5 gpc1874 (
      {stage3_13[25], stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29], stage3_13[30]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[6],stage4_14[10],stage4_13[12]}
   );
   gpc606_5 gpc1875 (
      {stage3_13[31], stage3_13[32], stage3_13[33], stage3_13[34], stage3_13[35], stage3_13[36]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[2],stage4_15[7],stage4_14[11],stage4_13[13]}
   );
   gpc606_5 gpc1876 (
      {stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11], stage3_14[12]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[2],stage4_16[3],stage4_15[8],stage4_14[12]}
   );
   gpc615_5 gpc1877 (
      {stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17]},
      {stage3_15[12]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[3],stage4_16[4],stage4_15[9],stage4_14[13]}
   );
   gpc615_5 gpc1878 (
      {stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22]},
      {stage3_15[13]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[4],stage4_16[5],stage4_15[10],stage4_14[14]}
   );
   gpc615_5 gpc1879 (
      {stage3_14[23], stage3_14[24], stage3_14[25], stage3_14[26], stage3_14[27]},
      {stage3_15[14]},
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23]},
      {stage4_18[3],stage4_17[5],stage4_16[6],stage4_15[11],stage4_14[15]}
   );
   gpc606_5 gpc1880 (
      {stage3_15[15], stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19], stage3_15[20]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[4],stage4_17[6],stage4_16[7],stage4_15[12]}
   );
   gpc615_5 gpc1881 (
      {stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25]},
      {stage3_16[24]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[5],stage4_17[7],stage4_16[8],stage4_15[13]}
   );
   gpc615_5 gpc1882 (
      {stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29], stage3_15[30]},
      {stage3_16[25]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[6],stage4_17[8],stage4_16[9],stage4_15[14]}
   );
   gpc606_5 gpc1883 (
      {stage3_16[26], stage3_16[27], stage3_16[28], stage3_16[29], stage3_16[30], stage3_16[31]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[3],stage4_18[7],stage4_17[9],stage4_16[10]}
   );
   gpc606_5 gpc1884 (
      {stage3_16[32], stage3_16[33], stage3_16[34], stage3_16[35], stage3_16[36], stage3_16[37]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[4],stage4_18[8],stage4_17[10],stage4_16[11]}
   );
   gpc606_5 gpc1885 (
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[2],stage4_19[5],stage4_18[9],stage4_17[11]}
   );
   gpc606_5 gpc1886 (
      {stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[3],stage4_19[6],stage4_18[10],stage4_17[12]}
   );
   gpc1_1 gpc1887 (
      {stage3_0[12]},
      {stage4_0[2]}
   );
   gpc1_1 gpc1888 (
      {stage3_0[13]},
      {stage4_0[3]}
   );
   gpc1_1 gpc1889 (
      {stage3_0[14]},
      {stage4_0[4]}
   );
   gpc1_1 gpc1890 (
      {stage3_0[15]},
      {stage4_0[5]}
   );
   gpc1_1 gpc1891 (
      {stage3_0[16]},
      {stage4_0[6]}
   );
   gpc1_1 gpc1892 (
      {stage3_0[17]},
      {stage4_0[7]}
   );
   gpc1_1 gpc1893 (
      {stage3_0[18]},
      {stage4_0[8]}
   );
   gpc1_1 gpc1894 (
      {stage3_0[19]},
      {stage4_0[9]}
   );
   gpc1_1 gpc1895 (
      {stage3_1[14]},
      {stage4_1[5]}
   );
   gpc1_1 gpc1896 (
      {stage3_2[15]},
      {stage4_2[5]}
   );
   gpc1_1 gpc1897 (
      {stage3_2[16]},
      {stage4_2[6]}
   );
   gpc1_1 gpc1898 (
      {stage3_2[17]},
      {stage4_2[7]}
   );
   gpc1_1 gpc1899 (
      {stage3_2[18]},
      {stage4_2[8]}
   );
   gpc1_1 gpc1900 (
      {stage3_4[38]},
      {stage4_4[16]}
   );
   gpc1_1 gpc1901 (
      {stage3_6[49]},
      {stage4_6[15]}
   );
   gpc1_1 gpc1902 (
      {stage3_7[35]},
      {stage4_7[20]}
   );
   gpc1_1 gpc1903 (
      {stage3_8[47]},
      {stage4_8[19]}
   );
   gpc1_1 gpc1904 (
      {stage3_9[42]},
      {stage4_9[15]}
   );
   gpc1_1 gpc1905 (
      {stage3_12[39]},
      {stage4_12[16]}
   );
   gpc1_1 gpc1906 (
      {stage3_12[40]},
      {stage4_12[17]}
   );
   gpc1_1 gpc1907 (
      {stage3_12[41]},
      {stage4_12[18]}
   );
   gpc1_1 gpc1908 (
      {stage3_12[42]},
      {stage4_12[19]}
   );
   gpc1_1 gpc1909 (
      {stage3_12[43]},
      {stage4_12[20]}
   );
   gpc1_1 gpc1910 (
      {stage3_12[44]},
      {stage4_12[21]}
   );
   gpc1_1 gpc1911 (
      {stage3_12[45]},
      {stage4_12[22]}
   );
   gpc1_1 gpc1912 (
      {stage3_12[46]},
      {stage4_12[23]}
   );
   gpc1_1 gpc1913 (
      {stage3_13[37]},
      {stage4_13[14]}
   );
   gpc1_1 gpc1914 (
      {stage3_13[38]},
      {stage4_13[15]}
   );
   gpc1_1 gpc1915 (
      {stage3_13[39]},
      {stage4_13[16]}
   );
   gpc1_1 gpc1916 (
      {stage3_14[28]},
      {stage4_14[16]}
   );
   gpc1_1 gpc1917 (
      {stage3_14[29]},
      {stage4_14[17]}
   );
   gpc1_1 gpc1918 (
      {stage3_14[30]},
      {stage4_14[18]}
   );
   gpc1_1 gpc1919 (
      {stage3_14[31]},
      {stage4_14[19]}
   );
   gpc1_1 gpc1920 (
      {stage3_15[31]},
      {stage4_15[15]}
   );
   gpc1_1 gpc1921 (
      {stage3_15[32]},
      {stage4_15[16]}
   );
   gpc1_1 gpc1922 (
      {stage3_15[33]},
      {stage4_15[17]}
   );
   gpc1_1 gpc1923 (
      {stage3_15[34]},
      {stage4_15[18]}
   );
   gpc1_1 gpc1924 (
      {stage3_15[35]},
      {stage4_15[19]}
   );
   gpc1_1 gpc1925 (
      {stage3_15[36]},
      {stage4_15[20]}
   );
   gpc1_1 gpc1926 (
      {stage3_15[37]},
      {stage4_15[21]}
   );
   gpc1_1 gpc1927 (
      {stage3_15[38]},
      {stage4_15[22]}
   );
   gpc1_1 gpc1928 (
      {stage3_15[39]},
      {stage4_15[23]}
   );
   gpc1_1 gpc1929 (
      {stage3_15[40]},
      {stage4_15[24]}
   );
   gpc1_1 gpc1930 (
      {stage3_15[41]},
      {stage4_15[25]}
   );
   gpc1_1 gpc1931 (
      {stage3_15[42]},
      {stage4_15[26]}
   );
   gpc1_1 gpc1932 (
      {stage3_15[43]},
      {stage4_15[27]}
   );
   gpc1_1 gpc1933 (
      {stage3_16[38]},
      {stage4_16[12]}
   );
   gpc1_1 gpc1934 (
      {stage3_16[39]},
      {stage4_16[13]}
   );
   gpc1_1 gpc1935 (
      {stage3_16[40]},
      {stage4_16[14]}
   );
   gpc1_1 gpc1936 (
      {stage3_16[41]},
      {stage4_16[15]}
   );
   gpc1_1 gpc1937 (
      {stage3_16[42]},
      {stage4_16[16]}
   );
   gpc1_1 gpc1938 (
      {stage3_16[43]},
      {stage4_16[17]}
   );
   gpc1_1 gpc1939 (
      {stage3_16[44]},
      {stage4_16[18]}
   );
   gpc1_1 gpc1940 (
      {stage3_18[12]},
      {stage4_18[11]}
   );
   gpc1_1 gpc1941 (
      {stage3_18[13]},
      {stage4_18[12]}
   );
   gpc1_1 gpc1942 (
      {stage3_18[14]},
      {stage4_18[13]}
   );
   gpc1_1 gpc1943 (
      {stage3_18[15]},
      {stage4_18[14]}
   );
   gpc1_1 gpc1944 (
      {stage3_18[16]},
      {stage4_18[15]}
   );
   gpc1_1 gpc1945 (
      {stage3_18[17]},
      {stage4_18[16]}
   );
   gpc1_1 gpc1946 (
      {stage3_18[18]},
      {stage4_18[17]}
   );
   gpc1_1 gpc1947 (
      {stage3_18[19]},
      {stage4_18[18]}
   );
   gpc1_1 gpc1948 (
      {stage3_18[20]},
      {stage4_18[19]}
   );
   gpc1_1 gpc1949 (
      {stage3_18[21]},
      {stage4_18[20]}
   );
   gpc1_1 gpc1950 (
      {stage3_18[22]},
      {stage4_18[21]}
   );
   gpc1_1 gpc1951 (
      {stage3_18[23]},
      {stage4_18[22]}
   );
   gpc1_1 gpc1952 (
      {stage3_18[24]},
      {stage4_18[23]}
   );
   gpc1_1 gpc1953 (
      {stage3_18[25]},
      {stage4_18[24]}
   );
   gpc1_1 gpc1954 (
      {stage3_19[12]},
      {stage4_19[7]}
   );
   gpc1_1 gpc1955 (
      {stage3_19[13]},
      {stage4_19[8]}
   );
   gpc1_1 gpc1956 (
      {stage3_19[14]},
      {stage4_19[9]}
   );
   gpc1_1 gpc1957 (
      {stage3_19[15]},
      {stage4_19[10]}
   );
   gpc1_1 gpc1958 (
      {stage3_19[16]},
      {stage4_19[11]}
   );
   gpc1_1 gpc1959 (
      {stage3_19[17]},
      {stage4_19[12]}
   );
   gpc1_1 gpc1960 (
      {stage3_19[18]},
      {stage4_19[13]}
   );
   gpc1_1 gpc1961 (
      {stage3_20[0]},
      {stage4_20[4]}
   );
   gpc1_1 gpc1962 (
      {stage3_20[1]},
      {stage4_20[5]}
   );
   gpc1_1 gpc1963 (
      {stage3_20[2]},
      {stage4_20[6]}
   );
   gpc1_1 gpc1964 (
      {stage3_20[3]},
      {stage4_20[7]}
   );
   gpc1_1 gpc1965 (
      {stage3_20[4]},
      {stage4_20[8]}
   );
   gpc1_1 gpc1966 (
      {stage3_21[0]},
      {stage4_21[2]}
   );
   gpc615_5 gpc1967 (
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4]},
      {stage4_4[0]},
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0]}
   );
   gpc2135_5 gpc1968 (
      {stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_5[6], stage4_5[7], stage4_5[8]},
      {stage4_6[0]},
      {stage4_7[0], stage4_7[1]},
      {stage5_8[0],stage5_7[1],stage5_6[1],stage5_5[1],stage5_4[1]}
   );
   gpc2135_5 gpc1969 (
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10]},
      {stage4_5[9], stage4_5[10], stage4_5[11]},
      {stage4_6[1]},
      {stage4_7[2], stage4_7[3]},
      {stage5_8[1],stage5_7[2],stage5_6[2],stage5_5[2],stage5_4[2]}
   );
   gpc2135_5 gpc1970 (
      {stage4_4[11], stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15]},
      {stage4_5[12], stage4_5[13], stage4_5[14]},
      {stage4_6[2]},
      {stage4_7[4], stage4_7[5]},
      {stage5_8[2],stage5_7[3],stage5_6[3],stage5_5[3],stage5_4[3]}
   );
   gpc615_5 gpc1971 (
      {stage4_6[3], stage4_6[4], stage4_6[5], stage4_6[6], stage4_6[7]},
      {stage4_7[6]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[0],stage5_8[3],stage5_7[4],stage5_6[4]}
   );
   gpc615_5 gpc1972 (
      {stage4_6[8], stage4_6[9], stage4_6[10], stage4_6[11], stage4_6[12]},
      {stage4_7[7]},
      {stage4_8[6], stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11]},
      {stage5_10[1],stage5_9[1],stage5_8[4],stage5_7[5],stage5_6[5]}
   );
   gpc2116_5 gpc1973 (
      {stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11], stage4_7[12], stage4_7[13]},
      {stage4_8[12]},
      {stage4_9[0]},
      {stage4_10[0], stage4_10[1]},
      {stage5_11[0],stage5_10[2],stage5_9[2],stage5_8[5],stage5_7[6]}
   );
   gpc606_5 gpc1974 (
      {stage4_7[14], stage4_7[15], stage4_7[16], stage4_7[17], stage4_7[18], stage4_7[19]},
      {stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6]},
      {stage5_11[1],stage5_10[3],stage5_9[3],stage5_8[6],stage5_7[7]}
   );
   gpc623_5 gpc1975 (
      {stage4_9[7], stage4_9[8], stage4_9[9]},
      {stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[0],stage5_11[2],stage5_10[4],stage5_9[4]}
   );
   gpc623_5 gpc1976 (
      {stage4_9[10], stage4_9[11], stage4_9[12]},
      {stage4_10[4], stage4_10[5]},
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage5_13[1],stage5_12[1],stage5_11[3],stage5_10[5],stage5_9[5]}
   );
   gpc606_5 gpc1977 (
      {stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[2],stage5_12[2],stage5_11[4],stage5_10[6]}
   );
   gpc606_5 gpc1978 (
      {stage4_10[12], stage4_10[13], stage4_10[14], stage4_10[15], stage4_10[16], stage4_10[17]},
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage5_14[1],stage5_13[3],stage5_12[3],stage5_11[5],stage5_10[7]}
   );
   gpc7_3 gpc1979 (
      {stage4_11[12], stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16], stage4_11[17], stage4_11[18]},
      {stage5_13[4],stage5_12[4],stage5_11[6]}
   );
   gpc606_5 gpc1980 (
      {stage4_12[12], stage4_12[13], stage4_12[14], stage4_12[15], stage4_12[16], stage4_12[17]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[2],stage5_13[5],stage5_12[5]}
   );
   gpc606_5 gpc1981 (
      {stage4_12[18], stage4_12[19], stage4_12[20], stage4_12[21], stage4_12[22], stage4_12[23]},
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10], stage4_14[11]},
      {stage5_16[1],stage5_15[1],stage5_14[3],stage5_13[6],stage5_12[6]}
   );
   gpc606_5 gpc1982 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[2],stage5_15[2],stage5_14[4],stage5_13[7]}
   );
   gpc606_5 gpc1983 (
      {stage4_13[6], stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11]},
      {stage4_15[6], stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage5_17[1],stage5_16[3],stage5_15[3],stage5_14[5],stage5_13[8]}
   );
   gpc615_5 gpc1984 (
      {stage4_13[12], stage4_13[13], stage4_13[14], stage4_13[15], stage4_13[16]},
      {stage4_14[12]},
      {stage4_15[12], stage4_15[13], stage4_15[14], stage4_15[15], stage4_15[16], stage4_15[17]},
      {stage5_17[2],stage5_16[4],stage5_15[4],stage5_14[6],stage5_13[9]}
   );
   gpc7_3 gpc1985 (
      {stage4_14[13], stage4_14[14], stage4_14[15], stage4_14[16], stage4_14[17], stage4_14[18], stage4_14[19]},
      {stage5_16[5],stage5_15[5],stage5_14[7]}
   );
   gpc1163_5 gpc1986 (
      {stage4_15[18], stage4_15[19], stage4_15[20]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage4_17[0]},
      {stage4_18[0]},
      {stage5_19[0],stage5_18[0],stage5_17[3],stage5_16[6],stage5_15[6]}
   );
   gpc615_5 gpc1987 (
      {stage4_15[21], stage4_15[22], stage4_15[23], stage4_15[24], stage4_15[25]},
      {stage4_16[6]},
      {stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5], stage4_17[6]},
      {stage5_19[1],stage5_18[1],stage5_17[4],stage5_16[7],stage5_15[7]}
   );
   gpc606_5 gpc1988 (
      {stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11], stage4_16[12]},
      {stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6]},
      {stage5_20[0],stage5_19[2],stage5_18[2],stage5_17[5],stage5_16[8]}
   );
   gpc606_5 gpc1989 (
      {stage4_16[13], stage4_16[14], stage4_16[15], stage4_16[16], stage4_16[17], stage4_16[18]},
      {stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11], stage4_18[12]},
      {stage5_20[1],stage5_19[3],stage5_18[3],stage5_17[6],stage5_16[9]}
   );
   gpc606_5 gpc1990 (
      {stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11], stage4_17[12]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[2],stage5_19[4],stage5_18[4],stage5_17[7]}
   );
   gpc2135_5 gpc1991 (
      {stage4_18[13], stage4_18[14], stage4_18[15], stage4_18[16], stage4_18[17]},
      {stage4_19[6], stage4_19[7], stage4_19[8]},
      {stage4_20[0]},
      {stage4_21[0], stage4_21[1]},
      {stage5_22[0],stage5_21[1],stage5_20[3],stage5_19[5],stage5_18[5]}
   );
   gpc117_4 gpc1992 (
      {stage4_18[18], stage4_18[19], stage4_18[20], stage4_18[21], stage4_18[22], stage4_18[23], stage4_18[24]},
      {stage4_19[9]},
      {stage4_20[1]},
      {stage5_21[2],stage5_20[4],stage5_19[6],stage5_18[6]}
   );
   gpc1_1 gpc1993 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1994 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1995 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc1996 (
      {stage4_0[3]},
      {stage5_0[3]}
   );
   gpc1_1 gpc1997 (
      {stage4_0[4]},
      {stage5_0[4]}
   );
   gpc1_1 gpc1998 (
      {stage4_0[5]},
      {stage5_0[5]}
   );
   gpc1_1 gpc1999 (
      {stage4_0[6]},
      {stage5_0[6]}
   );
   gpc1_1 gpc2000 (
      {stage4_0[7]},
      {stage5_0[7]}
   );
   gpc1_1 gpc2001 (
      {stage4_0[8]},
      {stage5_0[8]}
   );
   gpc1_1 gpc2002 (
      {stage4_0[9]},
      {stage5_0[9]}
   );
   gpc1_1 gpc2003 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc2004 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc2005 (
      {stage4_1[2]},
      {stage5_1[2]}
   );
   gpc1_1 gpc2006 (
      {stage4_1[3]},
      {stage5_1[3]}
   );
   gpc1_1 gpc2007 (
      {stage4_1[4]},
      {stage5_1[4]}
   );
   gpc1_1 gpc2008 (
      {stage4_1[5]},
      {stage5_1[5]}
   );
   gpc1_1 gpc2009 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc2010 (
      {stage4_2[1]},
      {stage5_2[1]}
   );
   gpc1_1 gpc2011 (
      {stage4_2[2]},
      {stage5_2[2]}
   );
   gpc1_1 gpc2012 (
      {stage4_2[3]},
      {stage5_2[3]}
   );
   gpc1_1 gpc2013 (
      {stage4_2[4]},
      {stage5_2[4]}
   );
   gpc1_1 gpc2014 (
      {stage4_2[5]},
      {stage5_2[5]}
   );
   gpc1_1 gpc2015 (
      {stage4_2[6]},
      {stage5_2[6]}
   );
   gpc1_1 gpc2016 (
      {stage4_2[7]},
      {stage5_2[7]}
   );
   gpc1_1 gpc2017 (
      {stage4_2[8]},
      {stage5_2[8]}
   );
   gpc1_1 gpc2018 (
      {stage4_3[5]},
      {stage5_3[1]}
   );
   gpc1_1 gpc2019 (
      {stage4_3[6]},
      {stage5_3[2]}
   );
   gpc1_1 gpc2020 (
      {stage4_3[7]},
      {stage5_3[3]}
   );
   gpc1_1 gpc2021 (
      {stage4_3[8]},
      {stage5_3[4]}
   );
   gpc1_1 gpc2022 (
      {stage4_3[9]},
      {stage5_3[5]}
   );
   gpc1_1 gpc2023 (
      {stage4_4[16]},
      {stage5_4[4]}
   );
   gpc1_1 gpc2024 (
      {stage4_6[13]},
      {stage5_6[6]}
   );
   gpc1_1 gpc2025 (
      {stage4_6[14]},
      {stage5_6[7]}
   );
   gpc1_1 gpc2026 (
      {stage4_6[15]},
      {stage5_6[8]}
   );
   gpc1_1 gpc2027 (
      {stage4_7[20]},
      {stage5_7[8]}
   );
   gpc1_1 gpc2028 (
      {stage4_8[13]},
      {stage5_8[7]}
   );
   gpc1_1 gpc2029 (
      {stage4_8[14]},
      {stage5_8[8]}
   );
   gpc1_1 gpc2030 (
      {stage4_8[15]},
      {stage5_8[9]}
   );
   gpc1_1 gpc2031 (
      {stage4_8[16]},
      {stage5_8[10]}
   );
   gpc1_1 gpc2032 (
      {stage4_8[17]},
      {stage5_8[11]}
   );
   gpc1_1 gpc2033 (
      {stage4_8[18]},
      {stage5_8[12]}
   );
   gpc1_1 gpc2034 (
      {stage4_8[19]},
      {stage5_8[13]}
   );
   gpc1_1 gpc2035 (
      {stage4_9[13]},
      {stage5_9[6]}
   );
   gpc1_1 gpc2036 (
      {stage4_9[14]},
      {stage5_9[7]}
   );
   gpc1_1 gpc2037 (
      {stage4_9[15]},
      {stage5_9[8]}
   );
   gpc1_1 gpc2038 (
      {stage4_15[26]},
      {stage5_15[8]}
   );
   gpc1_1 gpc2039 (
      {stage4_15[27]},
      {stage5_15[9]}
   );
   gpc1_1 gpc2040 (
      {stage4_19[10]},
      {stage5_19[7]}
   );
   gpc1_1 gpc2041 (
      {stage4_19[11]},
      {stage5_19[8]}
   );
   gpc1_1 gpc2042 (
      {stage4_19[12]},
      {stage5_19[9]}
   );
   gpc1_1 gpc2043 (
      {stage4_19[13]},
      {stage5_19[10]}
   );
   gpc1_1 gpc2044 (
      {stage4_20[2]},
      {stage5_20[5]}
   );
   gpc1_1 gpc2045 (
      {stage4_20[3]},
      {stage5_20[6]}
   );
   gpc1_1 gpc2046 (
      {stage4_20[4]},
      {stage5_20[7]}
   );
   gpc1_1 gpc2047 (
      {stage4_20[5]},
      {stage5_20[8]}
   );
   gpc1_1 gpc2048 (
      {stage4_20[6]},
      {stage5_20[9]}
   );
   gpc1_1 gpc2049 (
      {stage4_20[7]},
      {stage5_20[10]}
   );
   gpc1_1 gpc2050 (
      {stage4_20[8]},
      {stage5_20[11]}
   );
   gpc1_1 gpc2051 (
      {stage4_21[2]},
      {stage5_21[3]}
   );
   gpc2135_5 gpc2052 (
      {stage5_0[0], stage5_0[1], stage5_0[2], stage5_0[3], stage5_0[4]},
      {stage5_1[0], stage5_1[1], stage5_1[2]},
      {stage5_2[0]},
      {stage5_3[0], stage5_3[1]},
      {stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc135_4 gpc2053 (
      {stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4], stage5_2[5]},
      {stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0]},
      {stage6_5[0],stage6_4[1],stage6_3[1],stage6_2[1]}
   );
   gpc615_5 gpc2054 (
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4]},
      {stage5_7[0]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[0],stage6_6[0]}
   );
   gpc623_5 gpc2055 (
      {stage5_6[5], stage5_6[6], stage5_6[7]},
      {stage5_7[1], stage5_7[2]},
      {stage5_8[6], stage5_8[7], stage5_8[8], stage5_8[9], stage5_8[10], stage5_8[11]},
      {stage6_10[1],stage6_9[1],stage6_8[1],stage6_7[1],stage6_6[1]}
   );
   gpc615_5 gpc2056 (
      {stage5_7[3], stage5_7[4], stage5_7[5], stage5_7[6], stage5_7[7]},
      {stage5_8[12]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage6_11[0],stage6_10[2],stage6_9[2],stage6_8[2],stage6_7[2]}
   );
   gpc1163_5 gpc2057 (
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[1],stage6_10[3]}
   );
   gpc615_5 gpc2058 (
      {stage5_10[3], stage5_10[4], stage5_10[5], stage5_10[6], stage5_10[7]},
      {stage5_11[6]},
      {stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6]},
      {stage6_14[1],stage6_13[1],stage6_12[1],stage6_11[2],stage6_10[4]}
   );
   gpc135_4 gpc2059 (
      {stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_14[0], stage5_14[1], stage5_14[2]},
      {stage5_15[0]},
      {stage6_16[0],stage6_15[0],stage6_14[2],stage6_13[2]}
   );
   gpc2135_5 gpc2060 (
      {stage5_14[3], stage5_14[4], stage5_14[5], stage5_14[6], stage5_14[7]},
      {stage5_15[1], stage5_15[2], stage5_15[3]},
      {stage5_16[0]},
      {stage5_17[0], stage5_17[1]},
      {stage6_18[0],stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[3]}
   );
   gpc606_5 gpc2061 (
      {stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7], stage5_15[8], stage5_15[9]},
      {stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5], stage5_17[6], stage5_17[7]},
      {stage6_19[0],stage6_18[1],stage6_17[1],stage6_16[2],stage6_15[2]}
   );
   gpc7_3 gpc2062 (
      {stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5], stage5_16[6], stage5_16[7]},
      {stage6_18[2],stage6_17[2],stage6_16[3]}
   );
   gpc615_5 gpc2063 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4]},
      {stage5_19[0]},
      {stage5_20[0], stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5]},
      {stage6_22[0],stage6_21[0],stage6_20[0],stage6_19[1],stage6_18[3]}
   );
   gpc2135_5 gpc2064 (
      {stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage5_20[6], stage5_20[7], stage5_20[8]},
      {stage5_21[0]},
      {stage5_22[0], 1'b0},
      {stage6_23[0],stage6_22[1],stage6_21[1],stage6_20[1],stage6_19[2]}
   );
   gpc615_5 gpc2065 (
      {stage5_19[6], stage5_19[7], stage5_19[8], stage5_19[9], stage5_19[10]},
      {stage5_20[9]},
      {stage5_21[1], stage5_21[2], stage5_21[3], 1'b0, 1'b0, 1'b0},
      {stage6_23[1],stage6_22[2],stage6_21[2],stage6_20[2],stage6_19[3]}
   );
   gpc1_1 gpc2066 (
      {stage5_0[5]},
      {stage6_0[1]}
   );
   gpc1_1 gpc2067 (
      {stage5_0[6]},
      {stage6_0[2]}
   );
   gpc1_1 gpc2068 (
      {stage5_0[7]},
      {stage6_0[3]}
   );
   gpc1_1 gpc2069 (
      {stage5_0[8]},
      {stage6_0[4]}
   );
   gpc1_1 gpc2070 (
      {stage5_0[9]},
      {stage6_0[5]}
   );
   gpc1_1 gpc2071 (
      {stage5_1[3]},
      {stage6_1[1]}
   );
   gpc1_1 gpc2072 (
      {stage5_1[4]},
      {stage6_1[2]}
   );
   gpc1_1 gpc2073 (
      {stage5_1[5]},
      {stage6_1[3]}
   );
   gpc1_1 gpc2074 (
      {stage5_2[6]},
      {stage6_2[2]}
   );
   gpc1_1 gpc2075 (
      {stage5_2[7]},
      {stage6_2[3]}
   );
   gpc1_1 gpc2076 (
      {stage5_2[8]},
      {stage6_2[4]}
   );
   gpc1_1 gpc2077 (
      {stage5_3[5]},
      {stage6_3[2]}
   );
   gpc1_1 gpc2078 (
      {stage5_4[1]},
      {stage6_4[2]}
   );
   gpc1_1 gpc2079 (
      {stage5_4[2]},
      {stage6_4[3]}
   );
   gpc1_1 gpc2080 (
      {stage5_4[3]},
      {stage6_4[4]}
   );
   gpc1_1 gpc2081 (
      {stage5_4[4]},
      {stage6_4[5]}
   );
   gpc1_1 gpc2082 (
      {stage5_5[0]},
      {stage6_5[1]}
   );
   gpc1_1 gpc2083 (
      {stage5_5[1]},
      {stage6_5[2]}
   );
   gpc1_1 gpc2084 (
      {stage5_5[2]},
      {stage6_5[3]}
   );
   gpc1_1 gpc2085 (
      {stage5_5[3]},
      {stage6_5[4]}
   );
   gpc1_1 gpc2086 (
      {stage5_6[8]},
      {stage6_6[2]}
   );
   gpc1_1 gpc2087 (
      {stage5_7[8]},
      {stage6_7[3]}
   );
   gpc1_1 gpc2088 (
      {stage5_8[13]},
      {stage6_8[3]}
   );
   gpc1_1 gpc2089 (
      {stage5_9[6]},
      {stage6_9[3]}
   );
   gpc1_1 gpc2090 (
      {stage5_9[7]},
      {stage6_9[4]}
   );
   gpc1_1 gpc2091 (
      {stage5_9[8]},
      {stage6_9[5]}
   );
   gpc1_1 gpc2092 (
      {stage5_13[6]},
      {stage6_13[3]}
   );
   gpc1_1 gpc2093 (
      {stage5_13[7]},
      {stage6_13[4]}
   );
   gpc1_1 gpc2094 (
      {stage5_13[8]},
      {stage6_13[5]}
   );
   gpc1_1 gpc2095 (
      {stage5_13[9]},
      {stage6_13[6]}
   );
   gpc1_1 gpc2096 (
      {stage5_16[8]},
      {stage6_16[4]}
   );
   gpc1_1 gpc2097 (
      {stage5_16[9]},
      {stage6_16[5]}
   );
   gpc1_1 gpc2098 (
      {stage5_18[5]},
      {stage6_18[4]}
   );
   gpc1_1 gpc2099 (
      {stage5_18[6]},
      {stage6_18[5]}
   );
   gpc1_1 gpc2100 (
      {stage5_20[10]},
      {stage6_20[3]}
   );
   gpc1_1 gpc2101 (
      {stage5_20[11]},
      {stage6_20[4]}
   );
   gpc2135_5 gpc2102 (
      {stage6_0[0], stage6_0[1], stage6_0[2], stage6_0[3], stage6_0[4]},
      {stage6_1[0], stage6_1[1], stage6_1[2]},
      {stage6_2[0]},
      {stage6_3[0], stage6_3[1]},
      {stage7_4[0],stage7_3[0],stage7_2[0],stage7_1[0],stage7_0[0]}
   );
   gpc615_5 gpc2103 (
      {stage6_2[1], stage6_2[2], stage6_2[3], stage6_2[4], 1'b0},
      {stage6_3[2]},
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3], stage6_4[4], stage6_4[5]},
      {stage7_6[0],stage7_5[0],stage7_4[1],stage7_3[1],stage7_2[1]}
   );
   gpc135_4 gpc2104 (
      {stage6_5[0], stage6_5[1], stage6_5[2], stage6_5[3], stage6_5[4]},
      {stage6_6[0], stage6_6[1], stage6_6[2]},
      {stage6_7[0]},
      {stage7_8[0],stage7_7[0],stage7_6[1],stage7_5[1]}
   );
   gpc1343_5 gpc2105 (
      {stage6_7[1], stage6_7[2], stage6_7[3]},
      {stage6_8[0], stage6_8[1], stage6_8[2], stage6_8[3]},
      {stage6_9[0], stage6_9[1], stage6_9[2]},
      {stage6_10[0]},
      {stage7_11[0],stage7_10[0],stage7_9[0],stage7_8[1],stage7_7[1]}
   );
   gpc1343_5 gpc2106 (
      {stage6_9[3], stage6_9[4], stage6_9[5]},
      {stage6_10[1], stage6_10[2], stage6_10[3], stage6_10[4]},
      {stage6_11[0], stage6_11[1], stage6_11[2]},
      {stage6_12[0]},
      {stage7_13[0],stage7_12[0],stage7_11[1],stage7_10[1],stage7_9[1]}
   );
   gpc117_4 gpc2107 (
      {stage6_13[0], stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5], stage6_13[6]},
      {stage6_14[0]},
      {stage6_15[0]},
      {stage7_16[0],stage7_15[0],stage7_14[0],stage7_13[1]}
   );
   gpc623_5 gpc2108 (
      {stage6_14[1], stage6_14[2], stage6_14[3]},
      {stage6_15[1], stage6_15[2]},
      {stage6_16[0], stage6_16[1], stage6_16[2], stage6_16[3], stage6_16[4], stage6_16[5]},
      {stage7_18[0],stage7_17[0],stage7_16[1],stage7_15[1],stage7_14[1]}
   );
   gpc1163_5 gpc2109 (
      {stage6_17[0], stage6_17[1], stage6_17[2]},
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage6_19[0]},
      {stage6_20[0]},
      {stage7_21[0],stage7_20[0],stage7_19[0],stage7_18[1],stage7_17[1]}
   );
   gpc1343_5 gpc2110 (
      {stage6_19[1], stage6_19[2], stage6_19[3]},
      {stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4]},
      {stage6_21[0], stage6_21[1], stage6_21[2]},
      {stage6_22[0]},
      {stage7_23[0],stage7_22[0],stage7_21[1],stage7_20[1],stage7_19[1]}
   );
   gpc623_5 gpc2111 (
      {stage6_22[1], stage6_22[2], 1'b0},
      {stage6_23[0], stage6_23[1]},
      {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0},
      {stage7_24[0],stage7_23[1],stage7_22[1]}
   );
   gpc1_1 gpc2112 (
      {stage6_0[5]},
      {stage7_0[1]}
   );
   gpc1_1 gpc2113 (
      {stage6_1[3]},
      {stage7_1[1]}
   );
   gpc1_1 gpc2114 (
      {stage6_12[1]},
      {stage7_12[1]}
   );
endmodule
module rowadder2_1_25(input [24:0] src0, input [24:0] src1, output [25:0] dst0);
    wire [24:0] gene;
    wire [24:0] prop;
    wire [27:0] out;
    wire [27:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_22_gene (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(gene[22])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_22_prop (
        .I0(src0[22]),
        .I1(src1[22]),
        .O(prop[22])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_23_gene (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(gene[23])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_23_prop (
        .I0(src0[23]),
        .I1(src1[23]),
        .O(prop[23])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_24_gene (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(gene[24])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_24_prop (
        .I0(src0[24]),
        .I1(src1[24]),
        .O(prop[24])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_27_24 (
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CI(carryout[23]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[24:24]}),
        .S({3'h0, prop[24:24]})
    );
    assign dst0 = {carryout[24], out[24:0]};
endmodule


module testbench();
    reg [485:0] src0;
    reg [485:0] src1;
    reg [485:0] src2;
    reg [485:0] src3;
    reg [485:0] src4;
    reg [485:0] src5;
    reg [485:0] src6;
    reg [485:0] src7;
    reg [485:0] src8;
    reg [485:0] src9;
    reg [485:0] src10;
    reg [485:0] src11;
    reg [485:0] src12;
    reg [485:0] src13;
    reg [485:0] src14;
    reg [485:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [24:0] srcsum;
    wire [24:0] dstsum;
    wire test;
    compressor2_1_486_16 compressor2_1_486_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h114d09ad0772e27c6e807bdb06fce653b8e5b0f38bbb31880e562ffa71aa43b19d6fa1a93e6a766dd4c4ce79041513a1c1b3bec7782d71c6f890b0e93468b7ae4d44fbaf071dbad2c01c38d435d980498c436f8d79c1b016a2f98fbe2f73001e5f6a2405c31327c19c126bbcb570738bfeed9f8ab45d6ff1e33e36db8a3f9b692a1962c9d6a69fd789c28cadf5be270b8f1067c2c46ee106ec55c356781477d81706f445ea4db40b3cb172bbeb67953c0e48f92f63ab6866b8872c7306e5ccd829e31aefb663543033d4a1a00c4a68023b5da7b4da4cbd2638624ea81e03c2f8d3b6a284af603bdae44e126af221bbc94171fffdac4671fe8f39021cbd9bcbb2b4ef54021cddf0776ea542a2afabb38a4fea17079fcfe0d167e4fafa43f10b13d9e61bfa2c0ed439b82fa384890ea67a5c7db2447275bdfe147edbb3ac7df55361a401584fad0c861c0bafd3402eaa8ca5bc0d2adad9f45383e9a77392df7c8ac80384e5bd79cbb7efb953373cc3d7bacc258de1a03c804d0a5cf3a502c99871929db8d65915958ad1801c26c4d7bc57f025f66835e050607c02dda06f48cf42f07402fe06dc4517880f6f773aca4801efd49d0c824ef2fbcacc1c12ce290b057bcaaad0733646fda430a2743bf3fdbcc5d925346bdfc47c4c32ec64dff1936c88270581fd2f93601b9466b2306dd26cc4a768ca76c0623df58ee2f7d7fd4ee4cf47e32b56aeb659fb1f72326e380821dd116736e586a7d918faf3881c3b71979e8b16baf1f2b21f2d8c14e4d2f9a63737d595f0170b501beee2d5d9730d185f9b8d44c792d8c1e394348313bd893f4f5dab95fccff2af071cd467d48a6c3729753d60ee3cc6a567246d96d61e6f1b7de199c304e86d028a5adf67ede6fd9e75579d51e28507baeadf2c780ad4b709d6cf83cdccbee68846949b6e8c03113a241d11588c98cdeb19d455844e4f7f06a5662e8a69801e443ea40ea8f55d8feabb15c31ab5cbca9d5ceebc55d5f6bf8e70c0c71cf80772766590ea63a7cbe7b4e6a2518cf77e2d23c57a7d03c4d3f1151a99573a82c3f75f5cb0c2ae7b97e18555431f02bd168615496bbfa7d2f3ead1d42704531fead33c0b2e78c5735bb1f0063ee2890e5501fb4144c6069250973d2dd897f5c736d7aca3fa51189522628a28b5cd0e43dab1280cd2f9ed9f858588e0556b8af60a7cb390efb72df675110f27952d9e9d76a58d915ae0b5a6e7641c1a69537c147e1c2e073251b8e9561bb8e032d89881dbbce29b32775af8a54543aece6dceff966ee1170e295ecb61183d4a2643261fb7efd99c639020d6c3478167104f50fde0cd723a4d445cd508ba78040ffd974e0e6460a6f30415cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h5ff7a71bed67b18944ad3e49331f132f4ab901afaed3479332802adcff4b97a38bb08b3030032c26dd0dff4755c1d6fbbb0d9fe6c119acc6b534c020a6b4ba17a46fcfaa4654127141c1bd1b4f352fff412cd8fc17d10d896ef2989be09f9a02618477038e737d8f88e89cbafb134d57e90f6e80af689caf5c7953d2e43e84db0bfcf94654983c2083c83ead51e735bda23c6d80d921fcb8c94bc7af25c7a582ecbce58b4ae923905dfe7654639d568131c68c155c88d794106b92c9d78ee55a7ff4b13d3d71b7dd85d23fd12df29efcd4affb1066102d5617190115e2202dc94ee5e80354bde111e53085f464ae5f0fed5a396f9f7f781529105c97511ee2250ced131b0ac4d8c6f3334214ed0e4972e10d4dba24e500e4fb4b1b68e0adcdcd7f2e91197dcd00d95b2abb814f99020f22720f6b7a19c3af7e7cbfac46d237cc92b40043428a5db619f8e90e49670f6604f92eff5ee0facdcd427f36940f61fbaa649862d23e6b4125fcc6a17ab59347dc771b6044c654e33e1cd3e393a6740f6db5c8d970c6db791375185d1160e67aef4dae66d2647aea1bb45231712be56de23a36c45e445e09456436cb11a50da786f080003e1d13584f6c4586594ae13a1fd21b076cb9747be06e17dff8ed0b4eafdbbe396318fdd9f31fe996968819b9fd7a3c8417401311b6f1cee679a81483877956731c05818e48a947cebe9a707fc16416d46db8a0cf0a78e4bab736c67baedcd416adaacb383b7501535eb41e766dd39ba058c73772f5272cd22743967608fbe523d4cc78854adafb3b5d363d3ba8fdafcd52738fc09c14168d75bad4b022c4116e08b3591b452ab98012d2149d3516bb1d66743bf06e9bac4b9b4fad39c74e1f1810301afa04d60be187fac33bdc4b312d190312cd240616488aa3e1405739013343f39262fb5ec6a6f3745cd7e09ccabc16a372629bc226bef6743444b10f35af22cbfbb62586303b40843a0825a687008ef26a0fe98726482a7f0c30618048c899cfd55c8361a6c71349e2cb8dcf5ae996ab6bb50188bad3534b2040d68606587ecfd8de98e2bd93cbcce16e7a79ca68ed46b7562f78bf8f9e0c37b92350336745309c689a2718c5294e411da1d8dd1e0a264f8c7442f0d16e33e348b72452faba2016fb976e10b8e4d4f6efd266f6e09fc26e3fa874402fc60509f8990339f121b66ef319317cf5c04fd4f6d149f0ab5ce817da389f9518b34fae1155b06515e7681e64eb3d092a7374a52aee184450e3271e00c06f175efc5c0430badd52cb24de9a976be2f58ea9210f28b57cb27203d8536f2a2880d5453a7af51fb7831c9b1f42019f89d7a5321fcea0aa6f2522b14c76923084ae4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3b00cb27b247478ee6376761c99b667c1e1c894ddea45b3ad167b6faff25742e7a04ccc0a3c78d541dd5375d7522c492815a76dc8bcd8f18a083aab49287a394c1e5c1450f274f67dd6f7e927f8be4c638740154e238decdfa62b3b6bc9cd5317fb6610d4d4ea8184ac5698dfebc13df6a058821da5064f990c232aeede87d3ece52e57dd5ee2e0ac9bcb941fc79771c2309227996a49b905138958c5605de924da76277312bd8c7f2a398c650c6ca720647643c797acf47d39adbcad08013c368d79ab614d1ae44bcf7a3faee548540693ace23605b07fed866fac220f6c6bb4fff376137ffcef61b403a6781cfc154e3ffe91085e5dd21a3371197336e59507dce984dea1bea94e04ded10cf7daa2d910d4bfd8ff5b1607b2bebb0c1b91b4db61a5dc7eeb574063e0536d474aaed0fdb4f3db417cca9f8755d07e20b21d356f811f6270d879ab018ec8dc8fa573c23477e44f209f657535d653bc7e2e2974bc6cd1b13977516a824562d5bb627ba7c713bc4c86effe3f672650ca630deb9d783cbe3b98189b959b47671810d1192b94dfa8d0a4801327ab9b479e31746a95daf5e859401d2705935df00f073ed32b634b50a42d9f56c5bfa8e235b29cdae06661071db8ba36ebf4a56dff75a918de6357f563a8323f07df67ccad78534374da5131aecee6760ae8b48bd21c618ca56ababb2812d1481c39ecece6266f074fbb3dd164091e7e94222317f04757743587577912684d53eac8d21bd38408db63711a59981e08c42b75091fe017b3832242a90bedc3f5008a21b22b18600a86ebfef67d7bb4a2a6c11955192f28e904c3b21badf33cccd2f791027035e9e20a7d1bed7389e14b256e003201c49e4806bcb8c0c9d3342f278f275c703e49c106035ac51a0624c30c4ace4001a98e581cc40aa852d3749491f42e76794afb139d3c2b6180e67dee8442a49ca0711b021d52036f47bf4deff0a47d8c027c911a5727fbe74993c54abbbb3bff6555aa12303b58ca01b0036e9f381c350b923beb1a67ab0e9bd3574da28f2613b521990933e63837c8b70e5cc2cc571c70b0616a5a9184a62296ff16b9862f307ecc327c65eb1937d95a9f8c54c6490c9d7e2c8c992f87de3b2b0bfd59660e1d1a0ff03a90703284f5d2d66400d43ac0f782cc718fffb351577bef54739153b9f41fcab8aea172f481efe25ed9ff300aaad6a5d2caac20aa7d5117e742e9eef2318e7503b129d10daa8bd1fe6029b0074ed7790a5d96a95bf13ccf4fd1a2429fc415551ab54e9ce3badfb3b8cb06e47e489ee92f1d96c3374f68033f1104d60d36655aec7240258ed0de788438a96ff874bb6d3407335b7c0d934d31d760866c0fa60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h917006ecb1ffa859c7deabd893780376b31f0052b6b1c8f3baa10f849aa7abbb55c9aca1049c93471b947ff396668d003fde053bbde333597bcf7367a604b6af8779b11275e290a4c3f3eba73a1090102489cfe976d2d4874b817793c0664ffa4aae92ebe47cf5f6105b28b03f3ea5918d4b58ff501a7ffb1c2fed0916edf6c82e24bd4b3a431e8992e02b9a95a722d27674a3004d39525ab6b9be5ae14fe4d75a667b28bbef455b036bf62a1b933d314e92be0ac6d27c50e13501133ce967ba69b229f4b9f7f88e3ac99da7b4f61723e3a791d445ce8875bda846a4d7484eae31110f9b3167ea228449fa0942083d86d8bdcc7a3007480266d4dd9f1e32104c92dd37bc6ddc83e79b56c7510dddef57b41f9a0c8e47ab9b56892fe76b656eb102bdc357e5fb79d136a3bfc9bb7e62ccb5784b3d2651a00ff7c8ae5a9d52d7cdac093ae8213fd3aad0b6c90ea2d2e0ce687ad56d0bd1096964c2b9fe48f62d39e123abeafedc8a400f550f6f29a0caa74ebed69bc29913b3f4f62f261ec79cc5ac99352b8934335eeb568e60d77558794013812079a5c641191809473970d4d06f1a5649cb3f3f7122269fd17f13e364024ee8402a68524a4a86cc1c0b35dbc0055cc7a7ee763f72a1b42196080da391f05096b5fa757b1251ad7cf31953f188d58aaccf9abe8e7cfaff9543ab579559a90b7dc9577e27a60192dd697dd8cdf1037a846d9aef787fa52ed1085df7c9748926a33a064f1ad97787146051afd418d21fdffdf7ede72c02714328e2fce47e7e4ef837f560e378492235e38f96ef0d1fefcb1def83edb174f83003371c12b23c4aa431dcaa837dcf81b693e893487a10385dac9ec1fcd2874ab4b4a75a889365162109e9e6b20cd3ddd9db60318de8fae89ec74e783c5096caa7b557a862822c0285deeca98932a7669d4841232938615f13e44e98206c82de19850e47344f7a83f561f7a399bdcb4a095d9d547d2cd2b387e65ff0284501accbdf59ae808afc59b576d1d64874535582f586997612858c2aba1d0a5a89d80bc227610e54027848ade1c39e3372f3ee6c3b7a3bff709f0fb85e766636cd9f96595b73ce7be636f0ced413c30abfd583aa0be5142ef8aa52ad7343ddd82fb5a73c9c00576e3dd2f5edb9e671fbe13cd881dfc9f6bd7eec819db195908b77a37a1318930c7909387a5a86e0df938f60687c10265fe220dc17ffba6380b4c046645c9d1134cefd231c9c81aa96ef25c8c8ef279155c515a2a582e51c4632bacf2e859aadfadf78c42e69cc56bf83f5d16e0ecd98e015decf4b58ec0687cc77f146d18306271086b97be0d59f0925f8edd0527e1192db9b421405c0b71ed99e5d5b678a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h90d904de3f5ba127cf4fdf251df5447279542738990551fb668c643271ff48129e672db77bd0c77f82c0c7f20724dba8f0c94c0defc5129e4af3c34b2efcfbd3f84b19d0ee34def69964bc51bf710fbab134f9896023526a3012a5b9d09b18a5de63ad551e1c171a1576b480fdfa21a5a0aa3d7adf881b13a7acb1856322975bd88a466e335889272694c734b1bbb56ad082d3caefbb3c5ebac5c55cd697da40e34333c78b34143b5f97eeaa3fc9f7febb4db9e2aad5a3b0c7b191be886c8c059944b892f4da0685e39bd6bc6d1019d4c09f2dde6f040c7fb9d8b352c39439a98ce290db7af1b1e17a688c6cfcd3a5db13c577712c61e92a080e93340392f3b358218da9cbb28aab2e9e470af9e6fbbd5c8a9d6564dd83121830b670ee839525e437823427115ffd046e5f86f1ab650e2349c15dce4079d02672651fdaa271ffbd72470980e75aff7ee734c82d718d4285ce7ace4a4bd743187e0e6377e571743efefcf5f4d05365005d668ae3ad8c8c73c180a72b2872fe567e547d7a6b5209abe1579d241e480214a7573e3a4603130be9e893921f7925157cc5e21531167bef6e862ea6b1635cf216f9339e945ddcf1a421d70198c515c59166e7895e2d1b9dcb2216b1d9e8b0d35090879cb1441c55d0e4a814d73c3ad882af7e54ec1a8bc7b209e6d06d06d1b28f622e7e128e6a3345e5eefa25b3de1a26b5d159ed121ef6a4bfa64764235acd1d110737e4000a9db3e115bb88851fb438d194c18d5c79e277cc6ef27c592c07b5674d05b06227a9b481e32503fc59a2f1395a79c2c88be79ca55922031eccda9eeecd0986c536c731af90dda8cf4ad7bfcc634d732d0bcd31453c5f53e59964963606f0c964f788da82e700c836a55ee1da21b434ce607367a861217a3ee0980b4b0b731ed2aa6157c9e57b7a0927b043d3a63c12c192f62ae33a0dfee85ecc7a256633c8f03c24f592027f569ad78f1cb7949b3603595ceed6083636787f5e7e2e7f745bf538b4a926ff4515133e226445d62a9647c589612d26caabf4ba8a11db9a2fc598af9760d565d0195ad837c4fd3166c9b229f7c8fd7c64bbd6edcaa477e23b76ee4b61b967f7bd46aa4f099dfdcdcb9fddeef5f9fd3bd47c045810f2133fff6067dfe0682474e197fe27a10078915996195ee1f1ef8e7929efd48c1ab76485b7deefc7c3c0eae5ef7a0993ff3fd6fcbd419cd315f69027dfc569a304e7b2c2d37aea89dbdd2880765557fa2c1b25ad15f50d26b3086b73c969012f5b88db20d678a64a0ae5c0da531701e23feb9454e1f6d7a23acddd83ccfdab9be6f937b14533d5ce2daaa0fe3dd4cb259aaf4057ffde5f406ce20e02ee67d12682290f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h912162536ab501ff736e78f1a23bcb1e51e986ce70917bd32d0f3dce421ff01ce209e9134d6b2aa15fb91c3b02dc6f77559466c6053aa1e98b59e9bb017a046beaa7f065aa08e72c4620b92b12b7be65916caa0a5e7b2846e403a6d16b116ee93d1d32c27f97dfeff43d3e94437c805004d41035c5c2f6d94261a95a1d192f16f01d0cf5ae15664fc64539685afc9581da02d67618aaf48ac8a5e43514021ee4d4c412bebf5e7ad186e07fbb29340ed16e01947444d7cac5fb03cefbade956fb5741f4ac27266751e1f92996a1c16fd6e6625823298271bcc37435c7d8c465f3a2a38fa124b87c5a754a8e57da6f777985254d46d1fdea71202ba1137bebbf64245d73ed9feea2827b76ce61d7bf27c13cc717537a2fb2872733951c912016a61af5636e52d123efe41070a672bf9350160e354cd43209626d134d0977be9a673cb015c6379ab864c535d65a40698f44758d2d12df234e1a52dc0fd76581b9e5e9643dad68b815131827395d3d8cd16a94338091383937d9278a73746dfcc20de3ccbbdc1a56060ee69d836900fabceb2049362e6e7169881a79c5d7422966c0f3c1ad6e61a7597999c1835bb74682e1a1810b470eed69d391e900e9aab049111ad810521d65bc63ad7db1270055320f711e7701b149b061beac2b67a8587c716b1d5888f5279ef02cb3b43430d2786c98355a80a96f3f222c551ad7df2b4571961e5d0e532520b79c482e8df8bb3095560a66717a85699622ad379c166630767d92e0c73ca07df583da95531da4a96f447b34a90877139636b3612bb73ce3d6013e6fe101de518e06bbec32aec2056a335775930155b66407a6397bc648a0b3a91ee09bd637c0325d513ece9b611b1c0f2b71553b1b3a1e2466a8e2881540040cac5a35313675ea14a4b1282ae2746983f92caba5b0e5dd9449b95268888bbdf30f31fccd3f46a3595ae2e86eadec39852c6abc0a63ab9a35c93ab7b7b5ef3faf1394979af795b7ec2706951b11b738a7f60bfb5a79e3acca26edd5230af3eca277c876bb0b5cf8a78f771bab758ea5b5067529e85df1520d07a6929de379f552a344a0552f45303ed6d4cc315e5d550497375eace00e4bad11e7c9042055fec7d61db23188940a53cef9fd50646447fdf6c2607887fc054c7bed145186b6e2c7100a738a1f50144b6cab6c2ead695d52ecad518f2e1edad74391f77dec532b91f787cef0e8bfcf6b3b169e1e24bcf08fb00d0abdfda8b0f3564f9fd9fcce47e47305c7b686a494cb2340b43dea40467b834d273fd6c182769735ac6c2861572acd9cd51b34d577b74c24fcd40c52a1878063be072cf3f75d0642149cb807ec0589d4f631185d05d66cfaa4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd9d241a089ae88a23a74dab709e06b8f6638e2fbdbc2a6e7ae718b40e2550662488ee6dd8af66bbf7de2be3f33bb52af2a2ee1ca5b93111c4e70999f144973354e1da6972b31a791b2c14a2ac5f427110bf0533449a22aa40f68df1a11705c868a9bf735ec36c8d39c63bef56497e104c3a5db02f8aa8213d926dce5549d6e907ac89a8464d73faa2b5d856507f16f8f2b3747274e8781698e170d1d7ee5c336a34a03f9cc52a2fe9122d7685fda5240ca7ed65574ae838e11c00f74102dfdaf914d2ef082617d59a2a15127319d93593372ea3680d613ec6a4f835acf9ec86ab314a10cfa4932dc79d4363f4db4bad70735960030ead3ff8ef080c3c21e347edef91b561aeacc7ea063273b5eecc9d17f3f52071f8a8091e7c709d3266631bcd9432c0d919ef34e45e842e28580a30ef5810a88e04ab5ce0e7a347e3246c7dd0d551ae7c35dc5a1b841de4a0b14108cda8b328aa3a9b8d6a8f1d03ae784f30c1635feea267b95d9dab9bb99747728a709b6bb924b8a8808a3ec5112a559faea11d7650b15a28e2004af585a40203404b81e116d7daa8c7d9ad7d0d9f09493049254b0d579e42dcba504b18160241c69928251248c06bb555c0a4235fa76835b89b42225919460fbf2b258ecc46b35531542b377a0ba0e4307b8d5b04d9ffb6ffdc3dca7532d1d5f8ea75a2e9a348d5c09c1d70e3e85d3b02059b2176fd98adbf8c88f4c65b1560fa3479b0eaed73e4fa4bfe3a754605f9b4967c24bbf2f8639962ce9e992fbb506925d962ca9653773afb6bc86fdc674ada154feded61a3fe21248a932e77b3eb46dcc729c33ac593cc6c6c3505849f5895b49cff8b8ca62d09ea137f8efe05694541cd830bcbbc08407b6232b99f35b981d3a6e55e03c4bbbecfa0d5ff663e759d965fe72f646041115ab30c5aa0cd8b7cf21b1189c117907d14681f0353297cf6f87626085227e7fc1ba6e68d9832284edf27bb39d992fd5bce1865fffd76860af735720dbdfd69e5978389f5b47f8e5a2a6b35a132d977988776ade5d7e399e1e537da3dd741f93c816d3d840017fe593f4eb7a2e2e40d9d315318b23073b57f556189c6a276598f337da43d2e2e61fbadef7fafdb73664af81030af60ea8fc3f742a7b4956f718a7fbf042f43e7ceb75b0a24289ab6a77f8fe70a4f4c777afd814ee3ca2defb88d9dcf72b9d5abea6d0367de7095560108182637e938fff9f9ba459e798b9eff9a3881e1c7d10f3d6ed8a25a253d5ff23ddf3ceadabee0fd6d2c008ec4c97f28f60225099a519d1429c1b882ade164f3aed8da126f235811d0e605fa5463ea63d27821eb57b261e7b1869cb95452e0caee4ebd3e195ee58204b6c5c35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h463cd6ea3c4f5ed6b366977ffc41e379f5e83d380a19d0b09ab889f4accf4a498905a44b18e2815a9ad8936d95d707c81380588b2640204c0e210e39e6841d9a49219df312f040c01633422139abfd7150c0df8cb178a28bb7d29343151a76b6169c3d3a58e35e337de781ce0b994a6f2c2ba67af43ba1444702b06223c0fc647165734f37ec269e37b95aed538d684c4fd1d41ee4a8973241653a39b9a477c2b02f2aa5992f102f34a87279d826ce5602f013d548f684f1d6be3adac01b3ed4cdd8290912c260685aa93caede97e4b51a10ed15fae153f446edde2e5ac1d434bcd62eb7769e57c2953ddc825958b40bf73d708ed56d82441263564c909247ede559c53cbc2a89a9d756972dd759e9833a6105ad0b7e43c09b2dfca9697e2021f379f9bd9730c54ff6bf0849b0b57978467acb9dd3d32d4931ec3061d7454abdc763317b6c00087c7a66eabc57c22dc57dfcb0db63cd8cf17c629f831512740097688d886f70f59b7901ee24f188656634a3df205f3f0676a82fae1ff3256ef0fcc154f1d9bd99029ec09eb74069710379becc5a415983c5237ae6c7d81e4597e54c68ead62e5b687a7a29822f9bfb4e1a3392055aab9a32843e8df3383782fc0577c66b32e0025dbc0835aa7b9097aa984c961964a6f74ec318697a9ea9e13ad22e45b41986f9eb19fc35a78b300bff6060b692021b97170da7109d0b7e61832fae33e23cceba1a4f5ecfff8979ff9f04ce174154108d4d38294e17c468210ce9b0be9d6789f01daee1ba8a29f88ef769c236f8691c796a7e58dcfd30fd8d9d842946ea0c1213f42ebf5977bc5057b42e77b452355d0da45193e1f71f22432e8783a4b1baa3a5df4627489449a406b20a3a34c533c077f7aa5d09bf1221d643d8c4525274c959fa21201cd5053c94aca5b0f11ae85e4ee28008be8c0a8c42903191701a00de08fb8f18bbca29e3c2fec803706234be799614d2eb75f627078d0eed176727465208c550b314768abc6ff8baa8b10e1fe98d08848832dda41a8a409bf03e21f4bdca26a741d37412045abe4b22e129d03a4836b29365717315cd9b845bd4dbbaaf58e91e1067112dfbcdbdb1d5dbbf67bb3f222dfcb070b6314fcf2643c7f998dd6d92bbf1452fad7c4a9aea82d655032524ae93652ff17ef78f60123aeeeb82da45a7fb8834f43581a8ae44d37ac364c93e0d18e07a9a1fb7000f6747d8bd1ed7ec90a2703f27e3486ec89e36743ebf23b0527e374f63df5210f6c4790465a3194e671f45746b7d75c395bcdf529f8f389987b4fd501010c2530bad36e1216b22a7d4aaea9cd11c7b3686434d6bae3a9029164a4a18e52b1a0aea24a72ca5ce44862d528b7a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he56b9b56ed452d5aa0b84e61870cb20a3c7818b6c102a67efdb1afb50c0ba9db1a18c6c631c1a184187637de15264f1a81b2f53b6475804aa2ef7e29d5bdfaecdb4fa7241593e7f283613b18a695cd8e8d709a2b25e24526ccc8f3cae574cb06ce41a95c7d3681d58bc94fa3137177c522400af197205278293970a4cb868049982682c6ae6f6aa98a92b59a47d61a24b291e8cb93a58e2e7687e184b496f61eca0f66111272f8196f56b6b6cc17353c52f075d4ae533832254387bd7004c74fdd7324c8f460f2bd4148b1fd96123eb0ac6fb02ac2ed1a459a8534c9c3629e4e454c185e14536ff4e319a240746750b47d3df7ff4030b659e845280094f785f45d61df82206c14d63e0f20f4e20c0316ee8a64cc758de749986fcf127fe8f276eaaee4d66aafd25cf2a5696476cb891c0f44d2daaa85a0ba378d1a15cc770657e436fa01faa4cfcbeec2b6a2c12e6b1f8daa80c545ad573e58e25340b8db552195abf9d413e700ffaba3bc9a11369be5190c499dcd31ade0f05e8e1a5cd8655329bf1f544e4542eb520067145d8e95863c440d5302ca81b3775d7f8562159181888dad403663ea82bcebb7094a6fdc209f946d6bacefb7d936f58c694ff2203442aa2ba8faf2558720a1ca8eceed6fd2b72cce6927a3496b20f8ffac297ac5241841eae0c2f164e5bccc6b6572a79b3d2bf6688616110f85ed0c1435c23a0bbfbc53649afbafa139448a32a11c29968bd5d9719c7bdd00f48ce71478a1aae46070480ed2ea3133cf6d65968f7ae47137f396308431fe38274002c457c0c85dd6f35f013b95d7c309bb82b7e493eb4b9e65582b10d7268ba7dfe99fc6c808438fd96869171a4fc08775ca67d6130ad172cfe522a22506a85857168848ffecd4def7cbeb064a583e83564a9d873612c3f8c89ba349b460513a923ab3da3c33fe3a00ae7c903a1011735b45a304702a6968f60f3764dbe37b8e5fa9edc6772104f87225b9f74cf9a1b92f67a521b19c7d22740368f82f11be9528a6a84191d8f734872d394f44f65bfe62f3f6d76a95e1599d7bdb7e564862e00efa0575b719fa63c322e6e1e220a64073b7822a1a537857f0c43483c7cb231efa46fe31c6a710e1cd6be8e4cd1807281eebc7f8c4631dd697b3b86c68e22f3d713cec9e8c6b6d2b186a1c8d5adef9fe7d057ff55a530bcbc355f08355246097ace9ca852abd82f48bac15b95259ea130da36c00b2e46b40cad2bf3fd23880c6a533cbae435a7c7d8cd35a80f64a6dab80d13fae7b5ac0b3f3dfa11f58e79fb09ecd3f9e1e27ccff9f946283da6510eef6720f7f632b64d46336f88dfb08eae7f72dcea5198f7cd59e489b08631199351ee1221f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hbc77f24553eacb52df151b4c11ab6e0de2b2c66ad16c5c2388cee5de3b51a6e65f5042d5b12a188a2981744429e3c22ec9200cbdc044928b4bebdca7368d88732d3582ee1b22aa2bf7d5c318cefc90e67dddddd3d669b9afe870cb88f46e6c0eafc0ffb687127d708701306f2c012b461256641ea94bf81eb1fe5db47680c04b202e8d37bba2c109650f27925ca5db036f2b882c97b5bd7f73cd6700c9cdb0ca24a68d07167b3743f0a0def43407002b1fbd380d02c0aaf5551677f8a1ef38a6a8d6a1b48926816754feaaf86bf1262f2c57631ce5346260d51af88841cbe2412079b444eee93ede1dc542e51e38dcb4441dd63f5e0cd233c5fc112aa67f71347a4fb972453acd37d020258b2332f8db4a1ecce257b0d5e960ec739b840887f972b4635ff5b3261a9b0662d25f0a915207eb61199914a28c3a2f5638aa7436513db17b33b7a85bcac9a04c8d0e1625153684e5ceccb321e6b200199160989230f88ac063f45df60f9cfb87206507b55c4fe04108eef323458d333af974f9e2f0e7d2830952b62106cdcea06fa6427eb29496de2515ca20f317d976d7bc57cd4c74c9eb50b468c89b77de3fb102de54901b286a2f8c269f9e24f18eb28b3efde04cb5f9f0e58b194b7fc60b9740e92877e6f444311aededa8a45bc95b7df8a8c3beb7d7969267f2815dc385e9b5711a03372a30bcd8199a103451a50d11a9817d4e59717f4a1a44286280580fc1b1d10209c5e0a4f8d0a126bc4987770c0ed3c867e7985e6853bd47a267064a335b33e1bcd2fb440d27a1d604ccae176924159cadf1eb6a00119893ae22f2ed4ad697c09cf527cefad88fc4e9b2c382d86fd79049b28aa19625c6a1275fa14d07cf89a45048a4eb23651139226bff1399249735d29594b93cb6becc67034253646e3e48a1b87b0a791e72d0b441f3a8bff0c549f7215ffc63766485c9d4b716ad38216643f2fd0c2690366e7d13eeb728dd856e52a158fa535d5e96097b4864067ca58253e4ddd04461066d9ca2052264b22633d7571c0043663d6b7856ae368bf7f1480b896fe9de35774a2b6f86061ed497ae963d95e6582ac66aa7ebaa078d39cf9520a7fc83dbf75809bc19d2c67788289b19d881c6bf8fe09eb70058bd4f16883473e4e4078b3a2d4decd617400b075c979c51e44d779495eed4abd47ebde7487fdf2ea7785947e6855a09d8ab2331852e9a462c0cf5e762fda8874e681eea1142409742d393bd3c1486fe1f22a185d9ad5e9c748846c6bc07e1812190153e22695e5b53ad2e10080eb1793eca256727d54cab062334e87fb96a66464626f4f327bda620336fcee94c0d36568d5ce01b29e6767552d02cd3ba926fb434;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h77d31b44233db693e2507704471e70fe9c973d5077ba4dbe861550b9ddaa14620bacd7c766090cf68415567d5979d0596ced8ad7fbb876e6a747e2ef494056d4ee444a592e24073fb5703a28caf3217a685467dc15e768a9898a711c496eafcefb2b74ed5f70fcd66656de7b2918540acd1dbeb7cadaa348085098b473e966c6024698a40a0bfa9c269679980bd0394456bbeaca778c047225bf1c7b47366aef28d7516c85df4a2d61b9c150f395780246b10e0efd9942fec896ed26b23924ed41069f068b8a8319f8d057bc542d984eb68f8e5762c1ed5f38e22816a2734db8b038a9976a7010f1f415c088c2f425587d3706581246379fda8662052ae29658da70e0cbc6aedfe3df9f222cd21e3dcd9908e0798f48a6082368c7b646db91d7854d8be8b2b48e8de25466cfaaa1b815e7be5b430f243646e991267e19e359562c3fc233e28498f211ef1c595d181cfd2a15173724612d7003e2e99ccf14feabb0ab8ba9cf3b0d23e063664e3f71dab802cf3ac3651de7ea36db295631199fc048f1aed11cb473ce71e0b56e8697ff7c7fe51d435e40fe2268eed810900e41f2c32946e30b10c07fcfeac97bb080aa12cee22f1208d4790ac578c044d595f3dc1b5db0bc11de18bc371ffaa09f6e904013dc428adfb850e3392c72bb9d1b00becd20fafcd2fa303874e62044b4f3525bc6e138a9cffa42a0fa24b527aa3e0e5e01bb9d9658aac46c99a6dbe23bff0ad689c1988224397e2132c95546936387d1603044a5a7b861cc958d6c9ecbe21d385074118eeed851dcbda9902c82ad564c68007d76275c4ba06675fe743e7a3eea092773402dc5ed94a5272bd36a4a87e45f9dc5f01612fcac5b8faa4281d3d6b5d7254ecab455213780054e1fdf79495883eca8bc74da65de536a893b19d240ab8c9fecb71cb8c6c0d6bc6c7d42513c7d6b744fcda8e56562ab2431a637833a413233473e823bd6eb116eea69423bab43106a1483bd6bb0582cd9f909689c1a9897e217c0614e966edff2338a49f316519e68debd50946b3d07eeb1c75b76b16666c045c88ec2cad1d787caccfb1f0def602aefbdf5cb4434cc42e407242041b20f4daf55f66280c11aeb061ec947c9e8cc9da6d4405f82b62676c27e6193877e136c9c77ea53da85a67515343965fa2e0330a7438ac7fe42f824ca4ba2afd86e5071a3fd5924eef97e92b506b3b959c7e03cdce153cbf091dfc6e070071b77888bc6f396d73fdfed118326d6954e4650bf88510dc756353d3e424a32fd0c41564d90f162a08dc0dad0cbd6a2027a3df9ddf8c45fde439223a7ef1461ff866d2e4c1336b2efc5504bf7c3ee057433b31a02390176d4d82f781d5a46a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hc167243160aaed0670179653f16ee1598686bca9e24c26bd67fc625c0c292e381ab36fa3dfbdd0ecf24c0dbef68f68c57b32a41bfcbd8fbd159ac223f968bf8ed14801e3997befc99f91e6b15bec74dd96c58ea91b771b138b47e40a3256c6cc87b1aca532c1a09cf390be57eb418b92f0c03625ddeebd98ec54de0bba10a9b59351798e5fade2253ceaffcdcdd93a616ae2a4b48161251a4c48b0ed7b35988a44c1043a4fc2a23d627f56f9d79fca63ca847a11814040773559e6846b8bc21ac7e7c2da3d9bd78a2c692a423699925df6c6398058c80cc74185992aba32d1d134419b24fe9d9409d32d749a7ab071d663b77282fed97ec70620a3732e48c9b776a7d4f2293e7c7f7c8ec582f1c07ef07a521c1453ec151f1cee786deb09b676ac9e42ee8e755a3ce6f8123242b49e645582796042a97a8d0cbfd8d5421d86f9d697112c82becdfd5e477fc4d471d2f2cd1953adee3f1dccb96008abeb7552eb16b87c562ab2480920a02513a5d618b3b96d2680f32bfd605156669de9a3bfc89344c4c746b30eb3d2895e7edfd1486da0f7cd5794194607e1a08281b496b42b61c84b5c0816b423232c8c66d68a1b00d8f35c59735dcf17c44338b4326118cd6c5432bf923f1f3b6c583779304b68eec4dc9dd591bea4883f68ac4287b032ca615dc9ccffa9d7598c635f636405c91c71a7ba5d45cd368fa4f85c5c59fadbeff3ee02f93f0cf4940eb895c790623eac424c5693e3d2855ba902ee75119bb8e07a7e8d421e9ad98b825453df69b9c488c904ee811eaa5327946ff4be0efa1aa911cf50f3ee4affac2b50eefc8123d932216fcce394ac3db9ae69ec95c6d16699608c1b35a7c942116988056d9659a535f899b5ad0331eeae8a8570d935c2bad9f5e9ffbe11bb86758415259be17b169af919f6e309cf6ba2f88e64653bb16f53eca20639b82045932a91190989dd313b6767dd91b008010d0e992470c0442109f6f87b2de9e185c916887b6b9137aa8020d416810d0df510b0deecd4519621c8060bb2f82de9eeca9b95e92f2e81e2fabe9062bf4ab86264e0e49ba4339d9b9547646fc251b1e0f9c8e10ef6527fdb2e018bcf7caa07e0ac5d26c477ba0d784e92825f5ff84ba7830eae7b941399c01a3b80e56f2e017980ed3d4da1ee1c633d2b57439dc7a2cfd2e1515c02eb6294d765ca5a2930447d2245797f4bab9855ea311a39813e7aa8fb242e65b58fb002f8dc36eb1689aee1c476a6aca27b7efcebdd266fe3f0d07014e7c340102af07c4ed62197273f1767562a110011b2cd71f9ca4c52e5f519257564e382316041f73d4772d5a96893f34064b46e9dab20565c7825e5755aa59550966faf6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h21c51572448aa1a658ab835370a5ac3cf78a633c4e13cf4088400ad250c907568df6c1ef9903be1844c851f13949c2d39f177207792bdceef3aba23f91b0ec7f3786cd155132032d9e955c1c488d67e684ea777dc712b20e82fc825abae08b6e9e47601052d4e66d725289a28d771f29528446c18b3011eec8254f97f32cd1b677d723ee236822dd20d6882569080da170ae574616c50348c92fc561e37019021edf90f2495bfe6001b385462502b8f6dce612635c4acccc49348255b775fe4d3eb5f6281921315ca92b4ff2f759ce2d1eef251761f3d875e3981aaa49cd133e4979952a206c94efde7a42e5945916500a150c39c5af0e04ce584593ea046aa484843f7b56420b1352e88d2593b306ccc5f32d5ec56e6bdc2fb09eed45f8b4f7d03fed9b161d1009f08fec13f89611abbf04b7eb98e59ae34326d73d2cb95fc421d33b65a92608644c0e8aafb6526df62a73832388d43a3d1386fabe81246dc87306eb9851fa97a1438b9574023220a0a857ca3c97d5b06e9ea38ae6810f1b6e91b346528acb4601ef19e83aa1ac76d728182a676144ccd968ece7882ebade77a9b9b1645024a390a7c7c62bcc902c01bdd6cb594887496f494731a889836bfb809f240117551c936337e316cb52ba77dcb8529f07d7234b30c4cc72f2da35153301f7f04a203b8a762919d1a7abb491e0f70c73667ca55a22e35d6a98723540a61d732d633119e0081b1c72c49edcc131e6bf69fabc583345a15dc3e1ae06b345951bd36ba389362c816ec28dff663a9ad277b0a96f7872b4802838f1affd3ebc4762069d077b40c6e3bb61e1fa8d9ec9be07530c7af3d5ee4cae788d4b09353da577b963bbe47a063af3dd027fa57e70320e5bcf7b85c186aaa687d280dac53b8b0ab99e628bea471ce7b3bd3c715c18b2e7ecc0db1b9db1bbeb2bf2f5ecff0b02c6532feb8569fe31b60c583647de7ace13e5f0972db977094f1aa40703327716ffee90883bd2bdb183806bca2df13e1799cd20b2c99cce085bd4460ae17e3f8726789c88fdb5fc9805b12d217573a78232892d5d23d5cc0a59a870d3fc6658fc30f281ce22aaf97436549b64d5ac62a6b8f967268489ab483300958fb777f6c9c89ca5f5cff1b3602778a72ad784a0ee19def2b5d8690d85873a0ea8775503d40ff9620ee7f69369c23ed632daa2ceb2594faf6b77f45bc98cf5d7204c89ac68f65a663deba7e4150c13a2296c697034c8d7d31ce9a20314d52ee9647737504d69c550dce59817aee4a8a5fcda3337219a2c68294b0c4b30a670472628440f8930f8700f412278d48c6942389720ca4283dbd0ec2f709a3e137d86f25b6e110b178f10981bf4dd307eeb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hfc1df316747da0f2b36257aab2a0c6e499db4239c227392a645eed4a13b20c1e9e779523c350c6b2245e724c8cd914fd08a4b40cf0b3720adfe6111da7d36342eaa0a3cda72a79b2a4a9ba5b65519b9a584690cf37134fa26d2d50260404fc765dc60d60444040dabfd64deb83ef06ac55ca76b3abf272501ef0bafb6b8ad04ef498088624c075e2f0d8e975d42dbdd84a29216d336a265e9bd29b5ba338ec53477c4ed4916afaa4f9ef2efa88fdb7c2ee3cdbde9f3aa3395bcb9879c8c78bcb16e1c2ea685662173687f4b1d5360648a790d1704a122f23d2c0550a9cc5fb5a1962a88ff6f51ff52607adc1bfddb4fddfcd565338fc83ddb4dc37a33b29e7707f15ec1420f015b99ca7fbc6ca3ca04282ff0a9c2502ad90ad2a40d296d1fd59ba27fe90f312ee32b62ad106c6d0078ff458386b50791e03d2854b3103e2b8e8ab838a0bf34c8fd462a390fafecbde8f4067ab18146fabdc172b85c1a7749e222aab3c8524e6b5e935ba1bb8739c9dffac7a82d90f529412a1bf4010be8cb16c748c38ec1a05624c1ea44a3b1eedac1159b0d750648cb6d6e66b159d188c57d2028a7e468502c56c653b08e70c6b0675c7c12f207530c49732fb541992a1647c6643227fc4a3349e28b370b3a22710df22ef6d202cc157e2b3c3895b8260c795f43c27917651d6ddfee81082c4e44c76269dce54edc711f1888d48bc9d13bd3ad8bf626a38865cb4a72163b7385a95ceb37551c194f2d6ee7520163c4f5ad0a3a59546a24333199a4dc93348197eb8fda570d0f412c349f34ea5d0020cf178e4ae1deb46b20b01216b1c460594cbe118c3f16318b8fd2800e7d20c0ae480c240fef0f1f3711c5792e3a85dbdb6359ad11be5c58ef08becab4e73675b02b99b653e3c5408ad600664b128e75a43b6fae11b96e6b2d4db9948d19c96eaae38c82ea1a40947e65e15b778f23d30c8e72f5f1904e0fe8a650846813a2c1874dfcb18c1a6b563b5c6a6e6ac8ea8d11b9647bab5ce1378df573255c185c486073d060729902743d06e7dbdbcd32c724f93fcd6fd4ad9565e73a0dc1357433c8490e3ca3e0ce203965b922cff26d4b7afc3339cdaa8ebb5b9144852c200cb8662d7e3689f910b187ac60fb880e4c7f6f34ae8eaff893a8985537916a4b4f67b69d08647d428afe7a5299a15ffa08c6a2ff43f350eff0c0a946dadb380f79a87f8883b3d2bab3ef3eb4de1ce77c87b6b74e23576af61af3478c150729d17f7f30088c411f0156b74ada99a5a76778a905782fb31259b7fedd41e0efcf9bdfc83fe0b92180d4d9d9ee76cd06bdeaba098e72a56ead97209afeb1f76729e77ada433ce5388f73206df46749b39c5db4bb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h1b530e9069edda4dbc32f312e33acf3df41e0d481a1342433950c19d3e141fc433463138972ccffc8268fd975e5e25db45f1ea752ba82d3c4bdc9e00f354a335789af78bdb43b13912e76326f16dbb8da2e9196d2be699d2f38dfdb9013fcba35c80778fa36ec6b8a78f40b20e6a5d34391eefb72aa67b86b548598ba01d249fca82b8be7e5c8214494c483af140df38c0bc04cee85ff13d15d50837c9aa03e440a3d93dadea6fffc8dde3260a83564f9f7cba98bdabf9e490f1a5701da777e9403c57edd4d52d38cfb6541bed2eadd04e034a61ee3d62237ae895a688f6762110848ad7abdd789920c329e0c5c9ee367c770743d1e162217d3964290554692216c8e4b9e862cbfd619140c599f81000e9ea91aeb0f0180ef809c4b0419bb408283c1de5adba5f6cd8c2c772dca1c5bb3b1ac52e87b27a716978873ac9ae59e1bc00beada57337a9d075c896beea67bb1c284324b06e5f869fe3fc36fb0f05dd8856fb9b2775f0b8977b5917bedfa5c3ad72f30f0f9dc836608f150f23da2fbcf50fac10a81e517bb7342d2d426f7b13b37085e1d8075d440199dfb212bd8b988e4efc0a9b7ff84c814f5773a8a4b022e68434c396a7d5752905c48c2b4a8a79996fd3df546f3f2b6f89b966060485fe148101ee092649a36c0e85023d5fec54dae1e383558071179904d5d34b19da1c5d70f919a2f99974d2c247efa7b5fd68e2238c12b64337b17c6458662bfe46ec6d3a4a0b08e603f1bcd329f20f298d07618bbef2766c701a920e8ae0d9423d2139e25734f87a25efcd3b260376d13b50f4dce14501f37727900e7afe2a8162ad159d708e105eafde68031c40c8b0bda0ab72f24d81d5566141d80c952cd9f4dd99b2c46943d61b91e93460addcaa80bed42e085a4af84cdab18dfa8b281ab1b9d14016934a2af3b3df2451b247912e012c4a190aa6bd528d365fcf7de6a1c793f9abb36a2c3ceb4c51b4cadc6f81897f65d89286973e113735f3d1119bff46f3398c4f54103977da2004297cfb307acfc01c9fd986fbe81e61d7a8c5231f23e10cb471ad1612aa61b18585e1e3b3cb05794e45c6575bc4fe76a02d6bb7980b3912052280210e1e60d0d380d5acb76a08c9b4689386126dca7bc5df95a28a04a3d99c20491273dc584a96d8b33cc3c4c85b328b74a8be081490a44a4d9362a6bc5877b508bb0b62350d1ae2b04702e44705b75f1c3daff7a46e58bd06b8ed1bd6f212c5b3213085774deec9d970b7f8af3602c1e8d378259804bf2285d653212ae1c3cb2c88fbfa42200db6240ce491eeca36b7d72764c538ff168691bb870fad0f3a19d9d810e05123b22441b4f3e9e97279ebba01f72255e740c14f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h8547076acca76c7da8d0f982040f6db8e9741e4668c99638b4a5813978893ab828db93fc77393ce1bd7685cd05229e62ccca6d2e07886d45d0aa138825558ea48b84af300318003e044a81020257245ce9c9c467c6a5bd27a8b561218aa10c25b58e2066f8c78d1495185cf6b15dbf20ec76c6f6988fe50d1af9a2e9c493ac52a5b8ab3f7300e4ac0cb11e8e82957b21db79a228628374d7055cef6a4fd490b2fc1a1588ec9ea3eef85bc4f7e26cc42d3e4d6d1ae6e56c1a9ee7e8d5151b3c17c80a9db0595a561c62344ccefd254e7250620fd77f8683a0ff4255aa64cb195672a56fd1599d023e8b1fb66e3bdde7969c75a7b233fddbf5bb427e7ba880e23cfd5bf20e588186faa4eb8f473340b8b89b83cc3ebb14570f69eaa05d3a76845f24236951a28858caad407099dbbb930019463f45e0470fe118e0f310601fa04fad35881388ead5531ab676e91d0a0731734abf57c77fece602918d058b3028784c16bf2b6875ec09560d5570630ad44aa4f238dcff0462cdf05b82608c3430b900f7a38847e748b971b56b917939d5f3cc71bcc99b3558c9344e6424bef79ac44658e1140a87ddb6fcca5cf8e92d4e0ab0ff1593b91e10624b91cce8ffb74c2a513e9ffe24d973cdf175635547cd9aacb8fed0f2c8fb07e7354e17b5a9db5b82113aab5f35059b27599681a429c001aaf7252af72eda84d61f2e83ac5c4ee1e7ed39877b9e6fa6245573cd17c06d25c047deab18f684ed90f3011866a2daeaefe71c598e5afbcc2de966121d0993573d445d586b5fd8630943817bcfdc2e6653420b696698a4e59f146064806634ae3eba1d0151ae68274940f7a2f4a433271a8d94175f6bcb34111d18a3a603374c326a2aabe9bc70d754e43b51a0c961adf3f35259ea57cc0891cf2f40abfac6f45447b88d3b23d0f15e283b493c7cad4791977a6f971a01e3f906ffd872d4bab052480e22f0990d4bb7197279bf8d6d15402aa812a230e15be283abff6c56c5413f2dbc7809f4f88b2c7f88e8c8d36977a7a230023cfe71103f276e9136b8309b5afeaa5f0c0d32e2d71a8fd3f66cfc2dd1d9e63695b81ec88b4cc257fae2cd44e79bfdc44d703ea0a2b5e908282d038dd68b40663f15e21daa08356f08566a2fb080384366d4aacbffffc8bd34fae5dcdbff3c0944741bb5968130d387d0db0891377611610cf52561a55d2db35b2620e9acdc42e72d77de27ba8d972dcc0f79a154774fce880e322a32a9cd2d0d123f33ed6b6204a5edc94ec51f8a19a6470cc55a696bcfedd49e438dfa2034c2dcb81d1eabf606653ee4e709120871958a16dac52962dcdc4352ed7e0567dc8181eb3aeb7eb4cc3f072dc719d412a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h2e32ac6d890a55503d0884831172efcfe3f69cc5ad5e2edcc4b21a39d0b56687f895b2db81d09026fea1a9a23fb55ac85c7e6d9a3a03c0f0e3f9ada635ce431d706e2ce82cd3c792e99032a8510ed268bff48e3520d0f70463f6406175607ef05419799309957291e7949656ef865ef82b0869f11160f69562aa6a657df8ae0e6431e4cd6abe967ace4dd642345a8a90c8c7cb41303ef908989b117723010d7626fc4bf42d169d19ab79e35fd4159e1ef52ba4afa7fc731054536f1058e6d7a2ca5dde3fa3fbf7fa4ec1f1e63faabc1a625d524b7ff2f4d35be715149497271859308ce3023708aa28d59f00b6529a98fe6dbad4b6e6ca0d928aea157d552b032c0217b7f009677e2524013d7529e028c70278d5352323aa43265d9b3723245af0164c8c8eb19527cc9369f1fc24ed4446b961ab39c59e2dab58512579d2150503f2cf9ac3103435ec8df11f76b9f68f618fd6f99d61f317bc9b1ba06687e76d832ed8a84a8b7df6350c1f5536ba71231c36fe7f6623c04d611a1edb22f23a70764de06ee2ce3130a2087f4f35ce559de693d8b5068b4ba39ae4b047c14e812a6dba50fd5588149fa04ce93def2709a4146f2aff34d089f6b210495a842a21ba5d7d23d284b67e360617eb66d50f751b13b422797078d57f8ecc056c2fc6b849bfc647e7b01d940855b17959136b3cab060a977a1ab6d7de81a050b08280ddeaee54fe399cb0b4ff45da4ad870c7f7146ad10d1d1dcfc029a33187ad120fde8d4292b2ce54ae638b62080afa2e996702e8f893a8ae14a97d31b68d0c8e1567dffd4135595e47a9944fb23f46a7db279c67dea02210203f2d8c57056ff043947eaa6a5b74aa4ea0f03f70cac1a6a84501727f04cf77b4daa918360afdbb28ded7f87d20cab2277494cc9135445d3b765818454be5ea006fad0f486afff6226ba9afe49b4dee60960d8a3f9300d4cf55a07b458e9c8e2e82ad46471d226f5602226a4f56ce58af86b66f6fc569ba6d8c225bea17a853412e3929ddc95c1c3db9555aa1b39be6756e2043f048420d60cd275b87c6d8e30f09a64413eecaea12bbe22b05edd335e53ee6ecfcc522880eb4ab3a12574ca4c3825879f6f8d4e087612f52a18fef83f887eeaf3e608d4c3d913de08a1b18d14e3dd5d23560e124ba314288f6145e42f6fcc6e09e1a496301c6e04de4c5766f4cd2edef576cf120490b997e2bf4d96cdfd4a020ab08dfab3364a6fc9098d23506f5eb241b6ecb288aadef8f0d6b1716925581db62c33db785b16a259ca4817d6285b988e7ded77a0cd267f2e4da7479d0e48fdd534a4b3221f96958ccb793462560de382a6e3a20de97cf22b4e35a5de0c28d492e829a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h8a15a547b8d2bd8aa980733a619bb8984a68dc304c83df48912fd1b875cb8de0efbb786d74ae7fedc275acfd3ff9fd5c179aeb6a05a6ba9007ad4fa5975f8da9a4f7301a8d7cf6b5f78d43ae1e22d6e47dfa247f9fb5c1a07ddcf880c28ab4f36224ee4f1f756e97255b41be5c945bd77a792bcf7d80a886e3ae1d2235ed8852631e6f3158855c123a8bac5484d34090100f513bc0124c07e07a700d1699e6906308ff3bd270a7042ca4e08f8d9ad39583035f2f33eba48df3b04d3e5db0915536df6b12f14599f2f056ff1c67685a5fe73c03135106dcc12696986f8abb9803855507cbc37c5bb377d8a1686b473a4f2b829d0d612eaa712e448525971bf396df114e503d62deb56f501d8ca936d9e1730361bed7a6e059312f89ab28707820baaf832642a514195ab4f224718105840eddea8a03ff4a09374860f1165aeafdc9a74f4168d6694528a3aa75d09b9bb8470c4eabfadf63e0c01047b99d1391ae899e53cf9fab88451b9153d5061b0f12bd02889c7741123cebcd1c9b7329baa7781834b1cebaa387da6bde314e2025863c31188fd2ba7ccdd907dedfcfa2d40fbf4525353de7f862460e7ad6ec790ce7359b16027c62606b524e55d66ef845eb1f9497ae8997a645fbbf7393b4e6385df234bd6f3d7f2dc7f7bbc66896d06f0d0e7a6c2a4654a133a8d88e0f76fb4c714f6c805dde66e9f75f248ff60646487ce37d395a25cfd02cb7c27248268fd7b0565c14e27e33f263a6fd45da74ef15eabbdd16579f86f4faf815a7e2d99fc359e97cee626beea8e2d35346525a9d16494d70c738dc2c0b15c82aaa6a9c56dada788e1ba89d8155f61c18db8a411c18b52cfb813e32733cc30bb9f738903b0d59d329dc2dee408825bdf3117308bcbbd0e43872b399af0b0c0813d4a58873d5bbd5ae04a5b6fe7b4081bf2303233ba03a5c18613e84367194994fc23499420fbc95a340ec6651ffbdc54f0d7a28fb4031b6e68665ac65312a5def99f96d030990856872d8b8d80b46207fc0edc82558668741d39ead7a394d89eaec38f6c5e96272e5393d65cdddd09aea7e1f158e67d050be737b6eb62846e3da5a4e2350a5ee44c7ae54f41aea9d60e87d30215703cdffc4909b5a9e93e04bf2477b396b43994cc6985ed74569330a2f3090ad7b6c29e1d7173e653609e98e8c6b5b3800b3cc2269d38e918c2f2b2cdb6d4992afd865e5d9075a1667bf96323ea88dbfd2c47b4ae79833fb8153cc9dcd23d7ca73caaeae06a3eaf50a6cd03f77f388ac7695119e73fd9736e092fbd99383a6900f75fb2f3723a7e4a664ef3c377226b2e5d997e48b2be9497aa535c2d2fcc398b5571490ce9660a2a612353b2ffc41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hdaec0f6cfdc94ca236197297889392521f5f0e7c124170196616e5e49036d1d9165fd5a42442241a14f7c04159fed8be2d896d42c6137c057635521653be2a69ebd6bed0422455e138942d0772eff2b0537dd949586726f8115b56f17995d0a7d89930a4fe167121ccf0a9497bd88bb3340aceb534faecd8f77c43c56f168eaeba10dcc21bee7e50f5a7c5978ac904f8416f4703ec59d4183bac314ecc44b56ee23a17e47c9a1af0aaca302e77c1b6a943d57a58195739af9ca152e3969f66f7797f2661707b09ba814d4dc42466e51afe40ab030f92e54d36671a0754c8120823d1678c90610366ff55f154936a22134fe3a5ffddd8f454f1ef6f169e7c95110eddd44cc9573db86ff8e375581658252ca124f01a3ab9ecc05d4e5b8a8e55327f90a2af8b0ea3ce12fb254396e95b7f31672a36eca57a412616f447a2fc972733f85840afa3cbd071f12d55487d5c8d849e74932863f93e2256ea3c6d2027a2578ad6854128aa127025b8fd2dff32730eba73bb2d8e97b2a0af158808370d58fe119a0fdbdd90233726185f2aa58b769f64ebe8362a10817dd0a402454c5c6c339efc2b30b3b85ac53374ac9e6a99a385ef46331c93ab48491862a374d4fbb4804eb7776bd8bb14006a077f97a5bd889c8d45b15924fa3578a1cfabe5371a569beed787c9c1049643c7c99bf6491d223f45069f36d7c721035f653ebeb55b8ea800eac9e47e89b076c1aa08a17cb924b17e60ef2b98ed47400f62a846a8247ce100f17c1f2de06f636a151358749a83c2bcb09164f1f1530d295b47b381c73efeba540025a8a8577aae09fe638c7dfa7dedfb7acb6a224aa4159ac40053c8f1759ba4fa0454794e930bc36eddaf128ebda72b136fcfc4d35fa80b7108d94152cf43c38fdfe6a6baf7a1c8e8b5efb8e46c1f9fdf7ec28be55e41c8d57f476487db03f1fdedb4020a148d2ba6bfb465e9054372e5ac581523d4c4a373ddf1c5003bc5c476743e1778d4c4b7a729c97bb3ec143ceb2315010faaeea7c150d67a3a7d973abe9dd21d47fe666767799d9b39e2a2bdf5bba9755d5bfdeeeedaa937d4ee8dec7cc7e759e8e9b4fbb965ccf97b59c3cac6961d32f4569d0734bdb4eb14615c9877813327728f6759216ccad37e600de4b6bcdca90d32408c3262df3ab4ae1d898aa7cc0f267e71a93720fd1c78f74bb4142973017961fb925b2a2893de2cca7595efdfaf26c8a6c58f0f00c4611755b10794c6e011a4d83e99b56127bb1b60f58389afee23cab7ebb0b710b6da0577894df35dd64800f9f6b11b0cfbe6341b84f9c1d7ac6cde474cae895d5f7076770d7ecbccb3afcd9d43627754886f622ca92200d99e806d8e2895;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hba97512b47e8e3400aa235341fd37d1aec2b1a1a0de425948349a62518af224c9f0c42449b61e2d10c6ec5bd83d829a29bac130f02677fc2306d21aa672e3d3c46d876335f33eb1b752dc3742b172ff6e1516949c90f0312f1f3892618ab91c59fb0064e3ce362dc8c4ee16a146e23775b81bf7bc930e8423f0ea1b41a6b91b7d1b4e3915ccea40a84834844f5d2d5a5e26a6e2e4b9ad9fb2467e2ac92f11506d1bcab23daeac59f44ed2b0f5e42bf6d2f72f6b846de9b4164056316c712426ed8472f8d0056cfbd9f877283faa0b1f716680830912480d3b170fc8ae16a22ed097fb9b97ff0563c7f295b29c08337e05e0fa6c72f9212f2048611d6f91aecc1df1d401275ff2a74cc5ac09828d2d9e903211aea59476bfcc6c594a083335fd6e8b8e36fdc776a4909dcd1123735db30fd7116737de001f5048342ef204fd58192e859d366325861a3000ea3bd0f8549bf2455eeb29f33f327769c60cf82e6fee441be182369c964e9f02271b37813001b79261dc6230f6b3638a6cec298b24cf8c8801fdd3e3a0d331bb39d5628f2f647e939362b33c6dd7b26ce9af447510aa5e91405c8199c88c9c4b067dbed9e8395760750a86f15000eefbc19a8a30113e5181e74b6188e7f477cfda8b787cf235c816c9636753555510080189af286ab0e2cba19aba8f3ccd84a8e4f0fbd781d962792876dd3ce8129e4a3aba35b79ebf776a869a328d115b986e703a1b3521ecdd7c0f598e436fdfea3e88091fbbe0ce01f9908950cf03d1e82a7fc42404205c1d31ca48ee8416d81fda70440175aa51ff4a4a296e4ccfabe56e48b728101fd8b96b0417e1004465768dc9730d6385bcf42bfb70d01089379ee385f358d48a5dd083af89be0a4c8366203fb097e02b0666fe6bf75b56e9c8122e3000d786147e186ca486b614870b4ba6d60f1d1a695c51ccd10b13db98b808df7666661eb257d825737ce063ffef003778bfe249340f98c02cd5d500d79bfd5a24b7b6750fff38404306f2e4478c9d27b7ddff4ad4fcc70470ba7172e3ed9ccb7f10f4e63ff9e0b862406bae5710455be2b11ae0e2def82aa8c73cc37a47658c2bf641dfee7027ab337f2a3537b29e7fba9b6edc169b297d8fab24715d44cbfb7cf1b5bf2afd53f8a1e2e889b8031e81b38cf79bed4fe91d6699b12ec88db13d11911904ba5bd15e9b9790aa7a00513298609a2bad04e6293d38336b8a3876edee010dfeed0fdda644e8ff921653651bf18a070ff19095b0dc8c40eaa1128131a030c4eecb56ea3880b8f1acc5e610d22d77c1989097d7f7eeca80ad1b9ebef865f10a40d104f7f71add7a03d8892f0ac91665c03544cc02e6e48577626292161f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hcc487d0c93a56e05043b0b1505013c0f472fac2392b75eee5415cfe7f4b762f7fc0e22db4b13843111289e1cd0af8207e8c82c328b389a1da2e8813b0098ffec91db3c1da476421b3397928f3cf9c691435e8868c74bbb9731c94d6a3c7d5511c5a09e09c9889a7b6617373bef85ad21af8bdbb0c428128b309743fd3fe5607233bbb1126aa2e64d65ddb19c79e37ecd068b58f6a5a389df90e0a06afad58f8490e3ee662df835357964472e8f40a1ae72eece0e9206aaf22656a9045b47876d19cad4f8d627e69e4f04f0eec60c8866ae7e5ab4930a9ca065520e3541ee542606edfbe3d59982482127784aafbaac6c08e0fa331a0fd9dbc9550290c0bf92ac6438bae4b26d629e8cb40a57be3e471f12c16f1ead50ff42d73dc14dd38d44c46cf67b8c352c9121630a98ce471c014d7ec047ce34130b83a19ce7e00d600f7f42689758c5bab91475b91955f1ccfbd069b1f7885c0d8ce6e8e14105f788fbea1811b4c1d518a93694a96783fbe3d8d1f7b5b4c88a3d1fbd9fede5595c9e8fe01eb511cf066a36ae54c7b023f6f023cd961379cc97b6a550139239566bdf209cf21b1368c4c698b5698b5097feb46d4501b0fd30b95c6cc721a42ca63d133a8ea19581dffda7393ce032665e4a512a0cca7acb4823be6426198b6fb80d9ab6221443ab865ca85f791773a1893a36cee525799ea2fa665fcec6b60df28e9d600aa8332ea43c71e342602569c1bb917d01aed0e537eaba47932f64cc46abc2967883e31d79092393998a1b40ccb3336d3a8a3a244a08dc0b535b4c30516985f6f04c99740eeabf0ac7c4b70891ca160588ce075a7b8fa9f87568625c26b1d00d9e56d1bc740207067994ce447df28ef89a2de60428c40371b9a656ee7b2906a566b8a53dc15e6804b507bc09d3a72520989155a2e3a174058858a5d1637f70c5d43a3803982aea0eb28bf14cd5b7ef14c17ace5f089296ae51b29ab19b4c3b42049d785bb85f630b5f6b3543845fd014d1c7a168520e7a31f9dae0e65c6efa743d860be86b05ea2a2caf404db500bb500194b3529e6c25a63895ca0d1e07bf97f4ee96a1239686724215f1a974f25930abb858a41201794e2ae1e814f976000e0aba84c16d536db3cba11c17e64490ca0aa270862b3579b7da76af904b37970b69766ff3189bb5a77ae048c8043de81b4e4f9e76d1b970cae979c0648714011e546195e4e817be0bfaa98eb7ac6aae17dd1f587e60086d9af3124b4097606c332bf6528a4f0042505180c8c4281d5b98f173cc321136c0309489ed5a1a88ad66804b7f1fbdb98305604e35f32a5aa786213694bf3f40af5b556c738d3f7d97f28ba5f524b5229adc46ff980083;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h4a0fab4b6f4bcb930a0c28c19b83f548addad9d31b62a8af5914ba98aa25e1794bff7f69931fe491140b7fb39a26214120f146f9928ef55e4321ddcd376f3a7c77964316156324e3b4e012acb2f0a341614931ea473878662b8211a66023c0a4a25eec9bd2eaae171e18ede2e8b3c372645965eab06a349bbdc43d5728af4510445958b0021f107c94eac05de3fd98321c3b3ab3e053c45c372c71b6f88008d6692ea7c6b672e90c02364df4281a39c1c9c13bc11e98329a1b9bc49486eae3b7fcca8c551260ea2d27d39d71ece43720ae0585133aae16b6cd7013e710132ad8f6d50d1b9147c0cceac9ff10b386de519a0a916cf1d8760e369b8c734ba4214e7b2d063b044026af3b42721f3219bdc2f09ee2b4b21dc3acb46a3e4213564bd5dacf1bfb2d21bc79e0784e0f0e7381cc9d4b9e234aa38dc3e46c7ac3dbdd8eb43ff3ec2bf8f11e4c51474986449492a5e14aeac30147779b25f8c9564216459e712668bd0749ed9203b456f44407bbc4aaf1e279b78986fb17d85e06d799e7703ba48c019c768a7d52499da576dc7aa0b99a1fb7402a42060912e2987f694ef994cf803efc5de7fd852e48409e2a19dc7b0050f7851d7625708d74cc1d966e40390bc73b802ce2e1b826c64225b1a78c81e940b172ec33f09b266430c064477813346f0cf663a4cd9aac910bdf93a789dec66ae26672430b298d76110a5de4873fdb112c7038787ac42b0efe57b010dab9c584dec145649f74f36b4ed10800e469bb70553d5ae48414d4f4a80e0bcd2c40b27292dd31630768bd4ea409f306d823e22b7d8da3219aa91bc6d60e89caf05d95b0dd51ba11022d6e66b4d51562c04464e4aff1e1264b1a0c3ae0645ee39643c5d51b3939340dc1e2e381ed57efe6faaae0549d48fb66c2eea357044a6545bf44184712f41c7df3ec66cd1b86fa6e53be13acd87f167d4e96891fcd6047ad8ed28f0ee55dd8ac86249a75fdbae0c7ba6d685b86e8628a8f70c7651beab80ee0f51f289823bc5e23d0de8bf762ea60aaff06894044351912310e82e041a61e6f917ddeaf2ff9cd4a36e1cf1bd5657063c94934daa95e9f923c37eba494a2bb0dec2f51ba3621fa288bb51a8694094e2baeda4eb748b1d3498e6bcdede98df60638fd1d087bd6b392e71ae06eb998afdf9e8f4231cee6da54b180878b19076e792b55f32064b42b7f2ea778ecf0867dccd8e880acaef4a1861ba892b22e7132f8171c763ab8ff009979916669e1092ad30b26e6f7400308fd22c7f201ecae41ae644a66b6de70c825401dbff9cdf8a3b7b1f7c104676793655d75b121b560829a8eee0b477e4fb3853145c20eedaec619fc59bf2f3925d5870148e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h4d2db8b9311e19d7038eacdebb6cea908979c66b2aa05c3e141e62205e81572072c8a899d7412f568ef9d8b6ab6621b4c4974679473da022b8886c3846bff6e63d78bdee3eeac7db0c6bb96ed82da8278eff6b023f285bcef8df3c5c74feab955455e0b6d1027d6b8b7a82dfaa4d8c7523a2ffc82d0eab5da413bb5397035be0ceed6918755ad5e76909ecb4018575e890c17bd09045b4fd96ec346912703c04f3e60c50411606f3beb83a80948813a2b14abddee1ef84da258631138cb56079e0200032d151140f31255c99414bff474efee7ecc2110f293c77418d29427b1bc73c3dbd88bef36114c9b29394ecbe4679b653bd42c65d0251339b4ae40dedf0b00d52020083b5a1fc6d936f73e80aa6c040cd57367af997179e34f14ebd8de4e5fe60ac1330c3e3efd85a60ae0746e103e82019c218f8734feaf3d1dd04962f16343bc9fa630c270f08063768d1ac95d71e0af178c244b147aedffdbfcebfe95d6e01c3febdc883e78096b1d7f7e028e3153c861a48455bacc8e3cb5c0f05e25ff3052aa68e1445f7251d703904aa0581c89eff98c35c25e45863aa43393337df1eedab34795a47621b73ffdf6b07312567c196e0bea87d7c1cf99b60fea8fc732d8457a9485cb68b9d9363f3839545e8867c70fe69d4873ca5f9268569cb34d281d28c55bc86ac75dd03db5805d91c33ba6297975324ad4fd862fdffd0505d28ccffd7b9746a8a9eae269ea1d0a888ff5604257f634b9438666d66782d3ac6a0e3bd838c4d7092ad9ba913967aeb2f092cf0e2e6fbe2ca2985ca7f5ecf4e135d1d62edc5500cfbb03c419cc28af4f7f8ee9f1df329612904fe0a681db46b1909e4c906861152749456919c6efd109e20200c032ff39e9a6f5093375929f41c995ad5d2d9a602da5a443fe35e23b5ffc68f73e26cfacb8408aa3a7e23cb370f95075f063bdb1198cfdc74f6a0d2f1b43e13be03e4a3054dc98c8e4ba18eb681a217dc1460a852e17295892d8feeebf978350799c8c98d9fc819fdf2d6e7ff57a0acd87bf9164fd7106ec007e92031f4fdeb733086114e4576c90d6ac7f8d9fee9ac5a8802f0de534e4c6f4f26d031370d981575aa4a215b00b72c24821c65a463173fa150b3f1076006f5135b543e13acdf23794fd600eff9b3c46c327b2de163f197836b519b1a477e33c5cf0b83bf31448694c1b61526c90093f99643bdf7c95a76abc5a3c58f31eeabcf22f6d14ddffc0b613283ed544dc759c4a09728a3dcd7e005252aac3c25b7d66228c90acd9f4decc3fb930e71a9b14f82869acda18f939259a87b108b785f6d5672838fca481df315f9264575f682c713719ac4b545d068e4639c27bb0dc41fee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb6be0044b463333924c4cd2ede988a520e576556d73b219f6c01a5848d1637c2c06cb611ec49f0faa9f50424a5b5110454da05d61a77913c5e2aa41ff16051c021c3f6503035c5d6dcc70582e1edce5183b7c511bc15508dd3445b6e0556e04b539aeb44a10e17883171ae68df1c54cd26bce00e23977eb41e96d9d9e6fc0edbfef6649c2b3c40e777747743a0c90af211a6572cf0111c4c6519c074261571af3ff1ffdf59fe9b2783e326c02d170d540012af7be5a3dc243827918835e1cf468b0649febd5a0ef96e18861e4b97353bf8598d612210d27e6372cd1c31159d59601c4e92e7805526cf6823aec4631ec5f74b2a0762b7f3f81742519edba62d51b44f76a3493ca10168739438a78d81df098b55f02e6a253357e56dc00fd753d36ae7cf35ab2c58aee69a610bf6a97282840854a9a5346ba0d4620d2d8da7f92fcbbf6cf2a785593e946e9f80923a8106eb63faee20b8f3fbbf782cfe9d7e86b7a5206d77f1f94b6d389f8d35a8f30821ae4756d3bd5f3a3fbc6ec31405b4007990537901679ca32382231391aeb9588af4f154be2cac1eab3e932f8430f098fb5515cb665dc70cdb26ac4f8d91bc16ea63ec5592210a925ba53d69ba37f493d6786a6c528e05f0dcff167a6565a22e752a46cc26a260e0c54fa195212dc20396f9fc104ab85b7699b6ff843071ccdf509183503a84bb0505dcac18b3916154649f74545798d1f6270448e9e4f982070da5ff196183b8e9886f879b96476f048f630db3fb395ba98e1c7a0f3b29081521fffc8b5b52bd333b142c38c570caf3109fcad7fd82fc3bbca5d61e5265584de7dc5844e51b6dc936a4d106dd2e0eca2e36b5095e16ea096531f151675ab12956c6e4bcbf321914edcad78528b2f981f7238f42586c57ef26f049cc5b622b4812689b3a9d109d81d49179cd464676352cbcdc486b58344c08c46c2ccfea70874e531047e3f8e4e52e41db204c89c88fa3f7dcb955315b3bcd0486bb8b6a8e3e11173c7c2cf01d29987e9d353c08b4d2919238623007aaee2770cae9b4c42579f0ce41e2dac6d99a744b18b380da050bc75f1ef6d956365fd26685285ed8b70501ed5586abd792013a934169e0a8d0a3773299649f66c12ee353c2eec4fd66260590c089f976fb92994de69f2f12c3c93358b087db7cce3321c0406375b7a9b6fdcb8162ae17c41d3179cfce7968a976b37138a54c8c79387f009bae9529730460ba987eb9c7102a6e093851098ac78a465c13abecb41256d9321bb5249c8989ef7d415225a94dd2853c7f9bd896f4286699bd432af2cb328c4fa9e2e2673e8e5c9630e978e7364083ab42b5f9d3ada628a57e72a4b65bbd7b3157c4ef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h653786e5b0ede482925c613295458d3633cf911c7c370758524ba7a018052cb6b0ac4a02edd88e0b77e0e4c4bbd0980c0d4eef5ecc6344e177784887d648016bee3d4fe59d8c08ac801b9fa21433b5a3d74f41b1d15ab1e453a7e47353247d07f3e910846947d4c2c4d7484bcb31ccf4fa04fd07c85cd8177addc0bba3be47bcc9327f6ff61007ab47679b672ec26bf6d2ad63d49acf01af688f90363fb294f7fea9d683c56006fe18517361748d2fd4f91faeac164912870574aaf7acbcc7bb539ad6b5a0bf13513f5ebf59b7d405f300a58d5671b839163be96ae125ed23ed5b3d903c5a4243c320f0985bf14409ff6cd23482f1874c319efcbbc8cdacda1dc1aa3ff3ec653fc7390e8ea0a22c98eaa6c0b98500305ded7042e07eff1ed012af7bce83c7446d0922e15d67afc6bbd42b8063adc67936452cc26ab81ea712c8fd94414277c36c51708c707d6a64bad44aa6f477767b030bcc7a0b55f6b7a65cbc25c137608eed3496c64f5c916efeef15e47e5e005761674013035109be088ae5035051c22d7683fc55aee54d2b0a1fb6540a506cc982c89a9baba7cccd5d9ea4d6987b092d9374c59c3bafbd125c7e9d84e1568ec1ae6f27f9dc8bdc57a73bd30997b55aed1658109ecb611cfc781482d78cfd2486037871f988d6c9110da19c73a39561b2c8910f77c66fef67cc1d638b793166eb6636468f6c22cc054a9dd278e7f6bc84280023b77fc4b13c89069bdfadf1c86e1e9a998218adc2ddbebe2a9d982f6f96083870ec0d42e25c6bd5a3475d2bb887b2b85df718fc006247b1d120cb418dbe98baed6391a1ed54636a1f36d265cb40696b562819eaed233c20bd3dbdc35a6b393e611ba15ba121f60e11076fa0bb58a42253f34ec0f19a00d74bae3c61b51b2c6621c05716d6d06fd62d87b408fec52cad6de392e1e5c72e054b83d03bf19011a4e834055890642f270a6310f321d603d4738bf4415d18714a8f9e993d6391741b4a089b29f7c9c4aadb9de6af89c668d8be5354aed63661bd11a26ffe4e8fb051938c7d2fcd56a33d1cdf5db16ebe7aa7c06b1328e26974f32e9176797fb390d24297eec74f020dbf03084893fabd10058132c4f939e20c6f5c289723e00648ca3393cd73a11c705998b0973c05b7741ddd9cd16bf15cb7ddec892539f03c303bbb9e328d345b1aac35491004a69baa14fba517143e76413c9cc56c928f1329064729e1f0baf0b5610bd524f72f30b48aee1a290e803bce5286441ceabfea70863f3827c78779c5728d85eadb12a253d67dc0a4dea2230978bf64eef8ccd43822d983160e011770f9a6877580dd6bcf76c730eec6223d7e4436d688784c1a19774ac85378;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hebffe116c11f834b633346bb3812027e7a7a2eff66024fa16648cedd9efe2b5b6f2f98fe763f7198566bfee6a091fac186447a45a0f45600e9b71b863feb53f2f481bf1e3b7bffee2f4ed175fd0a2946b6b3f1d0f825e07e1c844e36797229a8ff639a20cbc2f26613d67717c38aa6b84c870659aeae0b98a8677fe9cd2e8de54db1fff09d86377124683fe103ec39a2928921f2ffcf6fb27bb3d95064c54f10f15859f9eec4353994ddff6d03054425b6176aaf49d5f3a477269737f70bb0881d014be03684623e9979e7c48851b4ab6cb1a5a72387e3eef98cc5c8a7dd93a5e64ed58c44ede6c52b00611e3a4254b01eeb9193dfea3de0b6653b756f8fdb992a9987a2f857c1391d4ef85fb285c3d589e465b07df70e1ed0aa5505eb17b77c96242c2848a29a4525e6d6f43b8bb0086c487e3ce41ca68e510f920ee47262d09563b416001eb1c3354fd2f4b322a4daf326da5a4937ffc5dcca33f2ea17dadeecaf5d6a35d144b250b1a565659a73443ecd2cbe20261de734f176108482cf81f4ed2f60f378f8089966b52995fa90f7217d8f12c2b2ea7a7fc171aec28b92a7fcf9d912bf84d188b504001f243925c0fd0ae5c11f3754c67120453fd09d7e3b84b2992d1fa5a6cf8df525351346a2df3c3dcc14f884a994de58b3ebdfa3297736efa8e161071e39e0541beea239b939fdc70e07e273a65ba2d14c9d5bcb760952c285e2a5213e4129fd7d6b7b29cf9288da548b4b0cf648f1e08e36d3bded08ec439be54a80e0ac3feb4dd009c44db5c4b2bed603c4217904cde39dfe447a45269f358eba122ea55830f29fd5b6ee00b203d624bccc0c9bb59f7c793276cf7e52d1bdffb90588dfcaed656d4180f3fcfb9b1e02391d3fbf0c79b20fb0528a36c91f0cd797d502e779e036891b084ca615ecc650b62171f7c461fbb822c6d2611d54d509e9cd7dd9da065636daf295c7e8f43c28f96ba09ce12df76af08527c7439dce63b645f26e920ae30c0d71ec501f8864801a56f6dd4006f9f23981d6b0bef81e6557325638556d2dfa17dac450327f9c324e5a699bfc141996b3e3ef7545948eee90c0249dd2191c67f9ab46f1373621033661b97b931da0ff07b2a2fe31c13497a5c6828727a56090e8edf0b0d219d771fceeca8a1198d5145b97f1916394a0629b76865f0bd3ec08d36e7d7ead15ea5563e8e13454d0d0a8d4e6fa2d837d0e22417e74eeb5364e12216406faeb38887151a20589b12729de8c56a43ad1881460ebbb1ea339862f7788b808c1a6354cac14ecdad1b44ce2ee6fae7a18e3dc0f433120a8b67130f39f299f6e841d6a4d202251352cfc016d243abd55c858c83304b875544b69f2cc37;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h190898d7b6003de73f626e6467113013751876a158451b718ddd94cfccd89ee98ede43ab07f9d2a42e90370eaf0b7331d01e0a71e2947a647054403f422a94911be3eacddfefd11d7f0687567d09f8fb896e05cb6ad4122dce26c89bc9264518050acaf7d50a81b2cc3a97896fd086bb06abe6fef53dc16f550c72b939c8af150c1a5cfd9a945136f681aa707b4bae9e007f5e04ae52461d0e6c907cd60c554c48ef17c9af7ae7cbc4ea8f5a380fa4bd5a502862bd71c2003dff0258d990928971a184de2a87b676738a74c2448d7a3e4378acfa769a417cf6001d455bddd91be76424c5bcb074640b6d53059bf3ce5e6e5b6d8d6e954ce72df9557afb22cb2cf92f97cac8b2c391847f6625266d6d0ab51f473e08c5a03252c819058973abf102b64af316544247c06b19b7079aa9c4059bbc1b7b0053c244e46333000f0a18a20ec7e9128964b7a2246244a7ae227ac7fac6246bd11bf57793d7ed48808f0285229b961ccfb9a63bc0f423b468c6d3a1364df14fccfe809298cd107d23781b7b407cad69f983e02ab40e6b5a4f4083479bd9e374e77dfa693902d037bff363bb71652221d2a8da9c4a57acceb5d2813dcfe275fc65e7c409b30d423567753d4038a94b84c473a89ea461ee134ef13a77e26a9c0a355908db4c7867c397273d51b0f487978fe6b3a375d79226870e6de7f38c82125eaf685deefa09f0771d78589b1eb86e17c8d752484b8b7690c9dfdc9a52f5046d3d9126a02507f6298e1580b10556fc551c7a9f9288ed961ed7e474dbbbf1ce34515fe2242bc46010d6331ceb5897e4151ebbced54b8646c9ea19407b5ffb8bb9749127a951c33ee611c2f8044503ab0904ef18f9d3429cffa4cc541e969e237692d2d7a8893bc4c13bc22a830a407153ae32cc840fff7ac0a985b319b3be1219b47a8bbfd2aea0f2c04393634003b67dee5d8d6652032400ce0ea9316a7913aaef3c18452ac5ac33b861ba93c8e1069f035905a8d43135779accd71dfe2b47266fffacfbcd822934d8f2c0cb7de2118ce7ee65a5cbbf94f54304b260fa6323561471ae85f4e407a81702fd4756056af9b3c9572e7682fa637852b00b7d712fc7acc7007b514d530155a6cb3c553eabfe4dfc76ee01b075cec32bea6d6f72acf0f51d5538d1f97a5380f38a756235d13460cc4bd88c58c9119b0c69dfefd295872de0e53c3cd94d9d33781a8ec31a5a024f2988439cd4d5bf44f95fd44aa4eb43c725febdd2610e1368dd151d52da590d92654ad53d6e91cb88ea8dc90f18b00c1111637345f713f1c373fb02f5dd3a87a65c82814aff03c0de31d543f9cea457c85c1d3496829b6ccc3bf310a998e78a04d5dea378ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h49260ec9aa1e8847a688b34c0a7103ff911d2c2313209548a66578cd356c87aa7d26ddaec24f2e9fc24174254eca2657ba01d1259aa06e0e9c478d5b5f8a68cbf65c255b7e8df01a0a403171a5799689524bfcc266f30e608a681e4fb1dd2707748e3e24f4e7e66dcdc0e26a574e21414503a0c8ba80198367c3c8cefff97bcdf150346e67e35caa5b613b6b9ff882f2258cc3a7aa092b5861253b7b0a9276660d178067e4c73cc6317f0a901869759301532b9df93fb02a443950432b4e90592806730e4a95d43ae33fc6efd61536458467980661565211fb6b9a5cab0aaeacc0fb253e27f0d642deac27e1c65bd68f74bbda5410301d1d5c9eed833255cfaeb0a59dcdec2a260fe624786cd15e948b27a187700c291315cfee8cf082b8345207a360be767a8848f8d315bda09466cc42ff958f0fedd168d5b5ba01309c55ed37eeda953bb62d524d2e09a756b6c3b1b0bd472f9dce1995d8bcc49cbdb6e5d139a9ad90643243d3de87065cb765517f6d326a90d316862170a3931665dd51c31024622b3edd9607e1d3e2d7837d9c72b6998c860799cf81ee581d02d98a5c796b9d53b66d942be984a2371644d9b0006a0b250de63ffbe700ac0544d01063695f6d4832496ce7115f753729c1ea74ec70bd07ed795a184e733e5bf238fe273f6d4b82a2cce2fac9cac0a0ebccf21d6e1a2234d15c8958917b575566b625947566bfb05c16d8cb0bcabd4e6f05244e8a1bb7b6639859dacd6c40a31c9ef8883502ae3126b76c183afd9389345b200781c39e7442b4a8d605650d866b4115c0a19958f3d93717066de162e8cd62b0a7ff4db7ee5b1fe4fefe0aa44c70088de9761d0a306626f6fc72016ccdfe4ce5542ccc479238fb6518be053376e8355267de67b9c25a35c6e9a37fcd76f19a6dc86526df979e72a18cf44e5c1b81eba013326a3d77a3990df25342569290316f7f95f6c94233fef22ae05b393b2e12e7e0d9a87095d72fd66e4f22ee19243456567cdb477607c10128d6d60a4a5b9d2dfd6c22a08185f2a01d9542b2d10a26a728373854eea2cfb86508ea64f4968fcbf9c0c938c04567926c077e0597754dd83f818e3df0ef6ae7fe83321bb8b2742bd7808b9365489cedebf10aecd846d3aecf9e721eb3c53f6709ea5458aab6ffbb54530ea2ecaaf9d3c0cb8e5cefd4bdd9eaffc536c9912e1e869a71b3cb4c3d8f6b54f25408ee6a04e6e206d9f59a8d3fa8beb59be7e01b032a1bf271af455913319965f005075ebc912348e177d5f03c40f52625b33a98f1c4d4eacb470d134b8f1d4dafb9964fbf327fef4b69f4f921ab451e9aaffe274fb07fac86684ded79d00d4a228e7cea11e91a33989ec0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h1335b0d6cf905a8ae6890245c96a65697eef72a61e99f127fc9be9aa8e90205ced906fdb30e007f74b51c182135976c35421581c9d4b2114cd0e88efb91054062a09937b4742e8164587541ca92c7efb35c16558ea376f12b5ccaeefef7f06e7017a846363209e5cf2eceaa94e2092dfd23ebf8a3620f5f06b788264e0a099c478ae5356c7e9d5894fd04d2537549821d521b23cf1ff3fcdfe8508a1d0e3697cd4f9ff542965e60f04623ac45ed1121625903752a9ced2560cf543d7349b0bde83e57fe996a2fb4f81c37c681d2c9aeca813198ce9809a271d69f1febad70081a6b1766bb84cdac69fe9ef760e42836589697dd51df109f4a73729a65bf2a739bf66a0de7c69e81596f90fc2b9424eaed907975224b7378ddc05782e3956986a84394a81ec84477168eb414fa6dbfc6695d84f03bf86c79af843e76536788b13fa8469aa935674cfb15bb5d782e92027e8139bad3c4f60613ae99aca0ed0c3cd59b97fd911fb0bc9bf15c1719270e1d9ca977c16f94c7252092f9295383e732127ed1df64d18282fcf0fc4c384075027e2b1f558b1e5682f55e4846cd341e17d2843976c2ce1b773c10513fe272c79d41d06c58808d58d5cb7a52be4533508ef823c63b93c969bdfa88969617f3289d6405d902d0f7d7f2deb23897593fb3f0bd99e6b8ff432329bc3829b595e0304fbd17f7d5d75d39fec55ab8d106200634694d5af136cba731409066b51a8fb2804c1f761d1f30300e66fe5ea281d58ebf084249717af0dc82a074522be7bfde3ddfee8be72c20b901e3b58d1ca19b7d2efc4a9414517a0f3d3b061fdb42e9465ebff8743a0357dde2bc4b2901b7063307453063623b0dd8d978617e37493b6c7e914e9d019c1c49a4eecc574f8e0aa966afccfd282e89fdebbaf4a1c1b38e3f2e1e59d801b206d57ca0b4509d2a50b12da35289e65494c53fdab19c3117dc7a7c18703b6e6c94a497c09b7d4f195c5a3366134d7c1c81798c03f1b240bd2c6bb0b6d60ae90f300b503211bb030aeeb48030ea23a6ce9b02984381848bb1c096d4478cea85477c9e298a96465aa78dcd52a1b900ed734b355c14765a82db3cd77e80a609e32ff44faba03527e2e2440e0773807ee75605007ddb0c1f4b015ab3d04d52671d4c4fcd4b03a533ad18a5274e402f6a63588ad67586826deee1b0dad10698dda4966bbff02a4dd1cfc200cd366f66bf14b746b156049b9afe2e2588aea2d039b79bcb96f90c19e39147bb5fc7ef7573543e7453502d5d753d2baa6089426d1078571cb847aed814423a32b3a0ffe6a31508c8c60e40b1cb96be9a753b5945d18b455f7d80f8dbfef54d5cb1e0d52b270638bd1f77969ac52c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h5aee6a3862425f0ce59ada7b29fd9165e440ef05eabee973a0dd9a4676e18faf6f6ace64db8943b24eca2b14e2dcf9398d1bc83536973bcef02047860979e2b2c2ef15d34fa976f3b5d90cb12bae18fa5fdda595b1d5a0b20f6d6dad07a9df24fce7391506b6f9b0d431451db0d323d1ef1e486e956839ced8e1cc6fd0ce241504f4c684be66614ef344bd65fbf5af8aad12ac7b747e2c5ff3a987bca0e59ca8ff0c41bba79ab19e6f998bec349ea0b9790a60477f0c2191cbd56e4eff5aa103b19b99e31a0fd1809938558584498965c99f6f50864e1c4897b8b20b7834d544246c0bca01cb2bf7efb5337e2f82edfc89c4495b19db502947eee2950fecf524460966bb1546686edf23a9894bb04188a50d5d4b85b408d97e03e05936e8197080af91549e6e509b7e3ad5a73052f8be32fa910d010d56d849fdc59ad096b6f7ca7c5941ad42b8aa1d99a9224ef07b410d0c981820f67b6868e156922d5e20719e24e31bd5bebc4352caccb11ebcd51cc29e8d3d8758f20ca2be2170e1b4e5a15b9417008ae493c5bcc6b06015c0e83ee7f4c288a2760294bdeb5bacea0f9a20b85a5b526e110676697855fb4e91e33c73bb97b3748aa368c11c828c88331261e5521590eef28faff0d9bf675c93d27eddc936a9305f44717391500b33c7637121741a389305021d15a9c8c2949ccdb9cc67cbb7263b2d4483b3929d238af02aa8af86fd90b1eed95a8d35feca82106c5e3affaada7f7c6e4abe5aa54dcc66bdd8ae3a91f9ea6229d2e42c4193495f58c8c370f4a21557bd8480d2695db4ba7609854a64cfb2cec1fd4e7cc1287d2cf8dc413a62f3b6f15538addde01c1183baf0da2905bb95f72b5b81f444b2ed157ceeca4adba6a6f4d2f2f833640e4cbeb0a763d6a6481e1826fb481ee095b37e810c80d173c2e013e9d931ac80310027ee364a637d8d927634b1b80888573ae2e678e849632557c29d24efa3e74ed9e4a8803dfee3d9a9f0d4093c5f5acfa9c23bf426e9f8f8445e08daa57f7eb923485837e1e72760fa41a829c9b27d122517b5df18238a097c9031f77c5fd2ee57fcd22432c448ad270c17648a1a643af0d9df7b55373e7b9d1615341b6a781e24c0b649aeae72e7e54fcab2c7ec3b239daadd7f34a91d4bd8ce892c8c0c1a235bbd02ce0982df5e2ae5563af02d6f2453bbcec06cf0aa05b5cd61713244a744f83fce4bbcbfff3e52770ccdcaab20e1296a029e800c6c1ce14bf283855836b23799b1b0f69d57337f0dfa3d713565eea75349a4e5e6c989679bf28e824c01a5273569d9f8f28a41dce889af3a1dbbc8f2316df7f83ca87e78cedfd3fa74941a92153f20fdecd9a9da8abd885296cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h655b7d585a5943570aa3f57d0822e5536ea8e48efc883b3f4db75c7c99a4994a952232dace20378eae9ea668cee18f0af30161ec7196d0f8916f4af175ff04d6fd1a6cb27607a5bee97a086b91b6efb5093e6a63e05729b77a0cef46ff2cb5cf0d3bed8c2d9971aa6e79b02956307949ae4113065aae0ac456493c404de15eb250270da05761b8b1c7fe5fffb76fbec7642310f450e61990d947d2a47a698208c7dbd63b8b6285d42d7a36d3f1200d7f8f69cce2e1f5c0a8da0c7bba7cede6f20b7784c0ffbc0d4cac4c3feec3dd92d68bfae60c11e547831cf405a8b5fd6a5fdcba1c115ead2ea6718326e16ec6c6a243afb2e52576909b044efa53a082245df98c9951e2efb0864dab3ea5557db52331360591460459c860b27f5eea0859f1829af80b5597b05428b7d97522cca0be8af501c8a42d0fbe25ccd4511432d7e79c4960f2389bc984e8c908f3b341086d5202a06e5c434ccf8949e2378ffbffaedcbe41cfe3f732c41abd3356a95dbdfeee3bff82ad430bdb86f67815bebe8f5d3fbdfda0727b1b630639e11e8d587850a5351c7e90a9dff3b7ff820fe137ac3beffde8d6abee1a887cf60a7ab9027a36754475ec53f49869eaebdeb5a4ac15fcc300a1fab91ce049539ee3cc2d454b50fa5fc98c56af26062a00fcf486cd82e10b9229fd9dad536b67d062e82434f15e92d50f2e7a5c2ff37e685c3124282e542e899ce2c861edb77e52e0e4c092d033309825b1aeca6e6e1df0590b7b341e01ec2fa7ef43884dfe3c570f0e662a1f8a1779341127430ec6d5550a1f9dc23025c56deadbab37bfd1665d61737c15e3a3d553bc22d7604e2eedb82221c1a12f9d119dbde258b4ffc6429c92f2fb170beee73d6bc34c988a4c3c7f2c69ec80331ec77db7058bf5a495931f284f95477eeec1308e70e3f442c73accfeda0ac831038f67388d0c90e3e90ad65c99c506fa2893bcd428ebb0432802ef6719dd40aba6f05b623956655a2a5febd69dbf9cd06ddd502cd7054fd6ad4c17614a3ef37fa92ded9ea067606552f539bd466a31cd03790f07837ec7d435aeac05c1fa0d8078fbf02e283a07fd2882fc81f8e9da7be827f3ca6511aa0c00cb3c54c696a68cb8e1ef8c8ba027b096d05dcabd66ae2cbde825cb27d9be8e86add8a1f65e6d7947d8c70d730b95a3a6a45394080aa0dabed5e9ee010a691c3f681e8917b20a0a82104aba1b2affe3f05164e0190f656a92c611f7e9e35af1eb06d4198c2211b26321263034cf58e2cc4dde40ad1e1bfcdc6c432e7b9e836fa0e90fbee7f4c13f068e8d3cd262470d7f5c085aff913d04e60d024c41e421d2ed99176061d0080a17559178be3b1d4f42e6a33452;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h57b2475bc76df94d90b259d8038719dc3a742f49fac52bc5fa2afbc624b39cf1ed534e92248d64296c77ba5da5a57850e33bda6a34c3bf585de2529046fb5116eba6d02cd955d459e5e6507b3f53d10364aa5219b530a199053b864beb89a0ed5d4333b9155b853dbf8f3e353e6cbe249d29ef392c7083fb463d8ff148e9513780364e6b09f2bf02456e2c4460335ef580a741c250df69667b353e2c379d496e8975d304d8eedf8218b095801806304725d2490bbd5a459d8104adcab607739437f833c43b9807e26235d2d992dcdc230809f3a7eda46adfad2ab9ea76f65f67cb675bc01851b35cc1afbd871b6af58fd4befe6632625ab2c59c9061a8d59a75887e2d2814bdc136aaf416deff5ffc3eb2e0246252046db56de1d9611029df58855760b5ff26b6609e6e5e3512435ebee3c49305fa568068b938e9939f2156a52b2fe8e61cc80d1edf73abdf74b65ea242701e59be4f7d6d374626cfbdea8d6d782917dc4beed0d1492ecbd9df5bf1b5ac30ce4d4cd050151dc1e319f445acad7fa575d77591731bc559735c49fb29b3ccd2c76dc65a593c95bcce8e9c5ced200c34660fed5911bcf9ab260d08e82f13cc13d9b57f430e84a009244345c7c24e823952e915eff289bb352be6b05cfbf074734cb02487f0c9a309abb5572ba18cf1c224d867bece599a45145a726711ba989b5576e30b424286d4a5c2ddc941a305be99e11d55d560b54310ae7b4f5df7ec08e7a691d1d9c2833bf42aaf72226a71991808011f3184e094d0a8c0dd749145c26991458375c8cb7da252ca6aa0899350da3bb21ba967fc44f9748dc8c623ded08a8ce9bc87adf4df0c30c87d994090aeedd7663d839c5f0d1a0dc85613a78db5384cc511573f6de549d16a32d6cb0de6461ece6d6b93f54efdc7e8cd64ef251b982e11d70de220fa0b9e037c9f0e262bd946fb2d0b4929700f02c79e110eae3ccff0c43a3b8d6aef70df6e62774f39fba483e18695469e0bc97227b99db3c45ef0e0e3a3d4952381ebee941fe8c01b25c5bb8c8ac6610ebd6c57f12b27fcf3add22fdb6303c94d82b06cdb90258f85db1a0968e8e3f39f16c00bb79d921b9fe91e5249d8f8ea8109a2700be7c0356a5a8b0c454197070b44ef762c221fb5d487313d8e242f8ef68418c4ac11d882a230619ef36b5c9cc04ada4a586ada8592f50e4bc7c681fb7f318c0e57970d39280604a8059210c297c2d15547b735c860211a018495a60cf147d77678c82e309fccfb2105d7821deae5e4c60b76350e8a4b3ebeca2d95b28ceea8e9ed218037ace3ca75bd309ca8d2fc6c59006908d89a5192d9a1b4d25f6fe00c62f916b067e5fc6f4774ef2ddc3f6737;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h66671070fe61b4f99c747e90a26f88235abfe6390ae95147b32df4a067a90a0463ef743f187d10111b2c1efd80de8645e2d5035a869bdba9555c94c00b9a5b7161518ccf43da23b16a9de4d6911c99a1c2c7e9f053da72103ea8dd6cb328c82ed7106b4f5ba1edf3ea393ffb608206291eaddf17543f83bdaf88e5b6a4ea9b5495040d3761329ff860d771b6e252efcbe01a0a01688c1fdda90017abb90c56ff4b8953c3c3cd57cc0cce719d25726f32e1ef7454f21b77c862b6d1a784c1130e8ad760abdb7cb36f83bff534c961e38276834032d5b69570cfb959fc923f4a595c96a5b3ee8833bef3866e07574d37d9d4879e7c1374049c4c01807c5c4e26a5acd4f8a4bc22cda0a2e6d8b074d7205bbad0fac758e8da59f666cab7614a69ffffcac517a411b1907508056077d6d8b4d528a91cda2927468d1fb3730ac3b5c69f372c41831be53ef968fd5489867394680c08ae6de73282d4e89e3f81b8537e3ff4a47e00ad9be9b92df7ab890d6211b3b7e1f5ee41cd2ff86dcff7d59c5c2f38f662a9f1d1bdd4a9a7fc5b87556c5a07b2fdd4bae7dc45ff17e7e6e932814038b1b13c5773a2f6c4aac724753b4bdf41e5f0eaf19568d5169123138072a801ba5ae06eb1dd93cf4fbd14b2eb9bfbd304dbec8c0f30a05b72100049a431cb8b649cc9ce9fa2f61fe41d7f64093e709387bb059e7b17908161b49dcc73b95ea6a1a810e3029faa00f04a8bae3cc1e48a6151c897f9fe2c497ff24a0866e272256dbbccb1a7a457ea3a6a63091cfdd0eafa7852ac6b2b0b3ce9c53be76e99ba8f6ef1d5836db20c3e39876e56af477e9794567c5f563558e0bf11d3c87f7909b4b62461a3b6db7c7b315a697c563a602bb918f865d9d1f78793993fa3b8d09e6531b13bb5a20dc1a8f98af64bbdc8ecb4f60be443da7e4ab8380b02af3d5c46be41c594975014e7931457e570895c93f236e559e1ce6b5d2e77494212d072f47e582f24d07e3b180c35f12cc0c596d846e8cb42d23405db8d4cebe94df6b94020c0c29f34aa024d95b80c10640a63267edb0c8f1f0e4b57ef27bf79fcce05f2012986588c5b5a6e007ec90e0f28dafd94013cd4e99a5c5040cd219c8ea512865474ad9553417d3a265a96e32afd37bfbde8c2428c80cbb237ea43025d880617e586ccd3185b8e67d87e27ab89abd7596d3c7343509abead0220f58c7dd7a5c7089375693582dbabc2dc606892a8304987f0bbed4b660e029e0638f18ccf22f62e10cf4f25c694895a15e88bee801540a1eb4811713f62b48d4507930d96792ae374e864923e39983eccfd3650c1546718e9c66de9d6fb83231373cdadf38ab4bfe04c462b372f0ec29a4c397c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf306eab56ed8c2751b4e3813dec90e48f5a5f0930cef56c23f59f46d6bb2c3bffbb7e56130d7c1ac809a71c5cfc7f2a7abfff8e6399d771c3060cdbc3b00cad893aeaea68df98a16996a98dcc434528b563a9e6c73fdc8b6d89301f2956ac07ef20f933bd9f9f88c3eb9f74c7c49c0a957cb22a1cf90faeb5c588923c1100c0bb7c0132267281166a36f23ab0690b6276ecfaf683b6b511dee5aeab57341d8a22398ccdffa3f4a79a760428a643f6a5b515169d372fd78bddb91c836c100768b262c08bed51c51078ceecc6e8172b829b31f0f57d8258b1b2f7d8e75e3ed8622990bb9aac126f0bd4f2b09c79ac4bacb82280396c2d290ae9663e7837d6b72119d1f9c90b20bfa608ff44780ecc8a7cf809fe2b737741fcf37bafd151b9fc4c1d9fee8827dc952bd62c6ea65b9fc8f1fb6dde29c05149e5d6e1396e36f3eef8a188b8a3de4ff44b0271946a446877060e875c26801802fcd34a47a302d78a58bb02c5b323ee09371885dbec3705c424f8c4c219071f23034a2da54a4497ec8d52fb989198ae3e95454bce0c4af8ac918d8dd4c7bf4243f089237cbbcebe6e7f5fe9811df9b8b33f09e7e5f3afc647dd6886fd41398eff3c3a8382135c9072b3aaeb62b6058f4e6303b8191aaeaf9a00e19e5faf5abd4d95e3e61259b1d9bb9f5304b9f1f8da5a6412a8848d8eda5060517aa6cdbc5e78d96c60c278b764beb7132adb2f032a297d511a9c4fdc7cb3cc5b488753ab06664914e05afbf5fe42a155d1a9979de7592594616cf1699e4e17cd5f24de1e000682758bc5115b9a111d77b5f8975de5a6a4f93a0a4f1f05ae0b3e17b09c645134aff0f883e60421dfcf328a37f2e55b6963b2110f29285838c55f3c45102bd0b3526a7848cd360364fbe8ad6dac067f66e535e42824a86884ef5fc29e9e47909f01cd80406f61f7226d60f3adcfd3823b92e202511afb108b93889e84d27ca0a718f00553e4d604b12892ffaea07c26a10875d82ec778fe9f85bf42ca2c01ddedb1f2f2ba249a657f70dcf9c8ccacec9ff48ab048f28f66a5d5c333f73f2ce171945ebba9956c824078ee4172c2f2172e2095aadac693ea8f863e6a5b1f28b67735d197d99fb62616be39e2a580e16a83875ebcc5ca70d1c233b8732a5cb9c59515fafa08442e6a853b1d4d0fb20bc5f0fe035bec86414cb95baa45164da5721e61cb857187eb8e692ba13b5a70bf1942241e1d3442c6a522f54b9f921c7da7d67dad31401dbf8982940f7849a27ea674e93cc0d9ecd5383b8887cc9d2d0afa00661b8427416b4e4dc40fbba60c0fa75754c7256201ca89a16ae078e365aed15350cfeeef6ef81651085b4709f122fa3ca39c3f3497d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3c7f43bd02272823397478f7d2040eb534a8b48f74e66e94671c796ca1b3b4ecd83cf4e0a4ebe29283148be37267e874fdaeea58c2589fa168b6a94e4dcacddea465e82eb96e2dd7f1582c490403c7ad7e7411a8ee366006a1741d33c42dd15a245d55fdcdadd5c99a626965df90074f222e4ca6fa5cadce3e270580b0f0b93f09174124239ee833f52182f396f235c3654c9ef24509cc8da9cde49e77e8aa5feb4dbc07bd186388aaeb0bd48f9d6a60dc138f2352a90ff302aacd6e323ef6267a6b9b64d069ba607fa061e2d1a35eb67d34695ab11c59c4cc7a76f9412663863bf96882dbffbc36a1759f6b138711fab33802561c443416f889918af9369bd653215a327499a0ec6daead5db857565979b13ed1bcaf85d1bf72398d1c49f0feb3c4a59f6683ea51d8b79ad0684a654a8c4bb0d3de4e55b8591ba4f81aca3aa79eeb218ac2accd9b2f95d4fe6c5ca94e18e5b88b66306354237936bb4d3e19108afa780198ccd97bbbde7a0f3be7e87eae64f0e98e3a290081e7378e9b6b739cd9f8f7f042306f29d21c7545fe406fcca5cee9466acba0d6c76c00943024477f28592f02d39eb535c803b85ea9100ffd281df7abd0d105fb1086fea2e884351c1f92a6f93c87dc5124942550f794e60ecb0ca3e895ef4c770edaebc16ca9eb124738b1968c03388cd2baac4ccc0c4b0536bd7b0edd30eebaad8a08de377675ca941d5d1b2620c67a2a017685c45fa0862fb35c47bb45cc88a8f3303847a250bb927404653a23b5479b0b0d22eb5ac3226075c571d0fbf65fd1d505c424f90482056e9d7cac280f3d524454286334e7ef601935467708065023f9c0c5a3c733e122366ab85a83563f64b4d6801a79abe017baae9ce12257f3e76140f0743a07651b0fe2442a9425990f20d828ca69b1fa922112e322553fa225ab63c1f93bda013a522d4ad414b95fe5ca95775241c34ef8b0ec7f532eb87736aced4f39fa5bb1768d055ff95f8c0d82f0c8c6aee1321fe7c80ac602f2034cdd0c83c96ba4ddc7937e4c8a60dafe180f0ac2de0bcaec5c5bfc22704f788d845cad232f5cbcb4268a9c2c414caab6e4e10f1e127be98c052e2e54af02bb8ddcde5648a8b8bc6d457aed15eb4977b5d34b9d49ba15086784b3730b75d47270f1e4082df7a30c6d3f1ad881d539d11590b3074c31785887418eae3d8dcdb72a4f0218f1612460e7615bc7687c6db4e1f6fd8002aad53de348ae2724fc6af9cf2307888ebbe1154a469b9014b8c0f7bf1b59cc5e594821ec15ee5579e0f35fe99f8f4ea727197bbd3946a05b0b79c2aa417bb9ed73401cd5be7e94775c168fd429421c556f5618a7a7195955ad165682a2777cbd32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h655c870a9c469dc63d965e241dbc36407d078f4929b8449665dde8da6171e6d3118a6310b4749751699c1acce125c6faccf1a3aefc11310f4262ecbe399b1df74977aba8e72b9b7bbf3ba55f614dc200aa8ed65a5f4a3909e612b55cdcf544dacee8c556c956df62fa3b34473f4f12804e19a1171517465e06f3706b33bd09775dfcac801811c255da7bda42c28c8d2fa152d50e446cd2295d0e6a19724a331ff24fb46cf99c11285c884aff0667aadedd523fa9f55d8983bc531d2ae6e0e9b5a872e9eac52e7f86b6db71e7a30a2ae1b6cb67ef5296fe3a5fd5682163f2eb2ad5f12beb43c891778e319c852014e628170cfff0b857304a5195cd68c1198a7d2ccf0d51554f09c05e6b3a4d5a8369e44ecdad1d3d6769d37a773bb1727b98ab85e6f611c4f76e911af90a276ef32a336047bcb87195bd43743bf2675d0197c76bb2c2fce3fecb4191c8090a37786175486053fa03213dd66469cc3007ef481532daad6d780c828bbdae09c5d52b6068a4683202fb9901a38fb69d8c1dbe2fa278f0ee08050781372b608455de892be59dca8ee4790779a4e066e6bf98880a2dbe0cf9da9f5cf84474434136c0ce8a7a01071d778c5a8e5c440c27acf665d047eaee5ac90a64596a826c7ccb35e6fda6f27f74aa7b965216013618a52dd94a0842a53bbd7b0af69afe167e2a26328a00e7a47a5cea79b354e20785fa2b7f5bd69968ac6d095d9e3b09510b4002bf17f8af0f1ef30d952992dcca508ed2c41837a6db7a93da0979b39fa03923533e3b3eaedf7c56d6bcbdaebe9fdb0782bbdaaa0a7e6189db295532466e204a3bcc72a70b14b8a4d3c4f84f7928aea11c157c284228bd7381a7ff92b29af0a1b385cce802aacafbaee94e45696dfa1a899ac474816889d59fc29b5696c34ec721aae28655c4217f16069f35e081ab8184ff4542f1c375dd0e2735329e91e6ff6869107abc999174956dd34b8c784a1d609e6e714e595ac32453fd925efde0435529aa1752577f6663495c8726c2c9a0814d06926a72232abec15672cd2761d6fd302c3acae07b4d300a3d9edca26493a2ede2273f09baad3a0f024c792327cd9e394571bd5a74dbbd459ef0538849362da291c1dc94cb2768afa6b648a9f220d1b1cff944286728566dfdaf4e15c460d0ab221bb222173567e9bb3a893f738814bab8a76da9a613177c7187a9b269170fd249dbe4609f9c8cfd06223d8c3e1179d72c759a55b42e7c8929ad322110232d3d55d6edf14a91f3b6b1816afce5078bfa2286d3cca364a3329e2c6d4588e78c00ef5a892edecd2b942cb08e841e8d9a8e106dc25fd068b007c8999d1fc2248f0949100bb04efd695dd54eb7f173d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hff85a2f67c58643db96ff3445cea5e2a66f871b4d1111c5d7f183ef220f141613d7b3125d07de5a1df2de67c7427a654bba173b48aa0a11e3ef2b4ddae847c223952ec47575d429976fa02e6d6489f0ca2e792a9abab66928f48c37ebe7f2aa6d5befe1557d48104f2a609328706349a86a693e33e2ee9a5166efdcb26d29d4e68781f21b7a3f072bcd80a63acfa03a4b5206974342d795229425fd546da01558366fd50ec917cb69982d3b33f3d6dbb4954ca15bf671c9b38da30d50ab2dcf7b416028a6e5374481b126d4b6843d34225353f5ffa520d0079b686f27e59f9cec8bbf92e6f7aadd2d68fecc2d70c1a3fcc4999a30649bab4e571c2f84260a531c6ee9883290a181c0d44ffdbac1aafb99570f2d5fe4d7b133d814b0035fc659162c661d0e0e51ddf4c84b31f6881fc185dd0157be80f13eac0d13f3336c0f58ee9901e6a5e9fafc3945c954096d966049feb47343141480405991d2b518502a1e72ef176cd2be80c526fc524734d3cdf16c4ee701a683e495e1dd94c38019e1398d0d789350f2d8bc1a3b58ec709a034b1626e6f0c83bfb79631459ed3d86e611c4ceae4fd95beca42daa2657c8ea5f2447dea9f5444738e8cb4c63bbd37c78fe6fe12458f4672f5cb782de27e04ab616e2d93bce49278f3095ed6ae5a30ab809dd799d91f0a82282b9a12429b8f4bd0c71341db0b777a24d813b0d304f4840492b131f52a4ed7d5c0511ed6f8247c5d6a2e48f15f7069b458a40d839859325119cc8416f5bd13a186f4bd544eeb57a5af54396414f133dfc281b97c6a470f5f112e13b8294873c270f6a49b2fc71bc8d22d40a326be2df1f4fa2383cf4594901ae0b0e9cfa779b90c90e7a07c1e6accf3d397069f70c1b97ea042c82371502b395f771b91dc5559cf2aa6a1c81debcad1650c9c3e2d749ea7dcbe8ef1fecdbe49e2c09e017b69ac4d805c55e49452d2201ac817a096a2f18786d23e0ee352833dcf4281652f6c2f4b2f4927843c6199d6f9af5d58ea3e853e4710f665eb07621685f5d3b0707da3638668c7e375c16d074e358a993b62e1be859904600ac22d81289564848b628b8a55bdc6a2b30277dca0d0c8307464e0058eb284875ab453c46960f056aff329ae2897d5c999dd640026cd9f57674d551a468405b6513c20ef505b4bf34cfdef17961eb69028b77a5219432d6d16b69c16516a2ebe1f37716f63298909dac6a4e190219fa65dedeab00954a9d76334176415a2831736a5bcf7f1ab058986c59f437f03fb5c0f0b34f5566a02ec2abf7b20ddacd7184dbaaa8c18bca9dfcdcfb79da86fe6f3af3c07bea64c8d39f3355937a64fe10cdebc33a339b891b600ffa8c3817af7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h360d68e80eaca415aaabf2f5b689a651457094e6ac95fde09661c099a655fb25100e9d24ddc39ecdafa827b31739869971ef1395e9baa6ae07eaea8079dc7c50f784761152005662adca362df1c1aeac679f55fa3a0337e2cb87208e0886e37578c820e6938c0f9f68d86912cb1cfe426079ef3531959ff75734f6217eba255f2e7ed362370002458aaae2797c41416cfb760973855a85a6d0be52161ca9668e19e52deb210ac79bdf3478ff2dddb8128ba59d5c9b737daf878f50a7fd2476581bcbc4610c29a227a53eedfddabebf753c2773a8ad6716dfad0af79ca4ef19a3bc342ae9c50c9af450ea1146202ff5133354c21e274abd1436527b0ffe315a853676439bbeb1abeb3f1c6e5c243e92051713a1559d7122dfdb53fc5ab7a507c4ec0faf4ad59a7bb1de9660c9fbe11eba1f44e3e05aab1ee7f5747d1eb2fb5f2e79d57242bcc7f44b1769e04a32c6b402f1e6f48fe089ff7fd960e85fce6424251acb10195f905a7a4c02fc19fa63583388670d5429e4d3349399bb36552ebe1750294bd021c473bc32d747f2c08202a875f0a160d2866c99995161058069636fd367a3f0b1f0e689e23cb54cf342bff359712c2ea28e98fa448195269ac7fbafa19b7d26831811a08d52a6437a5da3e4c04a4fa415253fc914e3e132034fa99b00e56cd1a9e8149d995948eb2dee4d9076773453f32a4a112a420cc92345c00878a71cfdf74ce93a2538e02615148c07b7a1882959feddf4f19b732938d8a071e89097bd66d67906dc188f00351bb0a6358f4a1186875d0761aaf0b0a652e917945095d2bf88e462de0e80abc9a4e29dd34eb15cd69d91b74f977a6a468f1677037324d17a3e693936ffda9dac22a003e2f1dcfebdb482a3e6abd4f4199c65774471843dcc66ef68dcb634bc10a512f52dad7375b25323cb00c3f14a25ba548198c5ba741f4a82cf3ed43da68cce78633a496d54d6250586516e5c5bc59a3a9d38c9fbe3dca2d37a58558ec60c0fa900f1306777b7e4080b6ff8c553a09fa129e745a3bc1dd8997962946882c64f5f300cf986ca43748a9d03696ddfa12a50d82ef937e9457c7a3dd211488c731f3410ab745aa44773aba0b1be2b74ff0c36d8db5e0f05af81ea2a259e7c1f360f7ed73886d9fb9cfb1220af87cc95c6740210a8a81862946add6e224d8f089db2d158f861b9b10a1ee7a49ef8ae6391f7927c2efec0a6fb64f8e56731e320962e311c98cca3ef1ac52ba0f690d0904c13baeada56c75dd639a00d962811302d8b8c83bb4049bcb0a93fad1dac467420de137cfed5cf897f0d9e82c805e7a8767fadf38bbe2a10df8f230fed3d21f9ee161f412c02f2b005d8749a12002612;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h8d62b257c50bd3da9ceff2e401fb9dd4d5e227afdc5eb2ffbf3541ae6193d73594ec81b727ce292366f012ab08c100ad6932acf0b25913ae7d647787f68a5483268558d3f3398784a52e0c69221e5a5261293b7daa2d7a66887896a6f1abbb77f4185e703c1e0e2100600c43b17adc19618729fb3356e8f136611a666ecd4a384668798bfdb4dcc2155128990b48fcc4f68c1a5fc7331079780c8b078f219b7f0808c88ef87526f75197064de18fed2915a71bcd2a6da07ea5f8c5cb6944384da103a488da2288792bb4aa60cd58a81e01d0e860b10abc16e239b8b220ff43bcf3e21a71168f5e08e4b265f99f0f8440b113df742546112a7151fef0d5930d6d108ba4b9eb07361cf25745fd0481d84f8e2a3e60837af11725621adc6e48ba4fa57110b82b1b2691399257db490a664b8893752cf55a840afb1a90d2710d7fa0e5cab345e8d1796b4587b8d025b26abf2cafabfd9be4fa8513105cafd300bf9a3766183a8651fc323122636b88ff92cb1dbae0cb40314753951dc09a9cdcd412aca1fb8bb601d9257b7a98192682799a9c24d799dd9abfe43413ae76435fb1e18f2fa32dfa92bd6053a1c122e6e84cdb2a851b4cca8c1a7126d333f29952db2eebe9f041cefda6b6d59b3a4386934a66df76d3acddc39548cd57066e75bf5eb2c98f658e2bf02d25752fda5441fccc4c0ebf077c214c3f756609b686e2fbf2f411a1b39706ebd7f0d9decedca59b1081e91cfb03c1df100cd5986532de207d9ba837ceedc1891c62b2ad2ddc022b0592124b883f1a4a2766a45a1893a1e622d2901151c7551debe7fd50864430dc8037b7d71f76e9e09cf51e8428614be3c843c548390f7239e6c66b01b748f0bf157d0dfd0e4da3ecdedb06d73fe3847cf5ab32b8acf920ce60a5d96c6268df1287bb027964f72beaa5f7d5cac643538e2dffd7c6bea71cad015ef6d11d006e41d5d295cc1b7e1993ea5e0233472ab24b38d78a16cae14aafd07d952352e92753dda2ca5642a0a7e664dfabd2ce83c1c01d348bc90ba5b61754c0eba156c1eaf111a6bc01047bf959570704babbef48ae58871171e77061c5c16dbaf1fa60c4eac1e828fe695831b249bd5c88e0abb869428cd0a10311bcc55b30d2abaf1b562a2b689688a1c57fed65ffd2119f2e7b80548a4ec2713e9a201f3d4380b3825aae4836091dc54374f5943bfb853da983cef3a54517bc17587935884db7234af82079ee3fa4dc5f8bb220141886975dd9a1330d02579caf765c333dafe8868438ea2c9ff5da182b48e72e361c031260bcfd9b18b94d5482f09dc597d188bbde69820b24ebb773de9a36285ac96e2352387a389147a8f89c1f06b917c62d78e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h4c867c7ceddb3a7b3f303305f90b6b0f865573253bc2d06d9f05f20516271a8673eb5b474ae66e75e28b820b3662e7483bc6993f2f14d12a0f70bef934447c0154d5f6f82a020d79bf8d9ee8985f6064fd53ff5f4d865265aafeb7dab23a88005c27022c5a7e88defa4cbcf3fa7d4662f82d681397b62d979b3edf75e0f4290743237745a2b0359fc54a90bbb18a8148583250ab4ebded3ad30448b8f7d36b2f0a17faab928af769a62d2b7bc35df656f3efced23256a04ce2ac0b3e03dd29699c5c92a7a282a0211877bd770166a213b6b254896fd630e92ea311d7920737ad72455d3125f4558ff4279b33d9d554570f0435c5434fa760ba1df48d4374617a9ebcf1ea0d3e0a811a9adcae0d8e02d8e4f35c1f621d9ef569fa5139adc8d4738edfc83c11cb684aff99e86e8409493f5b65735a900a49f3ad1ddb127a3e9c981ca54f64cdde53bef4f3c6213bba98f8e59bdf77c58737fb6f7600c8bdeb62645b3bd9f4fbfe6f27681eb5bdb6431eedac628a6f4338ed2e1e6b6773ed16acf2add3dd3b705bd6664a9dc2f925e937434b6a590104457b2ebbf02a6e6640c0610c64339cff678f15ddecf83c1381b3bbcc14afc3886bda8307adbda21ea73b9bc6498ec72f45f52feb5a34515c6a031de6a48ccbf6d8e8759bfc37e32bd19bea9a29e69ee4bc92f797ddd85336aaf15d174f6861fd61774d9773c1b6307e987f6caf1a3f89a16b9d48a19659c21e5a1cb16d62331eba1cfc0d9d3ca8edbdab8f28bdfbb952d3d00cfcf960e782233a2895982d24c01f45ea7170b8b12f80d04dd2cc4cc740e3d59042daa884159237dafd790a223107e905475bd74834cbe3367bfff41eed7d986c1d612f6844fbf9eb0ebf467fb1ed90164bf85f954b9eb8f2b56f179d7827089353cac058251aebb9ec1f0b4b686b86228bbe493077e3b8cfdedd82c981b85f96654d88f81743429c0c302dd356153e34ca52e21eb52d67108d1e2fbfa3bd5eb0348972fc9e99621bcbdb3edfc2597bd2724f547c8218a10100a16cdc9548f05cff638ccbc52b011f499801ec1ff67762e80667063583dc0ea1ee6ca750b570fbfd59be27006fec30e6548b3dfa4c187a2a4904fbb77dda64999665fd84fe3bc7f7518c3e997bf19f1f5ef92a3a7bfe885e8812554f8da80809c8a4d333a6b4cba18704285c5d14236ed3379cf1f5fccef05501fead4b1fb3f330790baf5f9d5751a9d94eb08a74103abe9b42badd50705c202c3f22458470c84f0f496997fff9ce80b755ba96aa0b68a3c01124da950f2362876de9168313375e307d6548842ee21034bfc302378b3294bb6fa6d59b20149ba0a380b748ac45ded57a298f14f9ed7930f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h1428f38a224077aec40f7e83ccd174830e4b6d6b1bf9682af25c7d5ad731c7c66345bdc136ed8cf48b214c9e26010b6035a6835a42382bec52e9ce9dc25bee8b357cfe877db25053a45c8be8c29cbc4c3d17165766704e8b327aac7e1f79de03f6170f2995225ab3e56add67f289ecdca2c8fe18cbb89a135a4893da32d332ca1b46d516700475d6ac50e39214136938ae0d866131e59bb21b5692ade97a0a5fcb79fc5c1c2d6522ed5197ed84d25315a7087a2c2b612ba375cdf46b1e118353fe7c966109ec74d61093098cd29be525564761e3492e1f957da0dcaa65e638ea54a126603fd40777e4a0c6d448e331232b2770a5a28c03f8911ab979153708195747c1c4e1e7fe64f851898e91c854d66022495c608406380b3b85d638a1ba27d05f807ba454fdc1bca73b00160ed9a245ecd5369a0732fd516097d299733a18cf626cb029f816413fb8638bd0905c3ec93728269e57b198020579bd9974c118e2d941acd8eb07c7e81429e51611829f828a3137af5d77ee84ff02acbd601772c124e7851d333c952ac5982afc21e850f9c926cc70e56c94c6038cf23423f0cd3d6a30eab5d8bf8a1f2385130bd748467be04eca1f028be1858b230adb005bd9532c4532e7ba81c85082cfb1d04e4bf3e5477b7a219db495b6dd2797d25440ef868b0334c33b1109d02dd4dff3e0d36d7084323c318633444617b8d119f9abde287345d9c2f244e9843be1fc3b59fb9c0752733924ac6dd64ae9e940516b94f4a3a7eebfc0e460d277002aa63309b35485f08b8115b07e889d325316f88d7194698b3dc6aa62173758877185415b2c26f348a0557d8085141c6557cb04b26ffb9ed852be2220e67f35c7988b4c71b3b8f46ca37d09e24728ad06eee5153e711d46e66657659e168f425267b439e4f45575dd9883c30dc67ca45570ac8b59b615ba54d5bc3fae0dfa0de7edd138a1a70fd296337ee84e21d5f1d122a6328992d93ff4354e530f91bb5e60d6b7772c998966a00f0e6d88ebb263d0601a4d128a1dd12b9fbf2e3a0f4e3e0c8a05e87fbaa0c929fb2d4aec57ce059efafcb712b9c20cc0b1e06701f4d026a3d119a8e93a69d8e88139461f0d4a3c7d82214d6c3f6ac240cf851e48d634b39a4eeea1c8934b862ef9a32eeec4a859891d562835db286a5d6b1ecd6b1bb7118ad3614d08fbc25e2e79b1b47c6e3ef33b59c241d2874bfe32a7233399f04caa0de3126f82dea9195b1bc69b7686cceea63321ac1012bd44a886608d012cf480b572ab8779f26723c43fcd7cea9ee60c93bf3f5ae8dd13e4e0960434eaaf41521f78f2aa097e4d1b94a69098d8c2b41e8a55dbde055824f71e1452ffdb4673b43b35dc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h452601eac61bb290f5e5bafb3317d053106a1822252149876acca9e512d65cf0fdaebec7779fcda8b682f1acc38a5b0df956bd400153e129d57d4eb17ba079837cc085a16879bfb06fd807f737c9e038ecd1ba2e63638244ba6ec87bb243511aec13834e342d379f178b45f906f2b39ee501dea23141230ec4ff158ae669af3dda9baea71e56e55d79b552fe54f06889301a76b42ce7fa4fea6b7588dc7a147331ca5f483dcb3676c5c33bd083f013e8abce6f797a897514d6ab80eb67f1b876bc1644cf234ed23175362a152366b32c7d16516dabf74d8ff5a6a4ab01982f457ba8b627acdd61d85635b56ce8fe4ae21c6d3eb4fedac2ae74d8b3d5468250102532034b126fb34dc81708199c52985fff0aa85eaef3d0703eed7a481f149eb1954ffae017f20a7d66a87354f4434aae93344c15b5a956d8ea3ba92f95db8b3c50a9e61974da18953683e0182c911d7f753667bfe7a0f844a0d9ebe67bd77744f719dc1fb2c71206358677b246618c112f5d48757a4971142758978fde2a2bd6ba5f63f2ee13fdacafa7611066cd3c4bad9c978884429a78148055394f43fd94941c91279c51b4c101d2b2a8eeaf07355150240150b1abb7c164328a957ccc28bc3d3a7d233d0386137b2428361ebe691e48fa6ef068b964e6994bf72f5216f4bf9173b2e1b16ba7e6f48977866ba1748c44f6b57237d35df4082e91be8c11c419304828a72d7ad1e1dc7d77f870fe464bfdfd13a2c522270450c9b954a6d805751c415d505802bbcc95be5e5426bd9aa807ab24cf6986a0c1f1b68b3c9600a0c89fa53f8f6411100fc22706a4c23cc55002f0f5e2ab206582e54cd1d3ff53c5f85c4862a1b3d245156fe1387a141cca49bf3276b1c1ac713b237487d75e7ead3baca6db992bddff7b46e67e39e65aa66459429a26abd0926f6a45ca0071a0349ad95211efc9082c1159bcb897627a3c7c6e6b76c14cb1b97da7fde3eba6b92818c5363704d18fe0e70863a1cc5527eb4ff28bb774236ab83acfb73896e9962ca2276a2a2f77157618107ae96a56e57f74cc41ae4d29fa13a3b3622de5f4ddb16e2ed88bc6f21b72625ba796cd064befc469d0d6233869c43995eb9c47cc306e157bbb872f4b7e529cce45db154c54939931ab26bbaf756c8e7ee6a6f2a31cf36f8a2bfbf537cffb287f110fefee376c64cee023f84888fcb9d0bbbbc0605106726946bbf77c7de9623aa539a7c4019b2350cccea59aa363bb5baa02942f17cc6b60efcb12bfe60ef6c0d02a8d384481ae97c65815ff20b017a903a5aedb9ac355b7fa822b5b06447392e256c84801aaaf1a75f7e71202e3e1d4eed8ba5fb80ce8fea85c0c342873f39a8161;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hcebbd5cdc039512336241e7724a2eef0b5d7124c5de64f1dd8f8a736274a0da73cef3e55f2820b58f567695a24bb7e934e247d557945bcb766ee97268985328b4f4892e56010895f9e788e7725d0a1f69cb263dcbe4878f79968723f1a1442531cfb1ecbc66084ef0f1b15869b91ea9d8313ab76adfe4de1c7aceb53622228fe3f87433f9289d0267167aff803a15a0778d0995764fdd15bfda9714b5d3d054df51697d7de24505265da2ee121a2d2ec18270a34504462b6cd9288549db979bfcbc18cca148a64fc8e02e5079be365239159933a527cb8aaff2bdc75032207f52b54e99dc3e81d0b1d2b6524297fed95ece35e15bd6d5dbfb1a8c659fb1fba4683970ac3d34b0dde747f4199aadd81f82ca717788db9f8e2b1d2ea0913ed1c09b7648c899b3b8c7c5047e1ca3fa66c018288f8a2ef5b78e0501b2965ef6b63735f5c9e8456eee4323c12d9abde5fb0a75c2e59c00f161dbf282ce77e169cec8ea03e14c5c708bae1c88d553839df366d6e0a17a701e26ee239fec575fe06febc05aa2cbccc04c5afdfb196ece2f1589c808b97284adc948faba9527786ce504e5845a714d3477d7c9d49983eafb12123b52d1bba2fec761dc4b10b35ae2926c85f82f316446222fd8b7c2925157f04541858d3bbb11b580d3030d752b4f26c5f64837cafb216d24d605fe8d2b3f9f4c343e499cf12fcd75fb34bc4d764df4e19df3a8d8342dded14a9b3385b7118b84b04145762135ea3f4b9da16a963a08b4461d52000e961a9d4d85ea7269cb66eda3b60f35f4a2d91409203749a1cd3339106f063d74b434fb795fd5231c60e5f198bc4d5fb7abf56a0e0b53a24d95b64913adf663f862dd80adfb38419c28fa7e060b2f010d2dc5e8a11847d6076bf17ec9387f585791377e44cfd8f12703f92a096341892ad8e8a9b039d001b59e2f2676cbce24fa91d6aef4c27c30375f3e3b6c00048514f090176284b14b046e7f343ba695496ae4d3eb4f47df9e874985196b69f898216489f6d9096d6175d4c591fcb7aef70219233029b1f75ce461d92c1fe38cc2492ef6b7462a6e10bfa70b91c0d7c6b7d8ac13adefa2e3f3881ce1e0314280ab4d4950f212e7e4b541d1c1f7653b7016ef6e5224f219626513cca4cb9060e1195b4b3d35804be3e43d06605fd81584196d5437cdf4ae1c7fc71bb90dc13b14f497cf8f0e4f8200424269503d06f2fefffa23bb63a18fd0cc8a37bd0b1fa79d3e2787bf49fec5c319072d1765a17a5af57b8e3ff81ca820d596851beda55f247c2dcc3c70df2cbbf60154797e870789c9e742efa9bc87cfd4e255f4a5db65d41cc713bac4229f5b0bf1a65a3a2836fe12791c7b544a8703e4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hc59878a9e53b16d9c700d979c966155485535fd8ae9c5ebf1bee14ef177362daa2d33cea5130316e83b7c474afa765d12f8590a21f6064cdb3d7cb61a10d22f2f0fdcec3462ea164416707cccb381a1ed2c0c0f6e4bd17bde5816212ed4bb09ea2d02933322eb6156e353fb82bf26e81eceb27887828f0d930b2bc27b695ba4299508f579c2a185e1a2f8f62f816f61f9f84ee1bc61af857d24db13005ab197fe8e865e5362644c55bd961a4f7d523c9241094267da6dc3c919aa1084a9ff8fb689227413183a74ad85db9c7989ac74a5e8d8df94072b9095e5fbac50b8c6b4a288fa0b9926a035af0269a392aca31c9ba3869a8388df3bf3f6d288543a4a7e88bbe908a43a77bd649aaa10e5826fb86ce89fe49d1eecd8d6ad106a191f257fdd93b2972b9cc85d98651292db052a7fbb27acbaa62786aaaaf2712470ef30944fa51df8d547e2a34c13e2f55c39ec90b3aa1f6354871998936b191fc3f064f3d16e81e093983f7a87508fb9418467418b39ee4146c4437eaa475d74f8d49ef2ea955c23be652b6e934ae7ad46f9c3d77e3322cb8c777b66a9d018b1ba6b5b1883e5430b20a3081539e031946ed98e1469bc33a5f8f21def4607035a1aa6635393134e98aacb25623ba7542cc82454be0c2bbce6074c1576fd8cb56703a0cef34055f71850faa3ffdcdb9ac5afce9815c9ea443c7f463f606e57bbb20ad5d8ba854e28d196d44fc8bd0e37e146d9b15c76c3390d123e7d9c93768a2246943c7333ad7081857bf0cca09df924144974e84d376b890c7c99d47a24d493fccf95e3166ae5c58b0253ef23ad66c0cf41d90533c0cb0decc4f5d487ce479c8ac0f2460d33df557c488c91f223b28dfb544c4f161c7050f5ade64e957fcced5c8bfe500fe6f43efe1876972d1af9245f05bdf15f6149e107f85224783ef9524e02a165656638a2963796ac7f7da5af34f3d5468c566f8cca7a5e1884ed07d7f40d40df24f6540b696f9830a008a12b06d0abe9962b0bb8c834e78f4b4829f8cb7920dc4f6fede1573235089d4e3792dacc807b0c6b9c68da3590181de9d66f4d3c8deec9c089379457d55fbaa77651efbe5c4989c477d4af4c44f2cc80b302222409fd17dee961e2303e953e8ed07c7a02d39d803a65c02aa8bdd3c8146aee42ca854754f9665bae4421c24a254065811ed4c4a0c7c261a472de2c469286f2fcf48749b5444d726069a5e9e490f23bf4ee3142355e3a73124d05f57ff0f33443f95f45fa26b80538e2dc75552fab5ec906bad28ffad78233612d30f5f977660624bc09bc7725f07f88890ec3da16d0d7d95b610a6c325cd99ac44208c92e172cda9be3e91c5d7b72ae56210448671a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'ha3c40a95412592ad143f690a25ff45d677fb4d69062cb86a379b69d7547c0dbcce417b65b237984f2ba9d895766c30396d1374ef5e5c0a8a357d870f91b8b34a56914d37dca17b0f0a07a761e546b96ff4676f4132ad611366ab5956926549d26fedb5816a1a044861bd8740c6dd59dbcec7addc9c8d27e01ac9acb52bb9b0d02195df84a061184ec1fd6f5b584d27119943419e7c6c5df2d9354e508c12bda9efc618eb3f7917c92597d5bf1c132b796984b83448a238b3b43b0bce705fc539728840b74b9663313b7aac3d9b7a309b4717525b54f20b5f49e02d1cbdca3055c8b2cf7a20c4bcd6b0dc638512a2f01e3bc25eb1873f161277883c022c268320007ca05b6a1dacc1a118a9cba8e6e20cb9867c69a47b140330392a6451c2fea020e08d85e03fdfacc30f1cb85f8e9a541c9c1d06e4c656e082829b231e1ea7918f10947a59c6c18472d98aecbb3193331e7f148558a7337764911649e9c3f31046e2b24cbbed50cecbee150ef21a584c52359408f66c03203b4a787fe96b3423c4315bdc07db146b972d3f6b3b1f557cd76fefd9e5688ac7d4d4dc0de8693590e48fd33a9daac3b06d55da747e33cce43dad9c15414f627e492a015ff3d4781e166b5805ec9b370e5856f08186018b94fda2a023dd7100d499f808577db6c2980c8caa865f4c3c2630cead2275d1e51860bd000550eae567939e7567f441341146e8ff165cd265d3b45717894df92b10897501dc0f49d1854e09f54c5beca0d7f4f82684330d4fecd3e531e4aa052d67aa85b329670be994b4ae0a4f6cfea514c5e94637d4837538481dd5bff2374a3119140823a81b03a355659db2dede3d31139c1f6ed2fc36c95c68d94754cc3b293453912dd6f20a54aadf29da66cc101798193a0b85c922bc1315854c93decf89c31f75e07619a2a9205b64a681f9dca85c3f8a7276478503b9af38c9150294fdc101807e4818f387eb7e5a522b94c388d2da4aa75ef2f554d4a92dd9df2413751ff1e6394c83d8bcd806c52c29e540779792b4261ceec0090d09dee7e1af61f2fd8672f444e9c0cbfe8371398269390dc455046b01727cc7e8932361b514a95989a55076823f998276b04752ec3ee6fe391aaba7e9477672e3727c20e8c9b7a3b2cdd4f128e87f7f372ed26cc5744b87129800e8d8d13bee5c9b0f381a775144ce1237b4878d07953f1c4c0aebf9a86f74871fe0926c7e14cf49fd213125d6768e1bd9871edaa1893e4535d69cd11e6de0d2f59bfbab1f22f4b987fb06a9ba30c703b0102ea6abc7fcce7e1bf4c2ea83689dd3f3827016f6d926a63b0b34ef8db1b507f0047a30c8356c9617c381e3964e80aa70dcb761073cedd8c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h18ed21e4d44b67411a152013796c838a74bec3a1c36c37ca0e369da0d257391b96c5ab5ba19038a0c5b96f159199cc419fc1772577716fa1a6afa06f5e3448b14b9c779439391dedea7927ee7e55ac7478600b4bec534522c54f272b6bfda1a95d669dcdb74caa6664b36f6016847e11c1ab77f1d6d633c5765c17153af2a47ff31e5ed229deb466c77aa450e5cc2defdcbbb13eab6a42759eda291d41788ff46727083e6d0d19d3d3c06f46ea3d3bfd4f2cc36027944593b03b1c98bceb108507fa964d45ae5540ae1dbee2bf76942c960d391bbe3f5beb79a2d664070e57626d524231ab13df41c06006cb7790a328f68e235debe21879f2ed125c9fce108f8c15dd772bfb43844fe4dcedb861b681b2c565fc82cf9b7675505bb474b268c0e7cff26ed112d4379237cd10ff04e51ca5454f0bda935862bd1b95359f7a3b7b2a6e39fdaf40ad0fffed7e4af0b48082848473e676d9a1f2446f953be0f0f490f598929611b1c81327cff12f6b36096a7e235f4aeaa8eda50900c671ce5ae9acbef1d0b0edbe17b98f8b007a356bd904154e8776c48ea225b18b9e9b6af562e06bf04489bfc58dad05fe5a88398310953520542b8c0955b2a8ecc54fd844304d75d44337e7a105d0a21d9cec1ab926c9fe81d9611b5fdf09ea342701043ed95d21665a3faa75d65216296b3474250315e5ce71f9520bf0eef7f737fb0fa4966c1e10de42590450a9afecddcba7306cd72098d4252808e24ca89a1225c29a39646635b22eb4976ee6abe6e689c1d483389081361d962747e46edcaea95295a96488784f70927e95049b80e4fc949bd5dfff0901c5a8c209c1cd9af96e32770db392e49399b2c31a5588fc01d7bace8a3371dd32680126964c434f1bf0089292d13e5df8118d4cf3d830d68a2754c9555625b0f9905a94a6ae7853ea366a12e6bd4b9a792b8cc93d5c64b061799674d4a19b433a31e6da6daf4c41d9685aeeac073eee960f634c2f7b1e83375a5075227bf22a878d8e30223f512a76617065f5b6eff3208cef2a5b54088b4af9744d0608b45f8418f55ff77449f949abe167a0c604a51f6e125761984335e4176b7b90ab2b96707a141221fd523e2167af1d76f101b7fc400fe719b7c54603a66fdd87284b2b23c4dcf2388ed0923ea57c10976d99d1feb4f1e0c02a79c28fec9bfd672c5614e9330b89c801f633338a1fe48ce09be782c82c2b1e6c6596e39d4079851dc845a9a0aeb7629baa813c0fe72d440574388ae6b08b46b93a5f61e6bb314a2b71161149d759f69292f9a9bdc8d8de610df3a642a6d56c82ff58eb8e646595fd7d3371b187c7ea372ad10ac63f7f09e9a4ef84a17bd9c1960fe5a6b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h75215d873c7e224b2bb32684e073388735a78bcd014ea2a847057112f2a0f5176f67dc20d1845405238df2ffe77b33bc1385782c6e35895832f0909f4192d8b8c48ba484dea6f30b83fa98f167d6e3b99d0cc9513760472012ef12530156fb3a2b0a0a653172ccfe4997afc01a83b540bcfdd068da58f1525001f0d71e54c18d4b2f8b670aac0726a2ca4e5bfd9c1fa3a3c0a6abb3a4cdc573fb4f55b3128f94453f8c0e2f8299a6de5d9129b4884d05dbd6f3af8d3f9a1989420491d55bb872c8a6ef84e307b5e58ddeedf51db7cdc4cc8e26bdf6193e4c62daf220f0c195c75e79c5f2a48dd0e72331ef115bbad1214084759437e44ed03960c128365df5866c054697b5f55cbbe866f6bfcd50db799a910fe140dc4105edd77793fdfd386630b69bce67a6a903bf07657d18686323751b1af86ae97b407b77b9f22b7161d58be44ce37aadc8eb377ba3a62d588166a8d33622ca5f9b469494266c18b2450a0739d7a57b7669d72ff638bdc848b63742a050285f5ab20103d5e4a0c8bc1d83e886f7a723fc2e7e70fb4664d7adee514d7e8b962bdf5740c470b9b43d4584682265437de5601a2cf1bc8c1b4c5c892dab8e0b10c03e3acdf4de79e1c016e645678bd62dc6c8318c4e46363ab66d002ac94d831e77df11c4656d8823ec44b4416270381d640d6849e70d10a6798d4db81b462c9d953ab497ddf28709365d06e6ce63d0d6452f9bc09898d93111c945cb8186fce75176fce9d9f8676aaac5d34544ac23eec721eeaa9a860457f17dcf7922ea8a42e8ba22001067bce79f55d865ece37f2bc94ee9ead08884b1d1dae2fa27ac4cf2a93ac88301744a459bd140c2a7f81432fc873094f7691bd0ecad4f5cbb3b4c60153759bda931c951473d6a36f698fad92cf4539776f48c30049402782f079987290d36e434f50c2fc2daa1ba9539f4e3fa1d2dbc58a9c49999016ea0abb48a74d2c886fd932781641331bdd73cd6e488bdcbe0d6fe31f412a3ef29e181feaaa5735f2e691b77c7abf5d53e95cf8f730828da0bd0b77fde0c8d8b724272494c04d479b7c0da8f56fb18f785fdcaa8860d13e81bce4738e3ef26a03017dc4e1201c38fd10307b8149917cd5d6b2c6dc5a0275b61d186e6c38dec794c33cdeef12678e5d5b405e3583f35b013c310276de3bb90793eeb605f2cfcb25c5381a61217670c4196e472b474ec488ba3074e1724cbd68954cd76fac99514f3d24c3277636e01f9574684def353950ee27ab9d32b8473836bf50962029e8ee0ee9a646a1c757418a4783e0c84f574a0076fb501446e49e3f70e5a950f659ce982a0587748d1909ee6e5155cfc06b8aa37ad539228239f281785b055c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he03672a2224b9d4fc21b3ea9230c62f25868a9a4ba2139c6f847714e63087643062e22ed01b5617450c0fed2b8f5f6047bdc4302a44c4e9fa58f874e510913d85c529dacb7b626cc091144f0ab90bc1f251cd0064e984802801e1e36a2fc6cbfb862d678baf493f34db23276a3695ca1a3990588bb42081f715a5213df051abc8b43e0a98db491b5a52979c69aafb150bbdbb54acf27e4c49656f7a265799e9e46324b586eeb2acf26be5427a9bb8af1e8913b0d9996ece7411fa9a0c3527dbedf988a634024f616f48ad01885468c3b35ff50d5f9459be6925c605903f58115a3628794da4a2a5ffe9c4507b8c723b791684d39c61fc362f1d57205658c9f24a4f31e2001a858e0d2e7d3db4e2fc7cdfc10bcfe1bf88da4aa83955e367a00deed3c51e33e23e0fd3b91a02db1d6c47881945f716a1bcbe4333db4de11a86028d72b7c17c5d561cbfec25c61e9dd740e533924696ad02f128ef52bb536e7f7e63cef870b0de84eb451603e8415e64cff8711b40428df8d4f522b88e56f0ed79d5ccfb1a4f03e2c17cb3972450bc93829e70155387b0bc8f285332b148aef995e364f3ed685b23138f67ab7d34cb9f9c1d6317f3cd8eb3cbcb4279e54554ca525559e06b502bfc67a49976d1ac32d48a28b3f2d435ecc87971a52bc09938004aacb55fec29e24000a19f85062acad5a09e7a652ec1d5beda50a91f32ecb8a90d984a9fef6ba9d9998b5e49cb7baea75a152cf3b952c3728b9c267c00824e87d28c21885ceb182dc330e4208a2177969c9a10db2beb6398f17d0e092a245ef3b38cc9bfa8a8b0f4f27b88123d055a2d353c1c438b9d9240bc34788370d41bb3300fec7aae6c875dcbe0232bb057b7d31067e265e501c3e423a4af8a9f0e1f67650542ba9ccd73e85f5eea7ba91c8bf155f025a96be2c242295cb7ac7ccd8ad00c0015b3287bd9ffca405cb0c45ac829171255f16b9bbad8829549161962f155803e19f803a7271cc7a5d8bee9414d7f5c442df477a13df396803f568ff11d7a6b93a5acca4fb9323066d9f8c935f2f083740bbd5d35b2a443643ee247c986fc8b7f0ac838187ffea6296f21c7945f7254f017ecca24ea9bb389a9694938907cd5869746afc2be9aaefc555db10f78359fc98739376b8037348a2226f5e5bd62762bd48f61c338c7a46b8a1130106428b75abcd1cdf77670b3048380252ad32976d83f66f66dfa314c82cdbc8643f385916a4751e72e77f0996fae760f3f8a4355460d651968bc6e0b97afb364b1f1d33671148665054d77461a39b4e00561f0720b2cd542a94d8de28f2effb74f837351f7d4a5e2b2adecc487fd62341eeef3fb3ca48c23fff6f4be0352f7388;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf674fcc8752f620fde19019ac8374703fadd9d0a98b376688bceb69abce1961dc212dfe3669fa85f0b406f6916064bc31e3f54e1e17637f75c6d0d142ffff3be8cbf9c89531ce3f6c2a9c90167b7607a75e3150559bc380165a09ce874adee9bb1431bf03852205f00885bd8f67d62fd1355e0d555b1e251919802fa6705f42977bd8dd6bd70d3e7caea0199bd87e2de2197662952704f9e27fda4e2103df989487dc0ec29e2134ec5ff6e826284018719dbb4b5255b684480ff371dfd4490428ce1efd5d49d48c040974898f7d273be4b2af28a283a91d58e383e94198a985cb821ed55370790e7fbacdd8b11167f2806ea34e0414d585e557eb38046e71f9ae3e3c9e627a47b845566c32753605f538387a2c66b356ddae249f46a78d4d4db304ff3373da1e890e0340269d4ceeee92992189343bbc71391c7373d0149161e3ade6e9f1237d711c623e33ed57184ffbe0e97319e512ca08f0284d796fd2864d7cbc1268ef93da661f0ec16cce9e0d3a43d00f8d7b3bcd9b1099578e5b11970cb521f3d1cb2a6552c28e70ee19ca60e30b2cab2a6be4e3c63c307e26fbc2833aeaffa049678069f90670035772fe4494e380d2029ae41e401a36d3a168d272ffe0296d35a254fe28d57759ac6006b4d8db81f381cbf66282fd6ff46f3a2ce690d90821bcb6d9631b6df357cc11f5e6be7945a0cee7b6903fec41b926137dd999cce9ede0e6c7d79337216d73ff951b688dd534ca492b764821af96effed8542818c857fb62d532667462025faf6878ed95fd705ab314384c52774df027362e85e5d43aa009ec4c9fbd4bc43f49f10f41c65ee58f9f645f891d5931afaf517d90db3f3b67ec92390c1e9b3ea0801130463124b736c3b12d75647b7e11513b2e34b777102c9d3f734c30d57707202032dbbdc350a724148027f052c854d935cbcb75612cc17185035d68128d3e5814c1b00d5906c33783fabc40e94b8e7c44713d4e4c2d5bc55f8d056c3f48ad7a83535e169181bc6024297045795c74ef0d23b8f05ad8ab21a29e34aa26aedea5143536f6702d0c2b81e701ac191c0ba745dd565a85f7498648fadec3e17e7a83072e070d66a5d589817914f98cbc1121d9e1f036839fe3e5a14e99cc91ff7fd8234f66c310c44644c0dcb03107045fe7551c1cc0cf7b2bddbd2532d60b7a1ebbc72a6b06b30b1f41f336c7e5f81de44f03f49d6a2b5e969daf15198fe8a35a2d21b97b40771e60bc70bac0b4525587693b2961bb35ed6523ff14bde68b59e83f2c9d73a826e36205ebd3fc8edc511db45784628d9bdc9be92bd24bd2a72edefe502e8534860d8b11cd07b0ade6aaabfb23f574cc9a1cbad65e7577bb56520;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h766fa1914c40d907cbdb37c0c05d2c35ab01704c6e72074a2d3ccadb748d7098188721c6c6568f5357bc53bad032b58b5136f7d238f62cbee4e9e38dab08c842c127cab7a625463a504ab8d86bd74d70c8f625d4954e0fcfcc9e7f818985f1da5b4ab0bdea2787954d9c9b7c80320a11ab1d2af49b0d345f5bd291a8d7f1a09886b07aad402db9b0fafe65dd68087caa3862e6769d5e5e10fa49da3f87f2c8ba8ca146f1a98f25a635743c9c33e57f472aaae70be70de2c994a2cdf88ba5c7bfe8c44696ff2dcb83f3339e2b3ca335761b9617afaf1fce54972c0b4c7516b3ddcffcde032d39916de5f8a7b0e469001445ce4b66aa14655f9028767caf398b2d43207717e5b35d0897e802923e7fae582d6abc1a59c4ca727a8c74bc5ef92214a920f621f69d6e336bdcd32fd603e607495fc322f497769c73cfeeb5f48c58b016db58b4f2609bb156b11e96912f0c09792addc97543ef2970c3466dbb966706fdeee215641587786ded4a6fd5285a3cd1fd77e713e62d82e8852600fe6509b944087e3a4e73fe16c01acddb9aca14e459b69e81d28f048df711a096ad39904bb4fefb2bee4d591eda834d991fde629b32a6184bce75fadfc014ec33438b3b34a69aba8da8467abc84bab30939f752133cd0760836f99852da68294d275cb54c532bed56ad1bacb199b83e17a4ed2407c3d953a5f3e915041dad80e7645fc493b4b748a6690523d894598f217688e828329aa0828f2a878be181271cc74c8565bfade0a01b0f759be7265372d000d54ab27ed4f8a310a55709a13940b77a8e6b6858f06bc6b68184944b5dfe319c32caabc7927c6a105edcff59d8c637d94ba233d9f714ce13a995d8b363d429521bead4b05796f1b13552ff8e935f77290391fae9e2b51706a2d99b999fc9eb164a397a51ec04e490643eed0f29f4f366791cbfae6189d481d754adcde090a0239a7e72f660c1399bbf87e6f5cbe85bca6043d2f1a0234ed5ec073b807996401c80bdfdca71e159be48fa7de9d8c1fee33ec7d09dc91f04122e32e4582c9ec471abf65ea5d441704ba663d063a643f5083f35bb6afa2357dab5bcc9d17debec83f436d9ccfd335f02c430b4970a2d36a24eb22dbc4021398d7c807e4bd88145746a739cfb7853f847fd006d1cdbb9f3b2ad8f71edaa717381f110ac1eff7e7a4dfdd4f949125771b743796ee6f7f5a896d61c19be5e5ca3224bc2b862643e9c71b15782880f69eb53fa84f515881e62047af104f3e2231bbe11cc9e773a52dee48d7538777e3b9634a6d3d7a2724ccbe0df3d6c94b963afea8407d1fde723893cc6e66be5cb8b2b5e2665faf0b09793b1268366301edbebee4f5d047db5f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hab6ecc14041eca374ce9198dd50fef5199cc4c2443c427591a997da400f34cd6aa6d81fa268c0ecb6d338b767ece201b2e511fdb8ff53f1b523cad6806e6ed599be4fe163b58b166eea6d534517ad36663a906c599ffa7a74831a86b21367b27fd18486749db6888dbf985fe1a1a8e688cc0bd9dde359e752c9c1ec3262092dfd83b3b66252ae619405ca01f1fd1b99f3e619b87a9bfbc4b2ea8350d0d4f514b4adad15478fcde9d732fc18123089104313f9f30b439e9d2417255b4ee2b6fe47058498eb696ecc4f795be1f1d9501e3a5d0ac2f2463cef6d49b2f93d962fdab17314bc2f780a85fb5eaf4e86f7d8de3194dc8aa022a36b3d22c00cdcb2056f7360527bdaa3f5f11ee4e8d09a0696570291053a7b5d9e375826723bbcd5c1798926d2b26b0a99e947efb74036440122663354629ff8c00f57d4bd9b7df49fe6ca91ea789571dbd2fa3fabc0ca65305f7d47914001ccf5848858af4583ea51d64fede21721d3e886f04c83708c649fb7dab6caada05cb363e799c4b004833f33da41a5ca492bde118cf924cb5a44569451fc9adeb4ae3e7ea6553c7d463b7d7d7700c4d92a45e434a2bf0f60aac306517945ec15f3f7a9206a3c9adeecf25e8e296be38c26bffc6b5543fccb924d7c0d3b93e0874e711d6cd9542385af1102faf644af1becedb515253efb31ba8253cb7abd5794b8668cff7d20fca668bfaa8d999f0fa5cec393b0383ff8910c5789d0fb3f0037ff3339c3d247c9640e15686e475b910a3c899018f6868a634c6955a389c5dd5725c4c33f08a6e30df04b64b5a74677fcdc031674de3b410ca766f3da82ab77a36a5a657cec17a8aeeb02bba3826b1f0c43cdea9c56d5cd28fd7a6b9de113a9eddef118e7e3f4443920babfad7bc8f2e51eaf80f7e9c886968928f659004c7109b15682f62ad201179d98dedd9726abfe80922dc089ac47c89e4e5010882c1cb26291af2d423ea12c30fcf3a0d8856ecc3249fc597e108897a1eeb336503369614f23355ba78793b63170a82fe46ddb450f252c51a2f1795c55c82600f9d23d77463546211f06e3ab5a13871f7cedd3e80690461e9d9756593f3ed9564bbfb8329c57e895d405cc6ec49d97eedd1114ef43137823a0f6b77a051f8c19e6d3cbca311917a2296ed466d49e9768e8edf822fec0bdc14964cba6bb576ec88f7c9c8a85b3db01bd3e7bbdafc75230fc937fac4e8bff6292648d370724514db826868d65d05702f02e55087de6665c772f709d28d148e068993a2513a8f8a9cb9ebc93e8ba4ff43478a2f5a0211e5d4e0ce479c211e38767ff9f4442aa321fd8d8e69bc2b746fde8f6decdf979972fc6ea82a01d3832d8a0a475d4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'had8a36089c897641e2056804c981cbe6a3a0de122abc8e5ac7025d105335a1e6586b308d986a7de0f8767586cc8d37c183359003dae386dffc41977c463951a5c8c47750520f5ef9c7069b8ba1eeed3993e1dd84dfab1b1aab8f7a13e7e46952b94cf7039f72a9a459e13ac663556206411ec50f82f9679618ffdc0a9f01d9b0d9599db8a5fb0f2879b094deb16ec70644185470eb20665c0b4a0e7ba56fe7172f4e21bf14555df8e5090c63ec462709678389b30702ef7f78144b23fee2ad37f27f016c3d62ed47d7b44023c692c3d666d6ae84a4eabf8a5c041b2c47c675dfe0239cd761f4f56c9074bc00e1ae0eba8c663d5657887096f85f2ef4c0cdf010674a76dc615e4a84d91361977d1b153ff4e1f0a122fcff2c7597d8518674e137addaee02f72d0a1f1c2b21ee16e6c50ea5d41bfd902938bb3d63fc477dc7052a835833a9e101dc49a8e7ce9f3c25c4b8bc78f561e00b11e75d8b9783f0b0a38993881dad2d5dd58e70cc1f2568acf917e19860d65c3f9253edb46893180c348ea47251245998eaa9358ae793206a6b792d8a356a23555e03a310beb6f5c41067e1a4671629770fb19b2095919108cd9648d849e7e04c92b1ad9c39b2722da4fad29a283c945eef4e680961d2e8eb79fd1faa787f32744e9d556df22cf4955720bea31e51479a98298ab6126969760aee84f5e656947e69b9297b6292d4b4932fc90c1f063bcfb876fcc72e842d075b9d3a9bda7094d3b8e3b55568e7be31269dcd081693aa9a077a2a002b80a2f1e3d82bede361bc1a7494be49daf9e96c3e406154286d19f77333c4b99c2e0fe31bfbd59101626d113996fe2837dfb84e5011f5168f8d8aa8beddcbe763551ead4525b82185bebb7baca324dfb3ae35be0d84e901b100e4553438bdbbbd6c8db0578acb0fc39a7f2ee02955d9f85a928493e7def771335c80d3e1d7c32696df8b62ccb8004a020e2403de20d7c9bbd775e837d47a3f0d072be76f714aeb78294e29582c3faeb4b55acadeef5ab3c15cbd03a45bc74569f9def6ec730ec50b14297ef1003ef9a06f08150f76b129312e7ce8a6a9cc42da4fc73b7f573841540b3f290845cd59bed60b90c637c43f3b69b96389e9e84c9c62a274f6fc0cf80c863421b313f14087a018b4a1917389cbd87b4f38b7ef3bc38856d7f2a907cbac925ef8022764a186aa4c479fa385bf6c7085a6df98ef4cef2ef203e5a521e39fc5205f677ae06200fb9deff91e86d6243945bccd32a350fe6202dc709eed3bd4d7a77b9b62e14b34f961bf49e7d697e41542d66de3bb7c6992db979e751c650742ff2ed3b5fcf2ef9cf9620cf70404f0e7de35e0c34c3c3998f66d8b158de159;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h30d67414eddff70f0143827000fdd1b7812fc891c75ccf1c29862fda007fc5cb9face1f39bd555df95de81a2bc30329f93720bf1c66ecec50da4a9b5c79ee6bb783b2443dcad05e3c4e531ca95bce8bed5831fc7813cd06068b2859b79a6282e19d8ec1b3af6c1300826b7d6e705cac71d7b81dc5265df9eea0917aa57b28612bc80ae819a0972c1ab75b44eef380e0cbeb8e4455d167a2c290d21df09131ea825adfc90fb9983f0e243ed9c213b5a2389d1f2c94b148bc4323152ca6b11293b616259ea3c79f891eadb117474a421bba0eb2bba4e9bfd175a6a7ac7305cb15acb03b57df77fdc4dcf22ac2642969b57ad54a940113a40bf70543ce6d6ab51bff9a3b747c6d5ffb0c3d2e178e025005fd56a703e499d5583815169f74bac2b32dbcce48ea8bbe5a71f8bd75c379f82e8517a6cacb1bc3c7d9eb01c50c9fd5d2d0736299c63a2d2600033d4f386f088e982389bd4fde6036e35b0f9c028876c2b207d3de61b07c74b0be27fdfcd9a7acb63e749ca0b12e503ba44a6eb7f5af2aa7cda370b770dcd9c2e9fa5d3b2baae5d7014227505c0fac158f1fee8b7b3c45fd91af195bb0a32155e1fc77aa5ab553c103a097dc3ab298d3ca122e3f9d169061a7f9d632709e66bcde46c6598cdfc22d4a706086ae592adbe65e12a68c5cba12aeefe9fff73af7a2118664df16e4e3bff56a1f910a19eee9f762449a4002ce7a235c2a1a01d30bdfb0c75f6064c77d8fec7418646f9ad690086bff91b688f14fb76359af3b5fee47751a83f145496dbb9272330e05250ca2eb3b8afcb081acb43afac3d0e1fd2b59b917818a5d0e2eea347d1657603309c68a24a77c02e26b69613087ebc3e4abb562199edcc6d48e74a49dc248074f853f6e2ad8a6e75c0a2390ebeef44f5c2da6e62871797b64088ed72546388944977435c6305aa0cbd8b0af9349d9478cea8fa2564aaf49bfc0588df4c12f0590a7960d952226da929d8c64197e8b55d99489b8783982cda785177f49e44477b457216a42a5038508ab99ac7ed4b74d70a4fa92f6df3bb219c1adc0f4661feeb65d18c318adec8037d2d6d1a32e4e707ea9e1c84fcd596c2e8afe27a8e857966339ea17d76a36b4c55337f2880aeb9857255e00e672188cf7cbfb8cf053322e28a225c0810e581d47d16281c440d81fd958ad50201b38e4c946118dc96f22cba6ee2f53f31d7232872acc1b34d64c106de204d2edcfad3e0471ef898000361649cf306461287d8bb83b01cd7cd496ed8e421abb308557301b75c1341527696d7ced4fd5a7186ca9e7bce476c2ef3210b2d5b474aaf21ce8493070ff543b5a5f3c95912725561e97bb85ad8436b5da57a5a9b102b89cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h12e7ad9b4a9099bc2f51091aa3432b29e3810179cd1de915db40b311789e297a3804b842d3ecf1442fc0dad1e21a3ca712489b30fbcd315f9cdd26347c6dade317c483cdc89efe62da851754ca57e9704aeae8ef5530e80f61fa6d8e23d2953326e0b6f7de45e9da964a901df19f4bd1eaa320d55a3cddcc21c37b1df7d36433f8135d0c583a50eab0af1bea477ebe7865cdd828674cc9519f2f73329ddf75097d70b43bafb71cb578b5bfd81ac6d2a027a49b5a9e43b9da35facec3478c2d05b8eeb568e42f873ddbe7910f7c52e5d8a5e39d5c3fd41722d5e61ccf939f2fddc217b3974b6de698f842a0c8f97f851400a9a2076cdd09c33f11ce79f98742783bb1c00b12e5170df6c7cf844622f82d9b61f489d31ab93ba5b98b17fdd3ab56a1622a8b2fd774a8720fbb709086db0cf47b6ae3fa4a34b7b5c0b46fbcc8a942e9c66dc92f3789a3709c078392a92bf21ffffcd33384468a9b38bd1925c6800b19ecc56db8f8f5b4011d1ba4da5011c30f8ec5b13215c80892a4de9aa761c246247abd957079a0e3ecdbe02fdba233747e19d08b5b8ec1d151c64e112ca776371855dd96eaebab26c01d3222b7f4c7d32e74c9875b3765646c70e4125e940188f0c5c20c3ab8920ae94e5b3465162d45af5c625683007f784bd5402db212f4782e7fb57f0826c4f1fd885979bc12072372ad9b60b7cf2ce971668ddb5d76fb6744d04b74b7d0c93c3a1e35034391b18a55588ac1ff61c3b8c8441d083023a145753e4d75cb267daafb1af25b16aa098f5c870f8fda45275674acd3c9f8aea278cbb98f10dc6c2283ab37857e4c574524a1a5d64bc47fcd12f1e0290a336f180800549c267b5a6fd0977a229c6de81fe9569c54d5d442cfb1a64951adcdedde82cc0978b21bf955da095dfc7ca1397144aeb68ef9788292df9c32a7e6e54ad0790933c79031f0b3df79282faf2904b0c711eb260126de88e91c51736273957bcd8d6db2cc93fad90bd55bd153d042ade6ecbd000b58b08fe6eb743a5b0fd7bcc2addb7b9b54681d8e93665e67af3a9202fb0534784c610d57e9d86b4af6dc4e5f69c3bcd5b4105249259a99b0a7ed37dfb1d07d3296779f823c74e0c8a0ee7d42e63ec7bc0593b33b4efe53bd09f9ee757ca8bf569304333980423d6ff08eb587505735750280983036ff5c0ab44d5ea6b327f8300c2fe54097632b8315b69134bb9dc22c37a37b1ad4aee26fb216f563074f0723111a08f5660059f13f10b6b214aa35cc81334ca67bd9e6358f9f6aeb3567276b383c18cc0334544843fa1100f8101eaa471140a3ffa064bd979aa7e1a0e4066d1933737461f58e228c7168baaa7661a237cc0a37af6e5185;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hff496a92cbd7c25842a902c906b43aa8d5dbf8a2f084bf17be6c5c720ebe9b78850c2f6e52a92cb64dd6a90a9ef95e810ac1c070b61b88a55ba24d941fa7b19eb551dd85d309aee23e1d303c7d0fd7e04d5b640248c8fec42f04590fca5b8bef3d1e5c2da97cecbf45bdaa7f9bab98fc1caad0710ef69ae57db9bca0e116e217dffc6da158f17aa7e9ae89123b3f3e3ebe54c69cfd14c7ef510c6297ef1ec8f7e131d351cf809191326cb981d026ac7a3fcaf15e23e8fb9b5dacae9f63a08bc607c48210ffdfc7bd1442a0864640b856ab24b011291a7258f5508e948efcc72e0ca03088521b5c2df87626eaaf2594f28b9c566d7ac7380499bb0618dad68567cef289b9e9a7761c1f9395601d963ea8dc2639d658c655a3efed6b7ac6d5b60fe2598a0115afbf3ac990c336fa2d4125a8c7c1d064cf18ba03b0e26295cd22662a21166e6527abe2aa66cde1737364aae4cd3cace7c31c031165df332b8bb6e0c922e4e1fdb886283212f9237c7380c2fc9fce6a93c3642edfcb1f1135918de9215f82cb89a13d66e88ceaa2ab05aa033a26dbd12f76074ab44e5b64a1f97f08641636a93a8cab9aed00e5e0abddd94b90e7edf8e5f37144f7383649ac2e04d2bafeef63c2f90eae1cfbd1b7ed293f11d3c42a4d0370fb4783e5eb2a3a6306b8f29228296b8994f78d9cd9e88d4778da3941eeb4e4a53f142b83e402400bf34154acd8e9f69d0238ce6ce833c7ea8698ea8c079cdc91da847e169419dea3fa145b2052e20726c518f170a1bcd26c7ae1f4eac9be22fc25be69c5c64c651552ad45bac0d2b20918bd7bc9dd1002516c8ef0225ddf3fff5195ea8fa92be66c847415089f2982e11a9b96eb9e544e748531c3996a8f66860957d4ca61da5d1b294aecffa5520fee14de4b557b7a4fa4fa9dd8d2b0027e30de55214c5e300034feacdff12a210894b8f0d6bbbe1b60f831cacce5d7ef3e745b96a83634d9dd34f140b6fb2e52caf2d33359fea7093873b1c9ddc1de6c25ed0c76dd1dfa46486897bb7b1076c629d2c43808e28b84e96aae7b1b1711886f7c05f2be8ccf81b37d4f27871ea43547a74c1d1399ecb4cf5a8cb49bfdb6e84e54236a70edc376adefd06a7e01a7bdea142e0c104b9239ada0c5dbcd7a18c5abb660905dcfb0e8c3e552cd867d6899cd8d1c4405199a2d7137e54f25b9e3e9e7422f132277c92d785b2dc71a8e0d19378f871ca7686c14ecbe80d883bdd3112474ca70a04b85031bbb5625bdb11cd9968ac3b476645e7003ebf25c659ccd57d9f87b6cc539bc0c9f15c543cb34142c46b86e2dbca2e80eb3ad582fc722aaab81d4f4c6c93b05216f665e418424a6f24ea142db238c3de4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'ha7db35fb1317b2279f57744918637736730c95028ba81a703828dda91536f344566921cd7432dddecf50263b2c900b0e120de9afaf915369e9c46000dc5ce94c84037c2985cd4c8d34e87215e5f6bf2d61db640c85463709cce33bd2bcf5c0db1bd74fcf3699fe677112e57a0ebb82b8aaf6d68b8080c3f10afcb8c9a694a1f49b96e5a724f621cf8f8ba59144f5d2432e1926a7cf6f4472f27791b752085ca53d0b5a1d2c94aea3dfebb44d28a309b9fc629482ebbfc95d65acf0a456d985551c96e112d0d80e231669f1a6e10248bdca10619534544a564f24d059436c5c19aaddcd9ab0c27aef98d98ecfcbfe18a5e7181c7412e2877473a9143ed513e94dba5782d4fdde1f95da51d6fca039c3c06a7be9279301472e762df55eefdbb2bc1725996fc2a373f9b0aa564533f014174cfd0122bcc4b90d3cb5d72f2dff80f46821bc41d18e8af62a9ceca9885b4e7d34f14e525d6b7e302de4918ecd0258771c5557460b2acada7ba1bb7540ad26dd57610f6fbe8b1bfc54eed8d0a65cc3d1aadc19bc13c1758782f8a245bda35b96a584c75845bbc124b6a53677adaa0970b05f003fe6d9b019dedc354ddf7e0d465cc280f31621d06f6d156c4a9b91652cd5f573dc1cea435b7556bc196c856e9c4405fc69c9bd3a00f65a5813da14b0880526c3d6409300dbf1822c4714bd45a4ea37c3d88654457a6e29dab385ee8ec1145a9b33afbb62051ceffb3d78f3c44241eeb07cc37c1bf880faa5aa292695d12d4054faf69064dfed3db5c47411b99684c2905b8c620198dbbbd4bd0bd4d528d29bb9ad930812679407f38ea5d1579e225f3e80774ec73808a805ee880234ad6138d7ae4dd94e016ce13233d86dccdd7ad4957b0923cba0a9d7b34a9e82fabedbb3aefd8e278ac7070c01c20235d56c11e2aceb03a8cd61723d21d377ba668f9a322b6a30971b78e8b4aae34c1d95fe0a08f56a592cba4c3d06810cbbf2cacf0c0115ab71d60cb8519c0228d2bbb11bf6b1412013c0de446a6c4bfa3065ec38da1f4d6bcaeb70b5475e643d2db328891b3007ea3f5b827af8f2620a0312c871fd01f50bc35734ea0d1887744512080238ebab765481d920908957f8dc7309f8bd73108e5eb876ed7582502fc2ebc25e8db6ad7c1f3952c100968a43577dbf988cd396a43c9ee09924ef83302677419faf70c1f014821cb7abe45f5e159bc2415494d6ccf36a0a256440610de997e13bf3992ec9afb0bd436da9589fc72d92f48a0320b4058b82d2830f7cbef8b565aecf3ecc34c42ef967f83edf9bc2f74d49211acb88a4d37f6e40191645fe809c9fb53b4734b12789f81be33db4569afe09a3b39e2bc1012973ebad21ff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hc395bd84ad868989e4fb460dcba2359d22e375928579ee0a4280ae9d1d9cf5d346cf6644384d36c45f84dcc81f486ed558fda4c481bee1fbf43168510f6722e3789f598a3010491360ccc6ed26bba7c4a8fd8946ef558d6ac59dde051c5555c790e92022960ff626f757982af21e097715eb99d39b61b5fc0d3f02049097be43987622b0a4e519b83e40955b27e6bb3b508e98eb3dae90b171c7f4bce4ec109c4e82eb0fb90a0dfc0911ac6019eac105fbed30b96abc386b429b5ca2ef9fefde6c847f043e070f3160fe2a87a757cac4e5a5b04809c347c5ddb11966da65580214ebb8a335912bd6c6d8602f5549626219c7c895a1d9dc84246701a556f957936c40dc2f9ff351bef3d15821b1b117a9b299b58499ff914bce80308bb2b1d26b044e9839011ab2b5d263d791fac90f78c561781b2a784436bfd98e87115a476ee6f9a7d98bfd4df3e8fa2e597648f6890aae3bfb761c3f48571c35a15fc75d3651952cda7c6a8b0a2e19f2e0693de41ff7a4708df39201ffc12b51fb53fca3df5fff3a4c58078883daeef78aaa6687798659af0f4b0f0e505dfe02ff1a0ee607c0e935e143a2ee9e16f3803c3507e031da0eb842635fe51a5ab614baa0570d3de33f5d5130e4d72c9501fe288c6cd94398e8eeffef804471c5544af9f5e940db0300aacfbca7c9513d6f055d1a395804f832a4973dc6d7dc783cb64bf96e4b00242331fc671457281201f5780c027be7dd84f4e929a8aaf355f80718ee60ee3bc83967d2cec97311ec8cae620c716cac64109b0f5e121d383271ca41002936d5664594b7053d101e83bedd7b19f4563eced54205b679a72df1b345b6c85fd9df1ee09684731df71f6f94603d212998d6fe5f89995de9391433117575bc3fac3abc4215a223f8026cfb60aba3e1d4b898e9dd2b3007b1c06ccabaab319f8a19b81c4fb53e549165647a443257a73d254f2c2fe997e3c8ba60eea427edc2e3c3731dd394c4ec4a0fa7163741404e6d3481734cfa7ed73cde05d9819236206e1919ef621be677e76ff07d5f659b0b2fd5816324c3aeae5f1028718f56434c9721b614f04c70bf7144fbe568c450a9d132c103ba736f20bfdd95f1d85a286700efce40673332f3703b14fec0d0133751de8480879c12d44fd1afac48402bd9c58a1b6600a604541b23a9b9a4de3a89c94a1e4a270790e606fb1b4496da3e24811f0cb99dfdcac40dfdcea57741391290efda4a5575edbebce76f1a7ef84e030c5d7c4b64ea50a06ed3769df42df8e2989e0bb5db1d8265fd363194e13081382850a076e8f29b8c09ac7fde3ad59a45a78d79f7faa36c8c21fa33d392b76460e8f87d8f445c8ed44c15fbcf95b574;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h6f19c426a7ab26d3663b85ab3900af2c3388d67e2fac7eafabbea3e53ca5b7b386d20a89e216d337e333f11c4aa8c0b8dbbdd4ffbe0aebb6bbed11844d8d49dcdff5e56a40e8d051034593dab90285869b456a884eeb1745bf0814a10828542d8d83beb24fc8ec59ea55b3bfdb6cda79221a964a422e0c5034c6400b6c96638602b5d477aebe39ad202a2a54824229c3664f136cc2da0deb4e65195ef465c226d5a4d8bd79d6d9e8ba5285c974f0bd8db8bd034249791633bd7e977b7dfad0f6bdc688d2e885e3153459ffdba3a5b24a08e264dbbb71f7154f5eac42fa4c6c8bd94c7dde6325c95d7ea69acf1d33853a1f48de93885260975bf4a4db3c82423ec4490b3090c494132cf2efbee5860dcf307b6f6531de2c35df1a9c10f7e6ba3c7915394413e42f69703d2ec4ef3cf815fae4de7919faeab6088837e725dced6ee38e4093af397613326fdde212612ea5f502c3b754edf9ce345cf30f79a5f7a9f701b6ce3d63de107f15e331152b3489b23e5d4fd6181a792bbf3427267a596b6217dbbdf60dafe69a878db8eead55c07fe9619a8e6589152d3353ed26df42a8b9e9bcdcf3b6e34d8aed562574478c162e538084980b7d3c06891762635d8b58c80dbda295fed07767a98085e8371b49f351a451a14978350f2c19548b9bbb8575b3bc74f1e7c91ed7b1d6934aca4b46d6ab0497d87d84667adc0d871740116b18b4be35b8b7752b1601d2fec34e66dde6d11b7ed8ee5410be0a474bb0daa676779c183ecae9d1baab2268ab24e8362bf7ff8908ce67e98cee56f6a94c7493f2bdcbe188c012f54d264a477cea19d3850fec97dd7b2fae36ae6688fb4a5b7c73dff09f6030eb6dbb0a5679407b42eaf29dba87ea56b5aae1d13e3dd6b1eb85b86f91957f5e390e432dd2fa8760fc8c444dd2e8b98bf43173d052d17c7d5d35a47460598e8973e244881d3ebc7ea559e14bac9cccce9fe010103f01a88061e7e2717322ec0fe34643273b42c514e007b9b8cf9517611ab43ae8581a9afa73eb29c767feaeeb3079d000a8cf401e521b8063676bd6211bb973226f3477efaa1adf7cc8c2a51e9fa84a00e0f83a55433cafaf308728f5c800f70fc5cea840410a0fc310abd60c2d8d0b1caa101264f6ac3a8d92123214a33d121c7b426fe538a3b4c05187536ed785b2adf67a628e40163b3affe2d60db66a1496c4da39a0750eeebb4610b759d77dfa528149360ac88db9ffaa21f76d37acee87faeb588a973f714c7b7f43ea81f31371bf799b78776dad70a1c209fabc9da85a3b1b3642f56d2d88a1f4bd0d35b84855a3b224f565d16b6ac0e1add8e76a0f9921c81f72e20f92910f702518ffb195a276a897;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h80ab11eb95cc87a4693d9cedd7d52bbcc12ef76f1c50bf2e3da074d203e60ae5550aaaa1caed8a8dca42b720616b60c2ca836dc24c21678f7585265a36c4d1448fb3db03fad9a7eaba882a3ec49ef7d3a5f198273fdf979d8d3385509faa719d0fbe9dfbd332709d5323d8d1b7c63529d81e768331e116823279e74ae5b9c91968308f8fe24cde9e9494d752824a594046f73afcae5aa6de5a5d2ed8f44fbb20d48ada7a82c202b0be181c7d54620bd270d349c1269a42fdd3b5801e2635d5855127f704db6e9865e66b6f56e6da8cbe421f1cb2bafcc13971636cf352629118d74daa0ca98a5e1fd7186553a3edd2a356b9b1eadb50456640c31ad6850edbd1ad7c2b622409e1c976f05ee9a291a7c6ef5c519518bcbb464dc9789f223585bb46ecb4df5c5777a46313e0c11344f4135dd47be300e8c364fb17567320ef51c889532eab88056aed8b88d6de7c720d5288ebdd1bd80707ff5ceb533398e777dacca6de54b49ae3837ee7fcf35c083469167574fcffbf7f6b8221725ba6b1e4cbdca29c05cc5b91a36a71921dc2705414f83a121ec92037731c8c524d9acb530171d033abe610932b1e3e6bdf11517092e2fb112f6afda2d1157bc04c70c474d0e89791f6b53bc5f4f3b360e4eeb1d498405a5db6cc52f59b2b41fe25c2c664bd30622e62fd91caf35bd08923bdcda4eb5b1ff29f7ffc2a8c407213b6a60f1713ec417f0685e49fa826c8d2306a8ae66bacbab5b06f84de81b820e7c850cd3e98c6ae59e5302b3f644d5c4be6787c39d5dea1d15d2a2d05fc75302e703fa09b8708b01d2e5a469bc5153e27240c7479c974767ecb74dd870041c7ba9223d4372786e3f9948a4850ed690747bb314af02d0b40b0e8273804a603af4602353f4543c09a89c32f2d9e9d5af21b0b3a8b4f95222e31c8b9fb09a672b7827e96a1ad623b624fc3259dff31fa768af01219264bef9c0a28a2dc0cad6b6ecff6d26b81957489b0885038dd207ae30fc235bd20b778b9645adb502748443315e1d2bfe429c42dc675664a6edeb833c66f1f6eb949b3a1e7d453ee4c32010e1289db2060b94655bf730ae57495ccc3ae7dc95c2181cebca7771ad60a2b32ee33bc0ff9f3cc51e854cf7b7d677a45f12be6547a2fdee3f05ef897fd33c70a5eed9fa9bb3772b60bebc4b10d7a7eef2016570ec8ed72612f44cede80c308a785d770286e72fe1b144174e077f6377c1d11b3dae1477a3e32c3f4e99e9f0d177ca086bd2fe8721a9c297f8decf94dcbc3b4cfeb27ee2723e9ab17a3a6a1631ec8a1c987c3cd06588392c85363512183f4303946260bda1195bbcf3cb0ff700d2911d5ba1c17a15971361986af8927801d0176;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'had3f20347b3f4a1f92df3989799a3dc5f3941b1f6d89744627c6e0e8829b69fbf43f9cf06978e495f8d63bc59dc814bd246331773998e93e0ca610b62f87bda254ad78dfe85cb40868b54821d068daeaf0117d37552bc2b2ae4d6d5f117d6d7def82c5806a22a99b3611ed8787f997c3111d8a349f2a1eb1a7941b3f015c3cc0c1151cfe09872b0dbc610e6ed228f8e8d24a99fe379dce621a3a311f84f3e5949c9f74248961e58b75fff24a463f1ddbcda9f5c9ce1c33ddc2f2b2d21fe3b5368f68d43105f4ce81c529cdeeac5fb24ad488253538c27b769a8c3398e3fe3f943f7035dd2b90bb4026b61d7a6887143175f635611d0ae1358952db0e47f9084f3f4228644428fc0e9d72e70240879cca0d3cdb1056e6c19d635b87e33865b34ddf391709c59fa365e7c8e55e639bf556743e3803b99a628c7bc107447b7d89833dae126a5450a6a5774557ebd027d5476af6e15988b9f9859dd1b3d1cad799572d6fa598b783dd77c1298152bcd8cb536c4f40adb749f82b876fce9e248447cbaa736d5bb47a9fe3c5ca07a34e2c8bb3c7c4c71c9f57197bd627542c67a778ae8a496c463de30ce01127e1a871513f54a6aa98ac85d1c44bfdc1b9de2283259fef74937245dc8c125735aec2ecaf3ca9b947e896488f5a441c52bdebc7511bff6eb69ceab3297b3c31dac9378461d190d8029aa645493441cf486679c2f481618c7058beb628619db9acb9857f4087e2d76be7069cd62c0766f7ab868c088f112d873f3aa11bb529db728684b8b454a82f52758eb72561e39d552bf7a9e64ee38a804a5af03ebcbfaa34cd572e75effe515426385f62e585466c795b1de620166decb3e72f5409b35011c2d64073f41238b38403ded04e6836c3527be738000d859e30a93572b2a39d2a312aac776cc7fa24aa5242119862f91639cad573c93415d91d46192b7505a0df29dab56b10803eeee7a70598faa1e6edffb1e2eaea6f84b4e94160b48ea5bc1bddf335d05b48912079cf7f48877e773a46197b2cd9a453002267ba3a6b52ad2917d2c6add07416f127a5518f451e1af649d9d23c91ef1014f9b43f18169e10745b26c357a74a369e4277e56d0ad0af73f367f68f02d03e33f1c7e792eb01a3d6c2a5c481d87de8226764dab6e373afd2c891bde4e072e017f22b9cc0c9952ba7fe21ac4a2fb0561dd7cf26538f35cb734f66296f1c18e4db5b8d3c3cfbf7c7ac3ac058cbc9df3aebe0a9880c5cbd1bee804053a6c28ae5d6f639edb6aa9e9aab82587b16c7901af02b9fe4d08fbc359864bec436b1e0b02296bd5e94731df9f7f11524487c7046d560ec81af3e37dcb121806a6fd9bb7839e2a7a11e874f57bc1237;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h73a58f889f86f68666e276115ada44de5306f20fd1ce6d86773e3e4796b34b28e64c4259e61933c6adc924373e2be50e498ca312843d126be80f68fcaeec242acbb32773d60c5e1a14204476db6367811a335eb289f7471e2b9d3660f8e358937d9d1e0e3ed8fa5d1b237de6c5a3710396cee513d83bde719f79b6bcfc09441889035203413a0c42e49f2795543f7b5d99d2279eda747bf0be098ef4edef862dec48678bc8633531a879cdfde5e4d41d5ad189e290999891ec90bceb40f5d2fa31b470a584fcdbc1d9c4d8c5ff0a03e474202b724413644d3306bd475877e445fc7a32f6c45bc61a2e00ce94fa4b699f7f2c5705404e54e9bee86427f8b6c30717586d6cfa230ba087e36e6dff0250f50354c7c97b71156592827150939a6345e5fb2cc30adbc30f0f61fd6537ed7ca7d3ca88bcae4a6d2da4636d7aa2f68b85e6a7fee5473fe8a9cecba16a938c5ccad9a7cf3e980bd2bafa1fd2e68d1e3ee6188372020e3787307e9f4695c5b474e04e848fcdbb5e7a324b89a456b4d8b385cdacfeceeb89623c3fb5e7d45e5b6f0e164ea39e495853c850516a3e6fd85dc2c177533ca7eab1dcc6a7532b748541e40542a711b359d56889e1373b43bef937a08f93e3f3cccf8aa85b72f075521c7c8a3281ec41a7ec34ccf0c8675fc11ccfeba8a6876c03aa9a553c8ebb301a7a65cbb941d0432a3dfe769bf48ed06dd13581c5296f0084b904a7786b2027eb2e6cc50eb6a3f5ce7b400db2f907ad1d4b175488112fa89a187e02def7d51d72bd3557e0c7a6c0dd22783d29d861a6944aee35a9cea669600fc4df18443219f21a2f0365d67c1245da99a7314cf1963eb35d8201718d60782eccd84af59a8cab1a4fe7942238162c8df3ceb3360f5e3751ee837fac9fd58aff8fa48ed740d01e885bb4484f4c8c2ce52cd726a4b5e879fcbc9e6e7f7e7e11b004a83b0a181358df14a8f86f48a59327c76c9f4165dd88efc52b408fa5a57eb55cdb2aa654b3732b7394b4c4b219dabcb518a86d2ee724417d5bd8d8e7a2c6a47c19cc09fd137de1eaa8d4ef6e70359c87e56aa7395307dd8dca4f341eceea7e18f1dab21ab9292b8e937f5dd994b7194fc5a759a68fb2259927d8b142a1b9a5dd7c95e80efd36f0ef6f7ab9ed165c0a0ce5cc6ded0cb471198f625c8d2d9b8cadb4a39844bbe5a19d4e80555523bfd29377fb32997acadce215d78d6d6ccf191c6ae14ee4306b5acb7c4b1c8eee4a250f82f33749e71b3df2419968ca5945fc7e75d44bd4e1d021951f83dd5d25980cb5a14be268c5df3886ed17ede64d685c0b9f366089103018e04fbd84a38260b087993948fedfceeb7fbd7987677aa548831e4f68c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h2e18850d7fea370d8d4a1faff7d8588b3e4b2a510b90a8525f247a69d70c9aefce6ed74e47caca1dd5e88653d97ca546f1f25ef519f86d5f21a91513ffc4d873d54d604076d32ad26df207e13c316a05498566c709ac08727416d85792a5f804ead2cd5822e5df5d5a6f1ee4addc370216fc385668d2f5e8be6ee10c606d08e3c0efd99ed051a19351cf62c49679681f5dbf7912c8f31b0c94f7b934a004224aad94e4ad5a6bbf8c2205436701b39f7866c9aa8e47b26b061f1b5fa6b58c1163c36984fe7cea7deacb15ac6e6835bef3133ccfb249b6a6cb34a940f0dde1e8bce5d18e92f0c38778c37eba13fd9a4e915a1da0a5e938f6f034d0bdcfadff4c2ddb641767bc479c3c3fac85278e99ac3a6f65a61142358408ff1a80a9c24689e55970360825153d739520ac5603c4dac8e89e47fbca1a8b6c6f78417d9b286a43b5d16bbf045e0179daae90b6056f239b69fcc3fc6958dbca321815e0a726e6ed993ee7543ea32cb3c3c4e5716a7fdf92b6c945041f7f108953322937de81332e9a64dc971fae45f4dec605c2998a0b0e9d6fe80a1ec93209adcc90ac3be99584630e79bb101a5379cb857491d7eace6d5b50d58045db6f34e7a2c7e4e185d548a6cd2aab3ca6e41351e6cb28767a6b39d8a2ff27fc81f9cca7c3e55c626580fb9ccec1e8017c47c5fff44e86bb0fbe1781dc439db588cb8fa63cb5fe00ca536100208ba2bbb11283f43dd5b3594664a221d083a16a703cc18d30f81ab9f5d97b396aeb15ab9667aabc71a909705e15b9df2fcd3630f8e3244263f86a04d64404787fb4b00811774808113bd1ffe8a0a3022a1d39cc05b37ed2297b8cc25cf421373d8c2bb8a65656d1f3978668edc3a207d28624364f4b877bdd51924afab5aa2482d634de646a56cf684bf3a267462ff8f38410c07c43a0d0502d56e731335e2935d84e5d3b7a8e31ed914f78c8263b328c7cd545089a421174a23b24dac8482d613aa41f86c306acc707192ae5c336f3785a0e0dd049ff9a8d8501bb3e91ac0bd65eadb2a48dfaf68789e9d99a88d6d6b7376c51a6a7e91c437db7cd96cdc7527e452369bfe6041f6579d83dd4930835e8f7b93b3c896b7ec82fc3abd636b2c169a6e6c8856428170d8d149d519513b02e20e5d35b38aac36d5c4346b1ea8b4c25a8766bc6d4a3bc8ac37d390263af10cef4a7f89b84e1b37f5a8b279cf60b65ad8746548fe397a59fa61567fd97e2904e57281a567f25c8b913eacd3104a084e260180010abe9416d9466e162c41a9762768b33348747755ae14e16bdc927dce7b622ad733d20a143fce48071d204c2ece3a984f42b0554b55410e1a09010a14363078fb572fab04f1ab8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hdd8c70af17e73d31a0b5c8b1e2d8cd8f908c159389ee1cf6db5e6431946623d7da462b70cfda77849561a80c57d8e99281dccfe4a21fbae0cb32d49aeeba25906dfbd5da80252d607f28418e14292c7499e249e32920e020198e796dde0ef109836b9e9fe58bf333f1e56ce6ee0ca1686245e0b04fd0213658bce4ff57e195aa62c519a1abd027c0af96bf63649f9e4b9019568bd9143d84db4ae9b61236eb66d77c8535a4280715a2ce7186f18a35d332386f6a266f4f063c307b0e82511173620f06063793c9a2b78f6ba9aca1fe5fa975e6835c8d83604385c24799f47a71214e3e1eba1db0650ab8926ecc2eacd09fe06a85ead72b38cdf640da0a5f7ab445db8a8b45ebe0842e453d80696b96c17cf87e8d9a0a286731bcbf3228c2b4d66d4acbaa5d6dd04291666e5167c905ab17a471cc82be12c3f186a1529c5cac17edee605e500de97be45054f7a80befc9a9a1dd2bededf6ad19e93f2a77d7cd3193b202fa11b721d8952da49a6c1e44f0d87efcc7464d404471ef1ed10d41d53f61a2800aa998aa83ee4887880f595885ddfc5118aa77c814be3d9565ac2b99c21487cc956866a949fa5677b5f520d5c16b909d27f414c81285249adedbaa98897735c1f6cf676934a2a9330f7032e01964e70e4606f87b33932c0d4172457d5f09f5a9adbbeeeb5fadde90a2835d7f2b92b14c998bbf55538144dd1b25b48ed2f4feaae5f27d2d46857c038cd325d600b81d3e1aaeb66ba681ec3f13aced44c11e136e4f09601290a4c15a0dc9d47c421759859bbd0e12f9826a01aa38a258f49c90e0ecd2ff9cc9a602d851e9208b0ec08426ca7aca907c58d356007c77767cee131f074f4bda9e572f5e7e4b01ab80daf2c85e46f431dd3f49922d87ffe1c2267c5934b70e15d700acaddc9e82657a572d7ad44a4076ff3c47220fc35401581f303263a8931f235e78a85656199f82ec8a3c8280aef1410cac36c6ebc4f71f557ec690d23809fa857c154babce97354c27625415b65a5fbd60abd907a32dbcf765ca7b2cb31ec14bd8920141eb25c8daaefc8a3e4781ca375aedf55eb86abc44d372736d56522e4b70cd437bb70526cef380f030453cc5d112e2bba29bae09917a3162e5771d85bde5f94b8de6df313881f49be0ad07aec4504b356782b569abdfe9bb8a449fe74f473506f3ccb132820f9558f84ccecc95bcf1d4aa466138427fa7fa74c9140a4abbaf3a96dfe90685b2ef9e537aee25a0ac4d4a89a06b90a61c5dd03c2e48b2e67024bc7c3aa0198a3df510f3f34f38e4220602baa58e367265c7322f5d17e7ecbfc66836d572953a8a6b0c1f1fcd9d3de4a42b6d33e245001092b94acc3f0210ad4002;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h914e0a5780cb4ab7c5eb8339a985228a707a2b6435529b84063ae954becdd6185ac25df27239c6ffb5c663682848b505767b1471b08daef4232b02ed7f113185d2c6f26a743962281d87f74f8d5f2aecb72e5e7b3d85406b62c4dfbcb82ae300b6bdbc9cc2aa8591c2f43a41dfe348c1106238861010482b6d35ca9cd6ae7a6e6dfbfe900d08e1fa4376db55e442411df63f1a7e7c816226a89ee568b06b73aac35a03075c3c3c157c1b74207fb1730e2ece90fd54a2c3fa723d99e95a2a9b6d1ffbfed115e1760c1c912fbebbd72b3c9f7816fbdbc157c16a7a574070007222bed1206bf8994254fbdf457ece6e43c3d08dac0585cf1500f1c9c83cb04fa4c1abecaf86feadbf193462c6b6a1a2e8e8b53c7a355e1be154e8d1b3be30bb36b1a6dcfbf9e50252a3b55c209440cb28b078a5a0587bbc07ff2bbea01af042e1fa446adfdc95452b4b5cb526853ac29201f350da422c690f3c22bb15924542330f8126709c5d6434bab3a46adfb503565575a894bc01c8835eebfa750a1a5785914d590ada54e6f9d59c2ddb552680aae2f834e4de5c204e5f4b41196eeebf7792e3fc8ca73c714bf0ef6dc2e4f8acf9bd15b9e4993f6cfef78362fa914953374e5c434fcd71169a896b5062ad484461d20ab195c9126dc6ea1ae86200c9d18bdb124762292dc177344340c505234e62789dd85339bf4142e51c4f11f028e48372f3630062757e9ce9afe5a1a0d5c4c9099143893507a15b40c33bb1753b78fc3d123cf8fee9dea6b05e98a969d3ce49ab10c95d52db5eb4fdca698eaec71eec3608ddd0ade77fcc7f507f9284741408300f87d0fe39a23b7f912c2bca0a28fa7d2213e5c913bf5026110ccb3244ae942ae9b93b0fa8018599d184f2ce1d48d1718040537ee851c298c33e53bf5255883cb9987a013e1548a97a9ed7758b9e8e78cfcf8f8704f9b330ab42bd61c93d58a0b432617ea03a7cae897a4171328c2d8ef49941f36ee12e7be2f6c50c25bf52a7b47c18868f53ab7354d5e1ff42d04d10e2b1d20a236b8d28bea3a684b82d6d1a4af9544f269a372bfb7e227771d89ec7cb7f8eaad598b3f61d96eede30a16532f3552e077aa5358e2adfba8be883f05d8b87fa91012de3038577d5f0b47dc3d6100efc859b125ba5162cfdfdda869c4791f1cc68b61ef8d4c87b3c813ca84f86776cd56bc10ea8096b85edfa51740bf3999b2245e7af1bc0a8b10bf940ca463368a7842b229ae75c10853ee77d4375d504a096e3d659a527bd3be289c45bab1b2c67adea0e0053a7c5925db4794e8179980a04c74c93bc4c0843345cbfea85e6a54dc8cf79e5cb5fe7f25b31a29935244bf4aaa26d053d9c99790bb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h8018237aba509346ecacc21e7e771e2ea9c6ec73b6d61fa2375c041dbca51906c8a5ec3915fde6ec18cd90fb6f0d2c0d34e9d56c56df1f0cd97d59e7800aed5dc7d3e7f314a3858d05e770de195c4b5aa8945bf554f249e2e959c5f6e353a6ad3149aa8ce06bbf9f590ddd0ccb0b18300017d9cc5e22dc0991b345c9c32ce4e7cabd74dec692262a933780b0de377faf56d07b1008dd77d89de0c7e5497d332fecaa7a1cc741ea73b55f912127fc441adda9e9c8eecc8197919d3a76f764fd57a68f057026fb1493ad9f4a04d692136778ce26db74c5530f2d766b3bddc6aff579c5842135572585e50f68edc72b150b1d136c82b98922c414b53fd77ebae576c97cb02f3255c4e7222eac6c8240f09d1f3b5237481ef00c4b9e6c0111a7e6b33f5d6b7381537e06554428dd8f35bb9dd03b88471fa912d4f877f29ff206a7dd930540428a13b71a38cf0b2449c87e53ed365265df53b924011d6838ea270bef2033b7b98b71759b5b7adfeb9256a393b23fc3bcc2cf954cd176911bba75e5fbee9009908d6f5c7b7e688c5310964ead27992df7e42b09a2501db924aec8675ac2a8be77f0bd6ca2598a4dd9853669c0257b06b0d9f47b5b0681ef5237f8fa442ac7ef1df0d63e1bcb5428171ae438b5154443c6dc74eee0d3bdb3f5d5f61b88e9e273f05193f71a98f5e0a9d73e3a1471cf6be549f31bba060faeb782818f75697bab54b9169edcc562fcef144d0913727bb03740545e393571d0df39718ba78e4bfb092c752b685434d49dacdac8879af3dadc609879ee368ba39bf5a8154f6a876e599a2f73e637c80349428368b2bac1381f44227e2ab49bf99337421ff4986fc2653efe6bd9d72d82fd7289bfb8be7f9e16500991757cf6b8ad28f0714533cb24ca42f8eda6d4446e99606b2fd35cb745f7789b8e968bf9693d550eff809815150d185b2a67832106860fa1a32544baf5cfdc74f6099d3a332288c1e47a56198ae771ad39ff7be6fa84e6e87dcd962bc20601e97db8a901728fdd074fee74f6c1b823ab766fd5b27231ed0ffc2f0d1ee2c604af9b16cf2cfc33ffe06a8d29583cbd8b5a9cb16598848f98e51692162947522587daea01bd1d389102217947abf4fda59031a8431723f29de2c3f797e76ad410fefa060371e0a8e28d3181b1e32672620244235ac504d69357b7af64e2d084d842f2d6eb7349343afa2fd46f779ef7974636b48dd9ba64031767c313b13047d30603c50268557cae07d7f5fbf4a1a053e30d55552b786e51ef64806582304e1e194f2b87554e3d1c5ccefe348a9fdf32ea9e4e6a860f2e4171e20f9f1c9afb9621ba202323914b107e6692c96287fb9a5dff5617d9661a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h93647f8a3f1a2f98f8f485c6da50824b13d16e162a59e2a9710d4aaa0cfb52a8738a03002400f95124302554b5f5421d1acede8065f9501843d41f25e23e8cbfb5e10b9e462e80ef6e65c41fe4989fcf02783a69f8129aa19b91f73b12bf2aee48cf58080b69c8b3337d99d8366c429b26a41619e4573e0efa8cfa11aa1c5181deabde81e64a55c8f4396070ebddf15468547abb9891d61fc73699abbca5528b2563f3500d591f2cd980207697aecd7777c22b743465e957f63e819d02a015360049201942e2db8da696f25abf66e293dbbb7fa806d0b449b3d7a35ad7406817a0e2319ac50b274f1f9606ced658a59df6c8a774cb6365d58b38a873b347e501eee309fc0fc983e3b6ba1c8184bde7414aab60122d3f0c60f2254df6dc322305c38ef4b46d55f68b315131ed45f104e328b0169f8da661ec823253e7bea67247a38c069124b5d509a6c460d3eac47b89de3811d41bfcc46d008a0061e103f518aadbe0ab3b57ebe8ae92cc650f7d3c7924714ff9fbd4fdf9359e4874f025664ef9cdda84748f89694652e35760350e67e4e411a03ef6326effd24ebf9cb05708e37d88ad44dab6143e0e094a9228a1ef4a3e7f3aec40c57bc2b5bf0d31e5932b8024a6ae7b3ce44d08922317e05510ab58f39e4baa74b87873a66133686109995e39989ee8bdf4ceacda332b1e76ca2916cb91284c13d9b7c9c84c3da7101f2595409f9ae7d62742062cc110eaa563f92234a136a835228fe60227453442b4e9a9c6ad27d9082dbdedd3c9ad494a3c788c3f3da3733d02145137d77f6ae8775ee952e82f4148c21687ef2c23e20f8a9defec3e86310fcdb965fc1cc966397972216c317368994fd9bcb3ed0146ce06a69850a56f6a6ebec3a0ec7f858f6703cd594253123ee06d5ed89595a374567a182e8f4037e7a676f249768d50311017b0497633728d5bd63abe07ab0bdabcb1056fa80da5156a377a290f74be6591a4cc36e46be3de262de1dbda51c1f526e901cbf085465df4f2d8f4637576d581f441007b3428c356a0c35003cf0af79ef81756d0729a19106e19d33cdb17f458f3a36780d3b60532892cbf44a6b8e4d67e1ec1db2e53b314274332f0413f78f3c1f9fe180984536e74d718eb1256e73ed2d5d0294246ebaf026644c0e704c6df33ac5db8efa59ada073aa11045518e851bb87e68ece8cb5b3989889c85c4cc03f6caacde2ed2d07030f880a824eb7f12a6acdfdec0c82b9acf5420cfb0dcef2d2c054328e5c6c7cb1e0f102486ae8afedb9375c97b137c613a11aa62f84fca959ddb2adf406cb8043655711cd679da5a65e1e528ed260d86c5819fe39404e5fb57d30cd377ef2d09ca7477e45f60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3905ad46afc7c0ab4094e0ddad9df2137cc9ce856eed820de53b04d04b4cf77d576e781c0b637e77d9094aa14f8906bc02d75fe0b78b35247ff26b899c1a0e9078c25cba75b26a31a2d46907c1fa7827ce34954a71c34ab3364ae2c64f4e9af70d828078a90ef6cb4201ddcc0ced4afeedb7974b6288622ada2a57cf9b7cf558955e2d45834fa58c7ef8a590693267bf1c6f64d6ca99857658700dd66b047728959afa402db01cc9b4243585647d5e72f5040d03c9a5beb3ae5c4a357be55b29689114cfb2434d51b17f638885c2beb66c915d316cc668140fde1a1ef0dc1be3e8def89258984c28c859ff217b4f0ea8b62168f3ecb412fce3bf4293fd138b50b354ab1eb863ed7ea080227cf52cdbbcdcb2479ef69442d13221e7ad89198bdaf19ed4a5604cc26e142c7b83acade8198ed03152f01488c89bf1a3ccae52d8b38a9bd5a03d12ae86cf2996982ca4481dcf9720c5ac0da024ea50e30af29d57ca9c0e0bee338c5aec5a484ccb22e80b5537d0a994238a29f07792ee085bc23ed2545956e7b8c008c33d3116e345b6c3187ad5a60d9e4016e3a12824ec5fade3f36bf1236e00de6fb325ce677fa2f6d6fa68dda8edce180cab328920c801ff061125080d9d7a54d00998d1f3569726cc421aa6d2f43a88159a4e6144486e1260d71c0700cafc1339301eb7dd00ec342015eec14c585c88b8f053de59187a44ba037af6e1c9be5b5eac0d3b9598885d8dcd8837ce5d15aa4a62670a6710779e25ba6bbc28d62578df6a9ee08a669919670d883684111820a6576d5ce3737b26def3e8c455a207b7bd9e1d1a5ee1970ff17b9dfef014fa1fe2862ceb37efcef7784e68618aca86934db049d8218f682c3a12c6374f4e3629e8f4dbb44de728054008a398c69af0e21f9b516e5135032b7a422a0ed15d62db291b6307d6b04c9d4ac0af9c7e43e6e8bc82fae6aa238f147f13ace9228c8c2b90091531980c21cc81c95e675913b94c5222a3bac5142d9a484eae84d6af5c451b7e32e6f7c680f4e78134da9712d0c209b94f148802ec4df8f5538043fc2ba29c8d4188f1ffd4b0a026243175427c91e598a3aaf95a4cf8087b70c3d5732015f59a22e4129cc4cceb5530a41b7bff0ffbd36ee481faf8b56cf5715c86528a586e95b3f8feb35d76b2bd96bada270c16fe84e4bb76bd803aa8fbf99173c777bc8599dac70d372fb7569ae78eff63890e4f2d4b16c8cdeafcdb80c7b3b79eb4a83e74f90333873b54320d459ff5eac2b06d7cd835836887aed0688dad08a69e9ab1810e25b1937e0ad722da49baf8796a2c5d1fb835d622700ba3297a6bdc48cf0e1c070451ed5d25a15a44c66e2e633b10ad450312ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h323cb0ef9b8526a8683aef5269a2ea3a8e2ed50dabb183901d7d9dce496134787d9175b7646e6581ff286dbcd5a120891e436bb4897b1b77ff958925737177c4b4d2600512b1f33fb2f630d8b7fbc019b96799e7099deead75e117ab81285b8b6dedbe96ad88e1cd027a74c2b6853448d92371d0f537a2d2379e566c52659b637ba5478522a033752a310b2e979853d8626baedfce267ae05b6984401ded9f58c5940e95aa3b5b72350811b70121935f6cce28d2e31ba3bd8dfcb72ceac0e642790b905cb331660c899e3ffa1a9cc4c507e6b7bb66c9d5211016b2bb10e01c1e063f067c47b26b285e1c895bae2bdabb74de110ffced7c62e05cd08e86562636bc0fd4711bdd139daffaae7098142fad713467cf5194f8567a2525e3dd148dffc76fb3c278cf657abe4c045be7d6a708f11b9471d7f680f6cf593f2116b174e10c45f029f20535b1da62ce8c3efc17c35490222edbb85003ff029ba4258d27f1bc61a9aa6933c90825061982cf7705c64669e73e303c959933344ac4e88216f2d4e8996bc20a7629138869439a4f3e17e9442d1ea232489a5fd112ea023c7def1cdbd24d71044b48d775cec94911b858a481b69089dfcf525ad6ff00f344212039e2d593a303150671ca18512d5681aece86d26d47e19ae93c816da04c115f098673b418812dabf32fe24ac39fdf83e6121d0102f1d548f744b7227a2b8e0a12c5139b9a639bbc2e6bfd5ce7e02a95d94a150ba2dadf328e15f2e4eb0b73d600810949460b01b19b2a4eb7b37069c7f0247ac84e9addc3a69eb047db64d0b487f80fac79a06fcb131b54396ac6a0a38bc955577d55b442ecd5eb4fbce43d6f22c0da37d31204117472c971a5b7acf3d7b510ede744605943cde9d0e123b2d273e0771b081cd4410fa6e4fe7a19c8a8239c53977158379820ab1c55029109999d1ea870987db6a4331a8bddefa8be84124af565116797fa0c6934a560e483e0c88d88e110327956d441c60a050f5ab7d8ddbc1a4e45dbae8d5f7c91208039ec18ef21fac752539c1b6807c8a2900ed584ea21b016ddefe69908a9fbffa90c5fab389b3ddc39a277bdc31b398e1e0768a66c776de2118811df2a717f1b37c245a09347ef388be4a9be8fcc063a45c0edf39634f4507f19ab36358ae9fb6655d841bb1914788ee1a0a4b7223d3949a5fba29eaa3c392cd08952a2a87df5f970ada969d15ea8cca1b842282d35bca9c635af1780a713c0a62c272a5deccab98374c0f3f7bf5a31ec68cde7c6f43ece938f78ce1cf0ac424660bb3040c427f641d4833a1d01ad851af533d006bf380751f1bc9b2b0fadad22d455857f131ba5a999c1409856f1f349c32666fa1dfd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hcbc7cdf862305e66d01426dbf4a9364e05638057fbc219b19ae68188d19fb4f3dd9ce9f3745b5b556eabe7072a80d4f4d94a1fd4ade48db4dd30327d136714e3b18792f7ebba1afcea8fad5e9b52e6a5e0410f227f90e0941605dd0ba5a8c6114fec2183a9c833934a7abf73242bf501e5b392bb7d9accad4284e5e5e9edd61fd71fff88781eaa2ed59388a71a88ce0ec940600bf0ddb7c5426ca5abe67af936690941b09a8ebf944c04e32803e0767cb858ae9571a0a0bba2b1882a0e4f9338883cb7431835af9f8fad3e9088339ba1f7e179a7c9f6c9a6d95a80ce5ee957818740aa161f5ca6e717ba61c361e93ac425904ffefde8c280d4a30be27c53395f20990327106cc74206058f8f7fc771b45f13d0c1e1dee5b3a79402dc1748c713f771b2553d699e1dc422a3507b27e08a1faade90c8c7225fc892da56759ae5eb6a6bc1f79d56c088f45d77f20f2ec30ae01037abe326a8481b36c2e50361b95e1a55d940fe34dfae07d36020ee4d025e4a0d51eb54a09ae489087151b87d88288586f959fa79f68e79ade446678d83b9c499e18411821c1ef4fa5c16e9beaf1f2423c183f4e8d7f470691c43d5e38e4c3bf052c708cb399f9416db5d56aec995ba24f4ede29d6cc747175c49628c6f01786bd61318a86302ef496e02679818e9cf19179229aaee6984d4661f63e9b411f5fb0e886c14865f7f8de39ee9336579074b80e2dba02dbb0f8d43b96d984b7cd003dac75eac7ca69566477a4ceb57312eda91d6c7db357f39302485555f0bd6bddb7e842870c10b7d94cd77e5495cc9671391d61bfdf899b620e38899fe7504b69e067b24af843171cccc20b62d90b61cb807268a54ebbb54859b4a5a158aec2ae64f41d8a239d7d3775666ea7f8fb0d78067ea6db8d4d2c87a9e81c3b506d8f11d0eaf0c290ff24ab28958b199776d20e49372f9cd8dba7038ca35e2acb4eac5938db6dee12275e21e1a6f4486e50c5f104123938b7a253acd7abf6883ba699e78d91291d34ac839ff3fcb7115016f1ccd04b3693bf59bfb8a25ea198bae6b998d36917214a5b217b77223145e59bf424940fe98db9ccd890866657d4af784929c10c501e33906bc36b31fdaf4dbac0a2a312c360e52f50d34c18de34fc708735a504f795bc7924819ff77dd455e2499bff8fd01b50e6d79b1566003c19de5f3c405af1acc2396deb9ed4c83811621bf804e580489b5f59aa68275e021ec5c7b921ca63c1a0b2c318de14cc9582495c92aa200eb3d07dd8f420086fbc10597b7beb60d0ab12523e7089c93fc2ce19f5512b65351b538a5b25b74bf7a478db12107bc9ca1b69a30228900dad6580994267eed97a3d5d4c530dd1b29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'ha6e3b2c85674b73e7481cf353d3c04183590b0f18a0048dda8be6595d0e4d3ab60f0cdb5d5b7f74969c295810fae483e6d3dd43e23293b83fe6d0f1cf76d90722c231befa73eba06e5bd0309fd65fcfc639d98d1eb658a9c2bf663313e48c5daff4b9171821ec0d37d6f8acac33cbd058cc715a6277cfe130ce71c1eeef0855cee08ddd8161cb26dee76981e0463f51800d09e6d2c0300eb01daad593889c9a38c30368ff73004aa494958985cbecf9afd0e415cad987054dba429c553da2ea2f18ed65b92637fde8996ca44b511be2594fbefe6406be2810ca55f11d7b57965287e5a3b21b44e0aa44f3fd44832f9e8822df1573a78f543c7505411b918e528fc3827e8d199832f21487495d0d1f757cf44a6cc13f5359603ceedcf80338a55ba867495136423f18ccaa67b77fb6b661d1dafabbde690e2ed3018e1488a6bbf241ca060087e00193a2f0a6067ed2bb6673f5e839487224087e6e1a9d5a62557660d5e50d72a9d3cda5f040fda73e78407cbdb619eb8e924ff7102767b4fb2a7aa880bd8ce95c4a4b41e6b4531416ac3cf03459f48a9b5a1a13ca117e660c318d772a52d887149b13556739e076a536eb41bedd242b2322ce67b8f45aa2bdbe5bcd0d9fedf6695cf325863bb60d1349e3b003870a53a453284ae645bebe66e21783ffc4eacb9cedf232335a534bfb5837aa7dc545c274b84b2bb7effbc203744be4c85702550003e144841c024b231d6536b51ff886d65dfbb4f7bfcfe4c7836cec9e81d98108233461599cea9030773ce34f0e24078e54a064e7608051e2c54f5f6257c91c0ddac64efc102ad96f4417f740754ff1c238b199152605bc7ba0946824904290d27820e53ba1617579f85d6886facd261099eac4651f86aa766405083e26bcb56f5fe165c1157427d8f22479caef76a8319e63cab445dac183ec5f0a3b7b38cb07dc533d5d0bb3a5da508be990a63ef8f8e261ad468ad909f565dc4ed33fb44ba47ad5ebb1c060a0f19081d3677064448b4b7d122da938adf6c13c4e30f903296544c613b57e736bbd51b628c81d7deba894e662b77742fbd1c6bd79c2764dcccf3c1dc6332592c246e9e15a0646254d787af983ebadf23d092ba419a6ce6e411860c7b23b498fd5feb5d91c85073861765432ff6cb6f678e64aa509fd55224506bb45d82dfb584bfcaf8bf3752dca462dc185fb98984cfc140e47290f90af3a25e61e3bacaa09c386c40cc981e6d20e8542a3fcf5f839e4c934e1c9fc7666210a1731301b9775c75f04d086a32aaa6962c874732c83ccc9bb369a21d04ea90309998ca8e4ff2cc2ce24865abbc03cc94dda3ecf760baed3cd6aae4f8991fc74adc9b8ad9b0d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h65c773e6be98086a39dad0757e0e589b02e5ee01e116f1dcc895d520259dcad1bcb389021c2bab8223ab3642ffd925a333ed6963b565bce392c9bafe07ab2928b7cdf15aabbfb19b742d92bfd5b9188e1d04fa62984fc57aa029cd2127662eb7df2a630f9860da14856ce9a18530fd321bf62e3bb9149509bb0ba7f760ab1857dbeb5616fdbcc7a4414fdf77f6529566c209854754827fff91a39ac2f4dea8c63a3d42d858ba8a3e3cbf84915687ee7f8c5a9bf1e16f85c30dadbbb07da5f594cdaf9ed7c756364f3981ce6949ae2925821c20c3eff5c4147b76246dd67f879edf9b237a1c9276d87b9be63de71bad96cd437f47f700416edba6ace47fc69f1dea19c753f4f5721f4f2cefff3c93632c736024943de0e7acbfda95c6db8fe023a78779da266792745ffb03d0f6135b0c067294fbca80aa53ca07b28e2346b8e5eaf07af2b043bd63c59849848011eee4f8f40274ba4daa2f483829f026637bf39268402b57f3176df22314e0873135e7c5df76d57c18829b45df7ceb4417c10970932ff3daff7edab5968907db176333d5f153e8e339b0ac3a76b0dbe633b4a9a7c0274f411df0d9c8fe68d14aeb3b6417404d2de5885e79dd96459bb14e1511ab0db9673c7adcdc2cb81ee7094276b412e6636e5f65236058ee0106e7fe5f3184a0861af10b5d2667323e4dd95ee13a635777998d899bb830c974af836ddf8b48fce3b12148a7a1c704853fcf59b8b2a9e3c21cc9ad986d05c7d59c184185323199e3dd16f80d1efe720a38012ced6603b5d7eafcf2c8e515c6f1d9a7b137ca25495ea9747b3a41f21c6ad32450da6cdc8b57c67d9fafd3afee8d273826eb106243c7872654804668cf5be5f3f2cb8adfbefb7bd6671c774dae2ac3c363b984800bc4333414fceaf03b90357e5e1adfd86b8af7c55543d56d97db28d106ddc9942286560cfb8c214c87d584f940305c4fc7411b1ea2f626668bd61e0a11e1d72151cc1280884d85a864fff6977506cb1b0249d91f541e4285ece0ca1c717eb01c590859186a9dec9a14ee77cfcf46b2cba1b86b60cedca4ed0dfc239c5d5471174ae7bd8d90a5c2f9b2a4a551e3a99bb354b07b95c1a74c6bf266a21d300cecc19a07708c5b6a6fb03b0e7fdc052c0d679ae364fa7be887d09bec19704e9cc7f696c6a9b5f619dd2cdd939f8ae9a51946930bd84391691183b6bf006e305f6c9018610b4d8240ee3fdab357affbcd1e5e4828fa4ef0dd4bd5c18988da83516e25ecf558f38653cff81454b80072e84eb6575f692700808e8c2bb47f68e87b82031f1d27815d12504e2bbdb5c9fcb71596db9cfee82ee2100b6caac793d614101f95f6b15be7dff174296921;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h15ddfcec35d49acf1bf8313a5d4b1dcae44ce2fbbc626873368656342f3d3d61bf62224e3e13d2b7d7ae8ff58330824752b4ef23438357a73eb30a0af902aeaa6f8d57bac3255f0ca6a31d8dabbe9de4690b8472876536af736d0a414f04d1f06febab313d85b7e39f60800565bd1da73fe89731c49a9a7f68e55ba0b7536be3adcf599083cda81e9b4a5fdbe6b449bee1d88599b06112999e014f4ba255feb2bffdad2cb264c93cfec5e83c9e83028e0b4ac6e03d3afa244da666fe2bdb3527cbf869980fbf011e13da1d40afffde06960fb92261ff6949e84d37bce4590d43a8ae8051c09375f2a998e88f2a1e73d92be8862fffd2f7160fd853a35f2cd5787226aad3a0c09bcce5eb742db929fa22c96636db02f01ab85b88afa17f4961ab103af8eb36e6519650927c88e05a64ae7f04fef32a569c4a75168e22048f99d28eac8a848687126a80945e03af08bf51364bc0f4f37e62f6ea8af87e1736de8ca83366abc8f7672f9eb7683253ab4696818a340b8af383837e0bcd60c618a171f465a9833aede18381448ae81659379c21f00bb4110e47b7d44ce76c4cb0c4d18a71aa0cfc2c23ea686bcb26d3b0187c4baf1efcb501206ffcf76c1c0f3f87f56dd7c28203d39264138e2f6645598aec58d273c1bd300392d3d42f76b927b25094d307725e09b937a9715dadf8eddf44ef0343ca935496e3989955b4d454d155f043592a9ffeb60b8e1306b7a4f8f032a9f055e55f8ba04064a3792159580eddad01934b7f29ed9a261651c4f1413073a993123bd7338e6745a10eafd3551720ca2a808c2518e5258defe0b825897e4dadece84bb001151d64159258857270acc398a98691625e2b01f1973c4dec0255be5cd7666b82d641cab6753d7b4e180621b45694d5fcf56be15e362591250d51c8686dbf4ce792f7738a65874325780ac7af682d0d780ecd52794a79546cfb28980b7291e8e8136eb675119f31582630029cdad025bcbad506e73afd4ae7c75e117da57ec7d90a9f6390d307c22aadeb3e7f29f65996504f8acee95247af6abe3189aa212ece18e6580b146b809653ab421e83f499ad7973a6930c037747a22a43095bdeae3fde3c45b9856130a008734e74a797c54fc7a84e21be98564b4560c884b9bba44b16c49cc403ae4af801889e62581ac9d9c58171095e12d4c802264c90b87fdb089ba0836933480edacb840c66982320bbe8aca29db54851118850583abbd49c247cf094254120d6bb2a5794ff23f3f696d7a440b25e1865555f1564e32a95a112b512b33bd2b3d91b17f71b8e8cb6ce1892f0687186f6d13b4b9128ed2e0195de43cece7e84014e5b1bc3bf1b648536a9c263e7db021e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf29d9ae158580876227ecd5cd93e09f08a6003a59ef8270d1a4ca06851d543db767aaf918e33675315f95604f5f6925336d0060806a6cacaed20571eee5617222bbc71e8b8648f50007293806d2e13c916e8e1ec00ee8bb10ffedac830b2034caf72202652ac74ca7f8ed9af62d705088bd61ed6d6e9c11dcccde16b8a408a6fc1941f002cc098b55c56f3857eff2e9f0cb56f12f2296be94e6fca938b45c305620c3b71a902ddbb8f49c54175b02dca437036658986bfd7936b28df5a0c20fc20e93f43f7a412b33c6a6cf9b2cd09c0d6292357e336bf68fefa4c91c66086ddf29a2decf0934e05ccfa9bda838de928d1f1f6e240d120793e2462977265c045ce03686c7812d760afcb48cbaa19009869cfaf7a73c7874fe098aa2315dc4bf2fe117dadbff946abdf978eb37cfaf0294cffc71c9386a693df5d9a03fba03f9c781b28a7e7ac6af761f218994d115e7ee4f446f9c0aafe7177b37879b5ebdc1df983f4e55525e610f1202abd9c89aff74756844810fa26e73b4009104a802ccf1b3e49fd1df37a9cf2d5115b59821b2e4179347f0af956723e84a6c2b53d73bf49ccf826ed31877af9e823ea65a9dea6b9899e660b818e7aa468fbf94cbadf17eabaadf6ad3ce1775813bc1ef88cf2a0a66af47158b197541d0bb0c4dfe8964a6877e4ec0439d8f8ee2a7eda51f93bced55399b6e5711206eab2fa8e9c17a038b51f0856c239c64385b2f2c17e09bfc86d1865dca24336f15a0495828f0305926b5b75e72ed0890007f7cb7a08058b9761f4edbc39583524804c045b1a0abc9b329db3cce9064802895dc3dd71539073e03540d6111e79323fd92ad3040ae0a9fafcf692e20dd74c4074161c52b9ad19e4144099e958d2ce0c2c7be1a3e279ff877e0f6b2c4dd138d06258b300107d9dfe1509e89843269bcef396937a4304ac5ddbe9fb92fedee5bfa29afb484c3855a1229aa023a772036c55600e30efede0638c383970c1565ad1261649262d9c34fce48586f0e99cc5fa6d9d4687a681900d7281e6bd204139128d5094a5244f1a1c6ea6e3953239f2fdee46003d4fb9ae006bb7596cb17fa56d10852db83d6e11ddf78364be150ca06ee9e10d44c6475fb600119df07300c2eea651de5b9a06ffaf7ac4a9a8ada4f4351d3c9c58aaa0058b7b865b266a1dd00df32255f128efeaa0951dd2b57ef7b8595340dafa90ad887f1e5d4e27a7d4735b535b308631f1d5cbfe9623f0a7f9dd657cea40274f0eabc9dc00cd78c4bc1d11c48ff19e538d5744a2f38d8fd60b1e90b707f2db056c648aee8be7b780cb47b2f9707ac0629be467c705add21f290cf24ef7d5e1c234d289f311ce5d3f82d7776b8183;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h4c889ae20f5bf204f773dd4a3e5a6982f784b66286de47c74b80ffb657edeb365dc2fdf95ea0a015bb36a10a869afd6ce4d8efef917912e64a7df02cc81511dd86c92364c38c74c9ba6dd0992278ee5df9ced4ca94fe730fec3d2470d58c505cb2d3ca58cac9275204e436374c8cfe83a1222de4f404b6c8f29014b2a2ffb67a413e862a6b9e0fe1be37b7e798f4dcc60f260617318355574012e8c64430c57400d342c4cbd5ca940deb6309da35d8b1cb7699dfc53fa11f9fa33bb445617500dbd57b8af0ecfc1080d210a0c1017a1f49071c19480b370e4d2bd59002ec027ce841855f2efbe94c25fe2be53fd4126e491cc6b345a316a47c91299610d150b1f1f8b896a86b93784217f5668f431904dd042e451a1024e76c16a1567648b553a8b2f58daa2637ad8beea1f0798d75c9e02b916085fc84985227f8b2d02d34c780d01cf4e754973092971f958c34208429af868f2f7158fa13e317f064ed047d66484097fede3c02ed1bd81ade9c3f78c2b62c874d21da9ee4a36d2a638dc05a1eb330a38184843b856900c49bacaf613939d8131de53b09c3e5b657c561262b45f5697ac21d71c9d937661b3e19488b658e7a8e36e62029e84c3f97928d49815a045cebac85a4ae6c023d95b3bebcc26ef2716c83a8b2c9a61eff12202b2caf29e5050c0fd5f5e70aa6b9b52ed7283f3e676de9934106b830b7b35c0537b5b50f0a21f721068948ef5cf29d27d90c21f0b568bf2ac8cab51c297ab34f2177a98d99e5fbbfc18da4c6cac9a852f360294a9db3cceed3e3aeed9ccd0b710a55ed88966c98e3b81ac8152b6c87b45f8f56aa42480945356f37faffce0569e0e6b4ef8bc6a7169dd14643bdb06e8cd196b8fe467daf6b5b9b24252baf00d6c9a5e843f6d9111587a9530ebb51bf9818089b516237158913c66b612d671c220d54925c4d4ade2207938638b968594d9d080cfa7beab019e330491e25cbef698964aa2046ab22a63525f87a3ec8a61cdc47fd81250be58f04a7d77864cc0ce811827de457f43c9f25e55d758f6cdf564f45ba681a35318b0fad7c1604b64e8adbba777127b31b11529bbd306b946dd77996f9131c8c989591e5010bd1994b28569e8e33e618bef8b85ba901acd34599d776fa9a6d1573e60876b7a3728ffef44a1d7511bcfe5e39a3c8cff10cd179cf5bf940b1705afca146a949a0b6c871c5f6bb1d762079aed300ab168ca0f0a17155b7f29ee9f93ee746679de9d059e33ceebf2be4cffb08a930343a6a8d2d0682734cb4e80503ed44a27135bfeafa4e0148642d24831773ecd210718bff7eb783e4651d93b443dd649c96af16c5f5bf7436c502d1081ebc61125172574ed1e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h21ab2298f9331bd6bbcc17aff7e7974df608f0cab8242e19065eb7b1c0c5e50338c9f89b2a99c732c1a8e6470fb03f83654f0efc3a1aab6f6b80de4c3548a3e665866ea33cd5137e586c4046c43e92331fecdd5bca100b630c7c7994e11886fee98109a450177cfadc5a74f04d7b388a1e38c8bf3864a3c2ec246d763569417684275f9e89238ba43dbab2f2931ffdc90fc53552108510b93ecc6aa63f15c64aba1a4841490298977158a2b6a45b182addfb96c96f92943d25bbef031b3029f224c3b0a88ca5db7286b7cc7e21f0256cde70a2ca0bcf9ac80e870273bd84f4830529ce11675a5bed8ddd238b47ae9d0cf632a3d1ef2e209b7a614790d60526a1bf4ccde61d2d1b58d07ebca412af3ac23826b83f0cb3ca83238e6b1bfc2b8bba4f4857d770758a4aee16388749d2b745bfac2d6ed6e66d5aa1a1ace3095ddab24dd9a281b00d9436d81d7a5dd3fda3f6f5af9917312fa41abff2c0b0cf87b0491e858417eb545251b8a250de90f6dbb1133c60955ae63a4da970f9942abf7e0a803893841727ea3375a2092fd613b88f1059b0bcdf2e7ba27d3246e2cad576abd935dd96db07bc0a3fe159d6647f333707c4c13ccd495ffa7fcdd9bbd1857a5b037eaf9d7b2e1282078fe55dc7307f4eb0d49f79d0c1b2c90f27a3acd43c5d11452728752ca15061b5f49c50871aaf14c94be5b0b62d66613b097b1d81d5affbfb32d5faf9f4b96bc23b3b9d084b5aed07cebc24ff11fa76af2d33ec223f5c1e54fb520c154dc182590d2cc49f2292bc25f8075163029f395c766281068b2d768438265aa5e3725b357290325bd8512cefbc527af1af26df691ac42b74977a0c913b6943636193c0c7b056f1ebdf8cb29701a3a920ab5991218c37e0a9740df61ce49fd9ab46179598386226b90a7cf7bc56fd01d2376314f828c3c9ecc075151b9f7217d32afc750d7e8ee13f1452dd10a8c2f7b42414071cffc5fb0f98ff869af42371fb797404399ef475da50c3a39cb1cb4bc8688c727c46388c41f20b3f0397e2cb5055fdf871925d9ec59f543a8ce45015bab1fe6550b1b3dcd67903e152b38e59f00f93b85e02761a2ed368bcaafaba615910f3aab87b98a9686cd1ddb9780f294a0010ac1a98590d4881769603d51a3d248bd805030c2111779e14c233623c6067bca114923357556be783af748f30a41b1d099598ae9f774146e938fc3e2d4d2a2875ccac19beaa050a0488d05d28ef82b0770ab66b75ae5d57b348891927c5e7981c67263b1b1eeaac4f60feeafc2e0c9e2b189a74f4a4395ba95dc7854ccd75c943d9a43a9e0ade20797f55f227bffc3df1b199092ac2e8d0ccfb8a10672820d3ba6c50f36e55;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'he4ff60ae9263773ae17a09c978c99d4e2241466deac1d87f739d2eae34d9e26dcfb8efff6a5a70156c21e53e9fa0697bd24c4c304babde4b06caa295d138ae8355e29abac3fd557ccc1365bbeed82ac5da28c4c32849cda60a81ef26109f4fdfe909cff59ba7adcfdebba9f143f53a871f32b2988b95f9300bc2f30695a02a142f8cfec143ec3fa7cc5d91bd05de761cb5d13c8319d6a979aa522b4c230fdb03ec7e4a7e2a7e721a9b813fadaec257de82bd6aad3cd8f65c3db7d13fe9dc2abf703a07a8ab3275a7ea8870602f7f6868453c2ed785b708fca4b91c432483c4311a3723e926fe66edf1eacf3263c61542381428cfdc7fb299f331581b808d88737628944b7017b2f6f87dd0fd99bc82ec0e9df9acf2060d52c84de058da90f35a66227cc6a1af03ea275285f9f648a04e9407520932c816ac2e69e1ebcd479f0124c3abc70b81e3d5e54b36158eff21b71fd9c8353e9522cca3ef6ecec5f9d8a3b129ba3e40c010f67d94111a89a121915b3a6cb6b27c466452f84f278a723da5059bb5be5a200a7beed6c1db8a69e9264ee72936c63845da227fdf7915ae5fb7db9a075d0b1b27fb2b9d4dfd84cbec4b92578cbf4a6242226f87bb7c080404028398b700b52f4e89694b0fd91d8ae54768f67910a22ae9240b7b5829a2f5b279415a0aad8eda62081e873a367f1c6139c8d628b84cd56713bcd769086a812369287ef2cde40fef5d8e5add8e18ce10f26d2cdfdffa3c47b59b9552ecc98b1d495e7061521c908087d136afe93d6c7ab4daee664bdcfa47e7e2233861936f50f8def9d98d3ccb4622d2fa72f365f05e8ef16f12989b03066fa046fc9a6b1c8e192c8d70e549aa4059b87e36e6e4c44dd18019e6175fca17eb1f14c8e914a24dfef844822a51a255596e67933ca4b4b6e7af58a9e613781665f01eeb4ab319c7664e133ea0022fcfb5429ebc10d91333c94f11dbca66e5e5a4c77ce455e75fac65d5f56ff52ef20b97da89f75e2ecd2672452c07de330a2c0f1938c30c8b27fe4ffd6cac2b71f731f10e021545bd8b780173a425de696527ad0185775d85ade77e39a2b38c52b0ee1276076201bd78c981d46d1f0f740969eeae350c363b768dee894cfdf61d913696dd824fe6151bee3dcfd863fe16f3599e381f9863bb787c6168fd0805eb9dab356cfb36bdbda9a427b63fb9fefcdce762424f045a8d3528517efec3f6eb0e73020152a5f90d8f3f0a87026e2e4b1ae0f2f915bc2caba81d321667b8a3ad2acfd31a870ac2c6a12c7ba3532a90a6f52b89eb1c1f558ac5562a7ed517995c0e7d304e1f30bc92fc12ebab921c1ba7d2dc1fcc14912e6ebf77be5c41b16fcab86cadb09d4865;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'had0ae31bc282bfa231f75889f66a176be7ad5519fa75dc9e9267a66051ab638e051d1fcec3048f4d495410ddf8e49658024c75b8f6b46549723371ae0e9119e389888f615ee189ef55fdc751873893de1c9f6e39986646d91f60010a61aea06a74947c22334f71fb097a277fb52df96983984a6f3345cd31c60c12ae2513510b5ecc5665671ec534d620ecddd3ec9c523adba000db69b2bd6787561b1b773b39faf6c63c4c429541c4e2febaa2151a1a84b81c0f42096a257d83838121db7a47b01c8b53f4b630989cdda5dde3ef1365690b7f8ee5258d61cf9e64cf88815949dd6e4264e4374d1fd728031b21fb90376ea4430ae69afb428d86043517d8d876dd36e6afded34169cd3b64333b29f654fdcd165631735be95f846a6aaad4aef8bfd78f36483203347af1e41a994f38b7eadaae2e462f350b0720822e2656b1a5bf1b562bc5ffa11f6ec70e2863ff80825e5e1438511a8978ada08da116ef76ea6a8e281394c6827eec434211d86cc237e76ece221bf7753f3b582d17a5778670aa12359140859009e31f7e671bf71338920fc9794d57007e03c4e7473c59ef6318575026a99f228c3f9217476bf844bc47c33dbf35eff697c54fe597be02d5ce8269d690a6035100827536de6574edb46bfb111bde2c986dd5176a8a50582f5a5f3c81e13288e38eb64cbc9e06a7e119a7810b36679c8a681c39dfd2b1c1b5fa576187b020a14a24a2c1465d2593901584aeff1f12c5dddb9378033d0d7ae27969f0d9d8ae193c737b297607fc01ee2db2de52f2f34d53741604bbcf3cad4b5c1a31200d354c1cb1c8933f716b3f893c86f542019b3309fc0ad0f5632ac04a9aff2a572fb464e348fbc4aa4270857693eb57facbdc465d5019c2323c26ffcea035b4a0324c795dc039dc4e3f4db5051d354901db2ddf72ba9505e02f241b41ffa6e957271140168f686bb30ef3fa7f6b43ccd6f929e6e43b77230a8947ded5946841a27898d4c26a85288507794eea4a1d3b003f120f205f202a0733af82faeb1e3ac5c0210a816788db352f22bc6067d357076b079e1269c217676e149ea0fade3354dbdabafcd71313235a4f9c873af4191380766c825d5dbe8ad57bb9af51731ccc49e3b2091026a545d0589a80cabc5b3c36ded4f389afb184666f0d4e0d394a140a25449363fea93e7154cb034e4920da8bf394d01e4300a7026f8a0c41bd97762ad3b0a8dd7f433d3601052c2e266358d82d543ca74714d5a81dface2cb1f02cd4b46d3f2b058562f53ba968bb74b4a87f1cd270a1fc105c3f8a9949ee424d090e1a6a9bdf833508e717e7b81aa91dc36100f012ac5ab6a9fb52cc36f513caf8d51e53caece0b7741c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h7a81836caba96ebf1bbded86ed00cf8f321954293fa84b72da8866fd9ef6cad79f687ecab8b12193d4138f54dbb40386d5b12593f874454c5e7eef1d4b2ff3f4823f4d06c797c0f8738d32e1851d799a857b01f5e54aba11be6eb0820bda8a249cc556ba7e12e27f09020c08b79af2fd28e0b806088928c703bc5b6cf2ec2f19a7c7c82d2bf12c4bb8901d6f949e560304b9916938d8ca7a9b97796ba7601ccec763a38d01a182eb4259b54a86600c8f63900564a3a87ebdd2d59fc9780806fb6f594902dad9be7f682823237ecf8d9108d53da5d04cc6c2b4e73101d076e6c3f44a31af00ae88a6acdf672705f25055909e38e95231e018b06d165fbaab565cd3c8a17f7f66195387cc693b074da09bde79a36d7ee68b05754a9bc2437924b95025a51b5bdaf8035be5b1c2be4951eb32160e13c78281dcc2c2544939f5538891047fa15d8658ae668ce5d835ca4c9b9e7c7395efa272f527c84cb3f35d61081ece15ac7c122089812a399a3949bc123d5d6b04e6616a39164b134023b8677e7623dc7bf2f34bbdff9ad576c923753d3b1d795c6eb9fc80038e0029359cacc7c847a04cc103750c2e11ec6ef2fcf0dce50b7710b7d3cf69301efcc98d8d64486904d5aae6efeb96fe89efaaa44d91027fdd96a41e8e427df28734d7f4794640afbf6e1b387fd816bd4b8652d4c996083ffd5e7003654680f5b7ebc3f6a418d597b88d77059c4c30d15b5dfc0c10f5f8ce12ba50a082c78381d4dfb70a8848e357aabaebb81d32dfe8c07748be8b652b170e08f93f5e0873e45f3648d663553ae30d928e32ac3d2f1fe2e218adbf8230200729d9c14654d70232a66a1767452c91d9d2f79354ab11440eb8f1381021f32a5f98ebd2a73b4898017b937eb0169006a14d3baee0b4c842182430851d32464620486a9dd3174433967529e7a93d8e584c11c89ddef6a4850dd25fbe56d0fcf53f25276596b68297ad75791b261f1ffc6bcd4d92c4c66a3e11a65f1fb17dd144c16de095f98b790cd26525b257b2b1884de14db5ad9ce4ec984b73d9eff3f42ba12c4bbf9c7d8b9e08bd694db40598a445b0d4ebd93c077f8a028ebcccccdd9b7f16a4a64d2fc1a1edefb94fd9ea67884f1cbe901b72fde1c3c04586b4af402ef03ea2607dc8ca70de66f3761e9749fba2d3a1f7929f050aff34a022b503c6581f63a7692ce4c1f6a8970dc849dde207ab8392739f379a2c39d8e59f78ab9e8ee6d5b51218f74eda22274ae971d0355372d80e6916ebc529c5d7225ad565a7b22cf66912e5dcabd94b0114222375ba14cb0ff996ea166fb7abe3fcb53e141fdf3aecdad0a9c822bc19b3e0d03f51a3fb66099e480c910a6187f71a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h53c708a9b06d61de9e7360378d1ca2c160c4d28b2aa77ad65abcb89bbdc24fef72ca113c355a92c3f64fccc0906bfca278179c52ec901e6d3a3cd33585e5ccc7f69dda51ce059a2968592e018c2e1187268b066b4cec13dfc444ce231116517c2b4a35af33248148262b9fc1c6c9399597c0c07237a81e667c6e4f7ed6f2fdb980d4c1cf8ba12fe50241c4f92769329b79f2fec0df2e6e80345cae6de4d16c969ba6baad09c4523c69b753f02210ca12f034d7b2015f0046a3409f92a30001965dcb5ef4523dfda41f50cc7b61106fd4dbd022ebb7c3d92191c281649bbadb5141e5d3c23d6c3852bc0ec5a75686c3b8f0688f8945fe85d98ef2c5ca0b86d5be1f93cdaa634ab8d61a0c83652f52b1938599c0198c35756fbd18bae4ec569e53ccc967f04268ba3950a3ab4ae8353d6417dc1bc68885604214785a7b56d21a1d38106cdde26aa2ba39751917fc46878ed3d2eda5beb1cdb08b9c6e586b2ce373da502f1c40ceb15a12349fa0e1cdce4e42eb909def06e53b6f0f76cf4b92c65f1115db620d0ace35382a1e9fbc768c5441a938dc60d391b3cc70cdd878bc8e59290c5648fd56ef4e31ee1200fd7073ba88ea563dcda2e031048f66152dc9a9dacb8082a7e3df4a8d1cc40ccd0f9d42a84cb70e68aa6662a9b6c0703a72c151d536ef498fa2c4d3b2e2392437d6e7cc552f96e24dae95120b0b6fa675a90747f9b6d853c5b8338c79d2be5cbfd2dbd6aafa1dd7a90588e1b95b0d5c663bbea392769b969acb4441a465a5c936b275a3cbd108b6ba51ed93e2fd49ad87ed2611ee3d9c02a56939000dce06c34544df388a8c773948216fd43bd969d0131370bb353878a1f60d70136d20cd81968e3bb01d20a961c410be5dda7465a84c2b042ef1c2d7b5b49e08cc85f0f6db4bb1bc2b769b0bdbb2528c880871ec80f731e0126505f7fbf5f2be90f99e469678241628c87aca22ed452d21c40a66b52d977122aab85a71774f3fcd3233b4b88c71a8904c90013e4b8f4c841b39063f460f87d6a20e94335c1e1d9b091e6f59ee85ca0c4c191f58a195111a3227bc8ce01bdff97383e335d2fe1fbc80480fc56dd68fe52fe0f9665727977ff93cc757f9629661b404d9edb2bd82aa54b649051d183152fe8847100785048a57f074a1321057832e2eb65f98d01517c2d188e69845e0b50744e1da9b0c3ebe0ed342788459ad4832479aa6dba7c0c97a0cb0c17fa5690c3d661dbd73dffb8b4af85e1d621aa1e2faef30e3381ee7b35e34aaa1cb8d812a58340a77071d43fa971162ff62c3a48a1e7871f13724aacdccc8ad75924713849b07e77a0a2cbf56f76d1ac90e0b3f21f7f0b828c2c77effa668ba482a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h3c41706c78e2bd6531de1822699527b8d06c8706bd47aee6d464c397bf4c667c02942a17128f431e5f5391c5e17d2ded3266e1792c048963661852f3d5223fdd1cbb43da329d24328ef41a9323a7f7c15161bd4e1ce9a304daba336d00208b75e64586179cb3c29f41932f57e39f5612a6007344b1786e92f6a67a918a5837c4044b0c07a826436ce863d6f156e551a429acde1eb757e8815751fd9c3d8ab540b5e60ba1d55326b0f01f5db702da27f36d122f6dfb3c814df7f2789a1f504cce26af0a3f963a14c8b2c65862b62f34440ccd10e2b004c30ede97c99feabb1e5aad2148cf8e45bd67632b810104d583e4ebf74f34e8f3f2abea7c14ac4935b5a7dfb267705e55dce6a071cf43aa744a44256d17920daeded9a0f6308a885e0a08e57278ef9cc679bb8003204af5cdbc1c55eaf84998f898f97cc30ac33d8e12113907c916ce7d7c6c92b25a4863ff5d5b54c763ae463f87779d7cfa9c4268a47aa0162eed986f40eb67e67c376435337958f27a33e0b108d98cd8fc91b4b1e335f48a8ddb480a3b924ac8e83df756bf4fd91036b5f6bc6fd51050f52e4143043b50b836418f1f1c0072c20816c4f2d9248fc30ac74ffe1cef10747639af37a44f60c87f6db7eef279b786859ee50a6b36e28e00a0c5bf8f3057b8fb8612812cba3765c2257e36c846603396f558a1f863ac698833e8475f1fe745d6878c684b05414eaa175494702bce39933fdade9df64a2002c031e64962b776eede11c8cadc96d090c1ee6dd8842f1b344df31115a9a959a54452e02af132cd358d882e3a3fd44ba897048e38bafe0e3d9e1b358ae9dd5a37e88bdca4edef2807fba3bb3b660727386e37b846747457dc74432ec5f87032067e234337fafca77b053e1765c44b30e74f72aec6f6b3aab27c09a0581e39d743e0119966986cb92601a6dd1b144b10cfe886868d8536f778297695d93d2a74b33027eedf7a04ec3524766a65f9289e1962461a1a664c8b71148c3b4080171d9baa5d90ab4ecd152c3e9f8ea63df040f7ca957b6e2dc832b0ee76b9588ded075f87cb1d4bc9c02d131e6751d08cd76fb04826ebaf03fc51048b3bbf367fd39d2c141e71c1c1f5e077208483e439ea7a9c95938f83715a826bfa464cdd9705fba0efe0fd879dfabdd86087a9c7cb0b6b136b4c3c800d8312bde4e483cdab94e69922b9ecdb9d23b503342ae2304f2595cfc84cbed7d6f58629a014c448269e6dfabcd8fad08a1659558c5cb3508799e819d4b9560a36d7546d024efe2f16b3ef83c31f5a2e05cfad0766402d05c0921ddb5d035928ab1dab5ccb58da06d1ceaed550ccba4ecce6577f3254985c40636e5f60b4ad7650e4c74f49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h52ca6f2f084d8d435497fefef08f142b01cc19d5219e68238c781973abc6f6e2d884a203a4e453bfa87c6097cc273eb3ed6262d64c4c6bc2f94ae9695e21b5394f35d8fe0a1f6f2d6eb0c7252f155248e196f30647c7bb4e2ad17c4a1d98b0798d42f4cfae5f7ccfba1835b5575c03de56791b53d3b2844e63e29cc53dac5f3eaab51ea2405d0dce0fb4bcb37926eb158d3e9cf3445240a300ab3ee2b6b6754d4dbfb7e77e02cb59ff94872581228244ebdb832f7f27849f0a895810b6dd6050e047c42305e7c8e9f81c6909cc13dd38943db20622525418e752ef688736de2d399740ccaa53b4a99145d2398723cc9e00207c38d7d6de486ed8684e002d253c03f11b66f5983dfe5b8fa974fc030f6379c63d97985a93aa2045480b3958b641be8fd9e109bc786bdba003972579e264ef3c559f1a17473b5fba7a9438ed4fd3317096c67cd1801932790642b0f2098a43489e32c55ac9c9d8e4d546d593973eeecc7704ba090e950a415a4947cfcc7fb23d4dc3a49b3d1e9ca1132092af16c97bf3b6a43f640ae419ed0ea73a775dfbacf53daddec6e240b1b744b3cf650d4580747f0e62dd7732a6930f8c1a8eda1eac5170d7229aadc4dcfd5a508babd38296e5342756d487bedb493005772a6dee7a8c99458503e6c9960d613383f7c7b1c092b570b2e589994a8bd92cf3fb4e45838f06faf36184e2404e47432cfa12358641a61d0fc48a3134727be9cd097cec4bedb07e675e8eb931ca41e2387ee22fc3a071e373c0083b3e13e1e3e24d7fbcc6027f881f8b80144ff7caad08ca3bd30d01b38154c08d5b7a33155763069986eb91d9b48eab01bcc29cf74fc42c8fbb7f6e49988775c1001ddc710b2c6b03b3636ef48c92c5a4acaed5ac27edfb4069aa33399122a3d06f78f0010c19698337b2abeffd3daaa9af0274081676c39e2837fa0f8b2bde465a2da2ea58ddd6ff39d6de1da716857c8507157eb3a5f298f4643d660db50194dfd41a91c2721c1396abc6639c267d3ece2265c26053a54deb8e2141b815b97d05ec7c78a04b87e3336ed4f5c67dbf325911fea8b1e704662e66cce0adc32b5eae848dc05f5a118866b008ce6311c39a49e6037dc3510fd77c4d5e2dce8a2c2c11cfa66343fb40ded9f82025e3d48e69c9f0c811249bb1626e05f1054295e9dc51c0a4c83e14bd6a3be3e4e2430afc4fdccfbce55791068d1eb26436a8cfcb9d21c0dc7caa110fd58dbad470b0875d5ba1097f81e711749b1fdd145635d7ada0c5fb9d95384a7674406767c9a9dd57a9ae25b2bd87a0228d23e16f1d97e5608c08d6f18ff4a5ac0ea34303c517400d5a9798662d2e8c0e2c10723c44198d72383beb379cd0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h406094d01363f864758acd343ed061f922cd80422cc96032e15dd9aae7af2e364afbf7734709333eeca19d6ea5760b129b53b879a0e29a3e29b073c38bfd0149f7e3c6f953256f0eb3f7e2e0811c536c9a6bdd824884cf77ccf5846c20b29957a447706297448bf24614336de27e18dcad3fc307033ebacb7d7a3e39e545193d78b8f847641120e8b960c9a94c66105ae8cc70bb99a7f89c7b370a3b72fa558f9ff0415b4a0368b4b0e006908688860ac037230ad6cccd088b8f119daa3e5dcf7429ad79124cf4b81bb117050bea111c88adc86f80cbc924e610407d373712866f28f3863d53f89c5864c8956ddb7bb986433bd4a0e4d410fb3a73f67a6f750579af00090e828c574b6bb94adb14deaf2d06827fc0dbe6fe06e93f2e1855320e6255e96ce61166fced2dac778bf9074ffab2297fa932f9f8bc69c7d43ab379b196bb00221322f5449d5359f03aecab0c6ab1bccd6a0c6b7f6ea2f04e56aa2c7474f94e3c269f5cfb42cf4046a87d26cbcdacce450d6df69734540c82e44dcf6fa09bb3eb1b30173bd1fdd7652589336728e1eb74e6cbd8ef80e59ed702a99c0ffc1b3526d718c325d911c72ec4211ba46888c5f5bbb3b3a0470625f32a2f1ca72551a8b7489fb8f8e24785da9974795d81cbb2d57b58a187b8f62863eaeffddc8f1c75af1ee468d883c0478f7ccae1d5d3e4582d3b7deda68f833778490923f9863087f3b26d9492205a71eb06832ac63884df006fe15be18b92d3913c6a41d5aa142117b1350319fb8c60b2c96fb81a4528bb4cfd1869980ebc631db1d9371d7f11e4549d50d81dfaf718054134f08df63cf84fa8ff791c026ea250f62dfbea2d8a9ff8c19a3dcb97beeb55f196f433e126d06d836a27bbf8e7e10ea2ac03e44edf368ff772738897ba966a98562e365c5de5c4ad6d4f2cb8f4bee35480249f850cb199659eff2d6295d7120a9de112178d3e9e1bac0c93c287d676abd54c2f41bcbee02c772466871a9608c6b1d49da6f398eca54f89ddbfd9904e21b4d0f993407f9c67107295fda8ad2b30c7cae5a302032329e31d60584402a698fb93d05140ac7757724dc752c775b1b85a86242d7428d09d38adb9984b9236ae9d5370458c1945b571ccc0de06c35027878edbf635381e30966403178a97b5697c49fd87160d8481258ae466f5f5b9d7cc9a6a98d4d5608f19ef1aad24011ebc8458fa08151ae280578e3ee2baf231d7566e19b7365da3a95e4971879f629a2889373e6363825e5e29322b4e5b8286a65836c0ae36f0cb2ad14ead2f206fc97d5e7a508d0bcb4b20a813fac78ef721b0f41da3c8a79f57afd70076a07bfb56aa75ae6bcdb2acb5c6a5dac2f57f2cb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hc2033090f7a5ab1b8bc5387f81ebaaf8d7d700062c2d7de2fee09ec09456182c4b0d3a0a2b0c3b8dca659f8043b40de4c822e67c61d0ea2220b3abaef4327e1e6f70c2260e839445aeabce24c4f009efca93af4c7af45893f09f05a4cc95ae36df7a6374f3d41b24831c4587066471e22243e54ddb8f754c1fc4e017d6c45e7706e2f9f6684550bc9228d80693d1977debbda554c6963302954df77551087ca792e5e5e08500b851dd92d51aebd7cfcdc2349ec249b1d234dc0a194aa1dbbec77d3d2b2ff4b3c7f0f20dba109b0ade3ada7c12707eb881db7660ec4d10922b7b681b3952d6973c80457cbfe07178dbf287dcedadbb62e89c8684cca40b0f51741ef0a305dc48f6ec4609df3dd210e7b5709bcd9cfe80a3cad9500ab68c8f5a264d5af45f9585e94ea6e77f4e3bdbf8bb027b94045f9d4b54fd076311a6c9c7f760e703c26c3575a1fc66befa4931746ca88a67f874287f1fb5a1ea0aa6b3dff867e73dcc88ed5372d1365c474c44fc040832df60b67a83f8cc043b9d8248908ab311a0aac934acf8637e8b44ba31e47aca35c75c7aeee48977f19ac8c0302a9238a5629a0e4de64cedfb2b4a3fe822e2f22da95e953a8b16802a8500bb555ab8b22ac7bca3cf00e803ebe7b20591da360f932fe489bf73e4156bd59a33a62d52bb349264cabef0363b987c07fe2bccb1746ab3f003769b0b1d76c698cd74593279081870d51ec0addcbc48b35cc4d86b3aa05c7302b7acf9b2f1decc316362c246466373367ce14566a36da9ea3efa83ae5e4a24221499e4d9e779311c670170b11962cdc3d176db5cc5978bb3f62390260bf298f7837d1350b093adf40d502bfad19bb5346b3da2bedc28df5d5be988eb1acd16c3e8b7e4d0233bde15bac1e2ad01febbb0cfe44b8c49dd5118c89a8628d1901d8cd5f2d699cae7281bf4806b685794932e07c0fdfdeeeb6a36b15845c5e7eb407f80c8a88c32498cbb5b7e6978f2f0d6f2a847dc497cd6f010d89cfc8d918f8a12fc75ed2e8fd72bef0ffd648d6471e3d8c30651072fb2aa85a87238621fe0597bba1400450152fc512d3a3d7f3639ce491c6254ed39f8dd5974562f2c0b7cb0de28f0b48f4908d3d765330e9dc67d85b910472a6949c384a9f91893c6107cf2e95c9ebea1d33ff579b28b0a8400e4df3ccd0d7323d52e4d3257803425e4ef91bf76369c9d8a8e8d661dad654e8c592b006478df78c88dc170cfe866baf23a5ad7b6dd3ab1d92a6ceb061ef3c47f683d9b0c19da06f5062642cd260414d1f28f4fc71e9ce62ba8609745300b7f4de8f0359e67b9e2f3cc15972c2d3ebd8a87e49c7850aaf67b9fcb572754948b51172bd30c56104d52c4aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hce6d4d868af1b82d9aa483b9d1fdbc8d7b59b0beda401fc2b77efcd61e4e252ce8b1868c060ab2b97430643310864547fea542a1bf55aac2c246764ca6d7871cfad6acef88531d52562421b545a4a6adee85b4bfef3b7fd2c084ca4a3cadfced3efdfee687deb4b55e4e23259091e9735d4046264dc916bf3841e32e04051c8b38a5a461743572bec8cc58e499556901a60f5c8c0f0988d67d4ae9ad54c1fd5b2b413a26fb015ab6e7d2c62bf7bd0aa0909dfdda4e57d413b7a95e0dd83f125418910456167b09b41d63129008ede7ca83d6b196ee0d071a1878d81f531bce00d3b47053b11daed38569ffe675e82823d8e7de36c759f930b7c6ee169d84b61b0b6d7fc596630acb60c88bc6af4ab7fdd8a50078e9872d0ba8265653986c9026e9b9ad29932e9207fe1c416dfab41a085bd384720239853eb8687ece15fbb0bc4fb8032b753fa95b95df7b931b2c9c7ea9a24455c624ccce59b403b063ab749f05da6da712ccb47664e7a81f8fb5c5bbec860f598aeda306a5abc661dd6999ffb01bd8d26c515570095e05eb44c4eda072be369ced22bcfeeda583137b1b79f4934b6474f491b28b288492b93d0ffaf6a0e36e0ca112874c5bdbbe87e83c4f38a7b44ada68794e48b44a46275b5afdbab74b398a664e9aadf0c0bf3545c054e7c65a0bef718fb6c6fa425685efc78b9b156bd41958e9cb6620449f2360e9aa377f0cefb291a976d0016dc62294ad6d8b04ab3b4c4de13a4822f0f3af5ac63a4c1141050a8086ade5f915759735f416efa01f874327813937814d5e734f4528e552970faba0dbfe09e9cde8ea044d1c3db8a07ce355b6a86c06bec8a85a2c0ce6b5a0ad6fbb1b612e844cbd54c3a180d60eb9a8022aa95aa9a55ae8e2291f95bbb7635bc299e35998ee43ccb4336c399443bfe0e7fd3374399aa2edbf911638cb2b861327627321bf17a4b64ccf488b6f6714e21d2390bdcc03f14890629f73f015d5780564fa10938d2a3056fa95afe58cbe01565170ff807f5ce8c18b79651aceb3beebadeafad5a28c324ccb0ef67cacf275520f9cff5127071206e5af10f0f3ffa612b10dfc905d14fc84ddeeffa78972d3f96d228bee3b2680356ccaa7c90d91a3e02a5eba73ee7c801844ff321c492c726ef04e8d2248474dc4fb141d3d8af2b08874e84fd69bd4d3085687e58c71b44e446d1b34adb3fc8870d2b1bf982b4eb052384abb8434f52ebcc506fe0efa6f8e604c6703172643b89fdd9d5bcad312ce223cb3df29ccc8cfd31ff4e2a32ac11c627c7acac26c9198dc7d2ff8db8fa3f1b94bc68e5afffecac5502afcfc6d2f3b03c6089ed2e92dfb91954b42f6f11b010e138a88596ff8a0ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hc140eff82390fe4eb170c645b597c02e05a0e49300a02bd1ff44f144ad76d96cb5394213542dce6dfb1803d49b4f8c4b6ffdd11fc6288945f08ac0503c403444fdc780900243050bc2678eab06103b9402661968fdca4504c8697d3e76c7bc2dd6dd76891372aee3992685e8ed0e15c51cd265bd87f4e64453e0e3def1ddb41cdb01aa5dd6069a337d41f2952ba334b72cf671ce018c9edb6e2f7dd6bbad69c9e518da4fc571675403b347e7b0c32bb99f8bdcd5dd3e380f644881a054b41e0022557dce62da67b76b024f4e2cc2987f082517e2e966499e3ec6c761bc3c59dd3a99e4c9bc1e7821f90ba90e814df08a59d1183bec87bb01d50c3f585d70d18f9c2f46cc1615d697becde154d7b1e62ccdd3d44ba6ddd7d1d55cbd6f36bb40e737515a09edcc1db9c2c8f6ba3b3c51cef86760d0ba892400ac1bea97bb16419207680f679f5a1d6f00baf824cbf28261b7776250e6cb98c8297b698108e4189a0dcca9e42b6987dc088e6db9fb929e298fa7b06ff75579759dad9bfead2422b3dad36face2af96480b203c07d3312061a5ad3314e497ea447590ce271859e4ba2d1dff0bc6b382e548c8feb00bea3259d4aa7a108badc1948e69f1f818d0d0b57382198004bd59f08f5803765ad47bbb0c8bdd0efc3938a5dd7b658750a6d831f4f4a24eb68e364b5382d3a5e828cb6e3546cf0107f74cf72bde024df1de6565f10ff6af197397415db2035570e193a44f83fb553210aeaf6f2f61521ff591def392329b4c35b9baac1c1a98b2aa38381bfbac18ff47d0622741277fbab87934275f1fc6eb586065839d8e2f40664a7c09d912d62214f95f328cfdd59778b4fa7a5e2b85c68395bf51415a99d6f263735d521c028cfb6771495954c66c914bc5a05c94387775092c0e54a3d877ff536737cd96633e9dbe35e95174ffe881c99be57155a26f9d9f164906003c27e16b0c385f2761e4c9245100d8f79f939d7a1eb50f393e17619c223000544a1f161117accc45fb0c224ace9b28ff3168ead6548ff584b25a6964311262ef23632fe71434d5cc8ea53dc7a74322a7998f2296cced1e84d91108c3e086b4dfe58879dfd3c9ca0c4d596535b5f420e40c12a706947d047dbff97a724c43cfa50049fbac32871cc4ef6e3ffa53b0b62cd7b8100a91c536c73ccd5f97678d0c39c193c172d45087fd42e7700ba185c57d3a745bcd30349aff4b1b0b2b01a1266d803c612a2acd940ab8a626bcd02d1309a7ab605b36b1a5f7b847fc17a401d2bf91e98ceef5eaebcd740da8de91e37b04fc85b378974c936b36b8e16d0663ca5dd3ec9484e2243acb262a98f16b032a92171a980b51d108b528f0ebfe888dfc1d68;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h76f01385332add6066d0db65b0e4734d67dc094bd103461f4d7adc6bc16ff9556299db314151cb648c8ab4c66573ba5ddff4bdfa80e2121e54fcbcde191fb3505b69cd5c7f3007adeb95e0fe765a4dba4a65b94cd509034a937c15f122d134933b270e26c567cf688bc7912465e53f93923bdd5432fa2e346612b412bff910a6f9efe67467b2c85a4080f2555739bf8168127b1168283b2491c9d729fd149ee9562724a7dc1c769deb5f2f7906b19c5812796cc528095f24467a650f3dfb3202e387952c72163633f27d89213c0e63448e5a31024a5cecbe9d6a759d2c338c585f404d31b1d91cba475ae58b382659951be1a3049d10ed5b7359cdb47b8216f459b8732f37afdb8d7059f5f7306ea5d458482f2c1556c32eb6e56261d50798c7b767f973555813315cc81a57ba4325e00e1d1c806e18924051f3139cddd95c9fd4564018929dfcc617b3f8de0d1c70c32f7627f5d594a0a3c075e9e9ba4690d435be035744605ca699360dda89b485ddd7fd6d41cf0116757ded95a443fbda48fc523bc2024264aab8c6965f6e1df80ce07aa52be2021a68c4c56650681296fd421b063973a1fdce7717f9fab557cebdc64ff1bd901eac1732b9162fbd394e9751b390cf355aaf93cc1e1fa703f2a04a864f7624cefff1470f12f49f5cfbf6f2fcb906d97c2fa712a6c1e998dc92c979303cb774fb2d4323c4f224f6b76dfa1f38415cb1d38556866bde67efe785acb1b5c36f3b1d97eb6bca9e7e9bba94be827815693ce9e0ca601d41d7267d565af1d50187596a9f7976b0c7999dfc71fe0936b8f626456ddf78147e48f4c55b4daa27cbebf18564b5b9fc52a612c195bb07ae5b7b4ec54519d5ed73f4191b1f5c024f66e0b5bf721a264b0780a0240d4dbf74511ba1f4c21b33def1a8db01418c4e028be8c1af1cc8a5518d59fdaa8d0cb1a98f96ee1510dc802f3ac190feca048b25c6e65b7b3ddb58a8350cfd5284720d758d7a9f385faef2b7ecd1bb10673e827f4313bd5f7c1c7dd0c39fed1357d130efaeb174a4996afe20ac7e28b1f2dd049ccdae607a231bc15fbc7176e0baf10349bc68c395900758618b71f24ff0edb794c83fbfb977205badafb1b6a258728b84504d4fb329fbf878d0b9f3a5d7269049820eb54caceaad80e66d9e138e1c1355ec25b9e97a1e22ddb37c60d97e8d90f20011c1086b3cdebf9424cf1748d15a5b59cca537f0d727bc6902ec303b802be3f13d1571c79fdeec1b08e7b8b938b31060462bf8892f6f60a40e401553a1539cbea14d9a32b3e3dab344cc9f4aa35adcfeea9d2c75ebd1940903db8f7b9a4952cf83f9da18f845109d18fe789e47de514c4fb0aac8880580ac8c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hc5afc1c25f1e360c7cb5f0e70ef6e59a5c72d6576157a908d6182a7b570b0aad3905abf4548b2ac6fea5bddd4634a8779619c0d5c279fd0a0c3c785a9fedbe8bdc74a4ad7b1395678111bbd8f2f787b495119b5dc31395e434a485eb405f07acc2665039a7eb035dda146c475bd3ceec369179919a982687b6834f82439d4decbe8559ed9df6e473af39c4700a388a18e4b02854ca4e8915baf9aee6ecdc36f8ec4a4aa51f3f19f677271f1e3071becd2abea26142f8710e6cddfc7c1934d9e0d771d19e9c1560e24aa04b6fd5ef2a41b9acdfa982207bcd851e682132ae793ff6e148201c3a6a532f920de5744a6225a44cbb6ac38261f3980b4fa633d343768486d7e12a40a1faba4a5eb0459b954de39e1405335b876b09a8952f93ee5063d4e62e464e54a40ad881aa7df281962484ec1f198f17a1eb297c3280c002caba85f32527f6e83ed1b382feeeaf26f3f32fedf63728fe054b846596db670fec8f398131cff52530e20effb834f4a6bf4df2b08a99045d5a8056fc7a57eb689c35df65b413fc4509818e9be776b01641061e4f23c1b55a2a8096998115e21f3536d310f55246bff9799af7f3bfcfada6d044b9735e3371519f37395af6256ba12adea564b557140b91de64398cf41cb9227e0375583e97eacb5066d3f2524fb00b8560f4e02b548869806dadae916eae08629e16fd6d67ae73af17d1235bb49d639d5241fff6be074fd41ddc464a51845442336fb69d2dd921a77a45ffe5481b2db1d98f287ad383d12866431b527d496af6baf89e8a49b194f9658826bed8f2bbf8525b525be194236afa3094756de41f0609fb82d25ad473d18a8a10a01f2995c68fdcdc17e1743683fdc0fe02614a89b0d31d53ebd9ba1b491f52f0d73c61b40fb23d4a719413a3f638ca5527944e0ace5bbbeddab33f0093e19f099823d5aa1b7f4e8259d0dde6bab6f093a0c1e5011624a41263ea5519a8760ea2220aa68ed9a9365443d81013c0556dbd4273f8d1a8589bfa92bdceda2522ebbf54e07e96adccd0ab170da2a633b84146684577d331e9664590a6853aecfeb682b3c9f92107bebb47dd8658b5d8f8cf2836f32ef506f1ecda087ec78bfc9772fd49f6ef09ce90e52df6384e15723dd45bd105282fa72d9161cd36c286ab883e7c923420595b7e87983ee40bb9b67c53c3999af53856b427521eb798ec66bbb694cb64f4c2cfc3dcf4797ea84cac08123c6f64fb2b97e75c2cd5e85f03a68d0b41b5f68bcd31d99cce1625277adc92d95fdf2524b12a0011b47c7ffd07a295938d6d4c219817e68d1e116da0bf8ac0a348f9aa01dbd0b8a4825a77b57050e84aa44036346580a54ded07e5a388f3d680be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hda6ed2a37466aa7be3fa93f1f2646c26fbf8fcc2486c472b40a54e5b1a85339acb6c937028e9ee548f08dc9032821cf889a3a4f1ed877c0f80e8ebf6ed81828e36dadf1a7f718ffaca81d3666dfe888659b0a4d45d437d497c71402e5e11716a194343daaf62f5d1b0b2cdb149af67648d16909f0acb506bca7617922bac05921c0e004af53aa11a668e6dcecbeb7674a4da5a6f135ba73633f9b0fb5abbcbd2799b2868aaaf06f44a50dab4f42a752a98754cd8d987bafeeeafed5771b5a1182acf73dea16a22022bef26abd31929816f607105144975604d1aa5ea7da44645bb9a08a952c5e8532c5e6fb6672f54108bb76ace4b9549b6f599c2a6f8b62fb9a2bba4da4f7073bc3be7b02ef4f6398da73160400cc1b354e454bed59962a69a58fe9be50bf551e3e41773f2ca5653855f0ef02a077e7285c1cf96df8a060eb5c7d6a39aeb155f16e45c57eb8c6e01963dc87fb805d17370fd145b2c0ea71cf34691dbc80ebf3401442868566ac83495a4290eaee66f3943f496b169a2fd113affda9968afd8b9c05610a2e9a61b89fe694698aee3d323cbb43dcf0dc3f8349a0c03880a644435e171097c3c91b7350e9d2590d69c8d438ba242f59bbef5c450c441119a38e9a3cd32a4a6cc232eae116d09231934dceb8b9ba040443ac4254218b12f98c273f9338b7752e549db7084248ad4b31ad8e3762f2345cf8ceca79a11fa604fb1302fe8682624e6db4bd65521ea3991cdaf60e555465da9a775f7a6fa3bacd5a82e1bfea22d50e2bb7344330e6da0742586197cbabaa0dda0ac756f0ab223cd1dd74067636e41674d10a92266df6466b10897f58212a0a3a9f45050621e2c3543f323f980593f9ae183c4f29b3c17ec83d42ba8a831338351923c15d348d1b84020a77be23c073e95808a6b528037444b26243e7b849c1740a634fd003228fb08ab8cfba602905eac25eac5481afaf7dd3de70b11a7298d8a2a9c8ee87322cec4b691d4a481c055cbb08d2bc64ba0999659860a6a2530c04f221e74b5bf910d38f6f944d1e6523a0c2f79bdcf85bcbb97bf8e6a24e155c7ca4ebfe070e93a71f7a9db52b9c677e01b826a2e0263ed4466f1f8db7062716e088bb398f8a014a0e351be067f8f32d699f6659607a91455781e9cb4cfa48802819a76350b78541bdc373d5aecfa105362cf2d8da7d6d2ea444e1753b60894bbbd2ee11bf87406b16c8473fc3b14246805eeed57b5e28f5f306cee01fa88a38f641435cb120d77503117ae5db598e273fde2294158e072236827cec63e4ae527894c4ac20d41e4f9e04377759f5f77c1048ec589f155b4aee2e39d1ba8e4ed8e355fdca0150ed4746118a4ad7aca90dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h8ce48ac75561cea08498554a5d398bf3e68684660c6ca3bf6917d180cdc19dc2851e354563d6ceb07be44fd452c46ad1184256a2181f65e6d4aa0fe4369e1366a6b84ead13080ec64779b4b99c93eac535f14f306f77097ca4fc765bc417f54e89cb0735bb2f3a5bc4b5fbe1c1bac60b73d8c8d7a5cb76eef7aba7a60e96f9edd006a3b45e039867408bf3fd3bd2e9aabcab458de32c790a2ba2f8368817f6c2ffcb09a8f477d45a7d354a05dfcb8a9e000aa6cbe43d2041d492adb54cb2f358193fee896430e76d3447a4904b67465d9488817127314d654895024f63ca51951e6e9aadc061ff3f1674270ff9d03d5bc45b61150745971ec87c3e8c122a2ab17610b056363a46a09d356c546e5f1ee36d252d64ee33c83b63ac80f9fe7907d2723002a19155c592e01ba31746e4148af935bccff90d08fd62c6870fe3dc29f25cdd496d5ceb12e590af45058ce91532110a05c74bc5db0b94006ffd91beb1865a97215ae3954c71df5ffa185ba4f57c15b9a5265c6c1f53a0a5e42ab36acba5b5dcec8fa2fc3a3fdbc34b16e72f83b1b900840b90f6e4f58b7439831c3dd8c71753fab3eb5378c202f73816719017f8de4321868006e287026fb1da3dd35941bb1e42b80a733a57e3f2b3a98d4774ec875765aaf44a5553c8769c17f73e2cd115d18e5b564d499583eaf5455dbf2cbacc19e3681f230a0b32c15cd2316f6a6eb49639aa42f10c0b60ab6ddb9b9ea7cc99f07094343f6b3d3989afa996203221600ae5cde5145af3498d3c4855a63d2352a8fd6a7d76ebb8ef34e5247f64fbe2db0cd0569193f756cd0c2d410dfd8f3ff93edabd16783bd0e918b880b860b4389358ce0195688a4969890282704f2a2e7562b39b419c722c60a4f2e1bd8ccd466c81e3f7eb7f8fe8569e5507a84f70929d6fe7efdfd8595ada2f0d93af95b5754b10f9cfdb4b841074ad67a8793b784cca3311d15f1a137e3ac336693a1d2407f6df7141a76b8e9c30867ac8cf1858f4783782bb5dcc6ee10391b4648be1874fd0182d45a6027bf3dc49ef5e62cd33bcb9b718305b20a7ba43f190389c178fcfdc05a61e357cfe712a165419fbc7f8e7dc22dfedf29155bdab737ca1113875696a703b5919f8ef622f048aed0f034f6548b573152e59ae03be44ec3c81de41b4369e4e3ba4e7fc5bbbc0e23f2b50498c34569dc69f76c8b8232685886dca3b193ece5eca7b1a2de66e8f1dab8743aed83bf18221817a3304384f0b5ef2d1fed7fe60c11aaf72eaf4746b1d3c1143f75e6c01d7f75626f7f84ef98f9e1989022fc78178601cb4c5e47d18e59615705199b8bb9e7f2cf0d409821400fad60b172349a64dc464f3fbae079b38a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hb270719e237d2b0a2193595621f1ebb1baea3886c39a77f3d84d9d55367f608883b58f4957d61950efe564f0d5b296a3b2e0e03015e3e4e00b94a552cf0537315d8bbee551334152fa82cea07ad19057c595447c288818d7556d31c73c29776e9ca259dac9caaeccf8d380bbc7a39391b8b9f3083359bb847d5e504dde1dd615a1417f20cf2684018a83dd0370f20c5638aeae8dfc40535961e0eb220b006b972792d45690edd53b9c5e4d3e8714b28e347dd2a9038afa1a51859274959276d62bef34b76e6fd9d7b1f93f1db4636f089fc9f497042718dcd410c76054eabe48e9ab8c307a24ccb459bd6671b55bcfb079ad119a91a85070e41d386acf0f8e823c39e3a8a45c92b043624bba68f49ada1a227636243004963c53afd20f0a1f566bc80e400c983b35ebfd7fc2a6f752ca6060dd349c6069f7075a40e84401f15cf9379ab8267c38226f2fbb7199a00ac9a8395f2e481f436dfd69baf6762889bbcf621b5f21ae020cc20153a05b6971428bdde1a71d766b7bd4be119788d48ca16ad94547fd23f93f11defa13339c7e069801b05cfae059eb260c776d9b3dde1b2a88065e010cca2c5133dd2940638b40a357d7b64a8d1b017c7d1059a2ec06aa6bdc7c6d25294f100698193ac123d3d1d79d6929ab04edb168482ba12fe8e72d0e0918410a1b0a3214cf762a81fe050b2cab3acaa2fe3e7ce564437bbcefeed1abe3ecabe3939d0f673a070962134353bf032539b5eb9bc2f1fa3cc2ff7af8a1aafe7d5ea342eff68b899cf1930b124f93ba0b778923c69904a3ac88e217292adc8655a7c4241d9e6646a623b4c436aa394129295c4c2db6c445537d041cf35683e247d71aaa89f8b6a045a54b3a62f5dcf7c2c5daf1f3adfa7ea3a2d88fb30598a6549d4c63a9c74b40c5661fa4d9dbd770e4756ac74ccfc3e98938c504cb6e4503ba48c86979e557a9eb663243b51dcd506a21f19dc003e69efb4321f7b96adcc8cefc1ae8e877bc0c74c9be391cf3ad409fadc166f7e186efef620edcf4252d3276247f4bcb9c96300b808cc08b7aa61d9b8af31b2554d6bb6a083e0581bde9ec762e71655f16e6a50ed1d5026da4229b2bacbc1c0204994cad404c2d4fab9a0ab9ba109fd7dabd8f35cc7a4940ce491b3d177fd8e3cd217da91bb04a106dca6e07d759a2882aa08ee069cb996ffe3810c5b58c01d6f1a8e61e00f2f6a3014e85b6450151d16bc8e82ac7d42c6cc6a59529ee1afd9a0719a8f4c9665da80eeef81085262ef705113ad52904ef7b5689a76ec512bff738f1548114099155441c16d78aed3fc6271449004238b25ad4780a5b790fc13f80d7fa718af4af5cbc3f546cccbdbaa2e5589a478e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h883e7535e3ce85ee0e3daeae44a1abd640099d4d00b22d65986e96fb02e322c3e80331301144ee6ad2a1fc5bd82bc16dd67d5479beab44c5faa0ded6cbbdb5ca3c322d1a9517bd3c73e12dd359b724e55b369c7dd6cc014aec59857f97dbefe2d8e9a25824b0c526ed97bedd85216860e8e2bf03ece5d1186784aaac189385b2e49ee1dc4bc8ef6d0d088a604d2f9ba0ce0cb6fcc0bb1b4d4c552c5d1d55c96fd6195a6f4d943282636d3479874053b897ecc4127a59e70328a0400be8962c4150d31767139003787c190cc50768008f12664a9276d7827ed39980207fc695b731c931a53cc0347b9a4bcd6831d7ae18d5e4808d193d006c3b1048746bb87d3448196f4f15865e36fc1dd42cd0bd80f5028f8c200f1afc1a58fb50af22e12051d6ea437da6ca779f63c57bb828969f5ebbf4144a6e85be18e4d0d6d6f39f0e7e07cc48ec260cdbd66e272ded379d65ee7d20e05bfea2ff5cb68ea6f90441d7d7acb7b61107cb66aba7d78d9034030aa0cbf77d28a1aa5882b96b8ded8850c10f70bff1e916966ed56745952500b9377468825af717180bc5d307d53567fb9169ad2754d3447ee34c01b6952c46f3b223279df0c12155e2a1513f35d4bbb2600abb00b01dbad80a5515a49bec544d161ad102adcd9bfc3070c3a8fe4f85a21387f159b1d745ed3313310dd0552efe8f4bc3f469886d741a4dc2c79e3d0a7b48f1887e95d61960e663394f6f7b44b1c1449ff8776103c185152fb3bb418b356af3568db4c88fce98ee867cca073b5411bc2d08004cc0b78ed13733894d4c25b61bbc82a402e05d5acf4b38a547b8d970a67ddccafd8599c85f5cf4c02ab1aecd67822318e86aec344411acefcc632543b4c16161cc4926d3ddb011ceddabdb706d300b147acd77a3b00d5bc41fd079bfa9eb215177017d65f34c282470e9217e96ca74f3cf13d1ffa34002a71c186098586efaf3123a5dabde3eb57281f0bb21b82b8d460808079a43d3b1d86d2d0b1674725c5d43572c0ce464296239ccd2662d6e698be510843f4206db8f20ac24d00f809f3e13d21818cebaa34c2eecc0e7a06fabd31c4f08e16fef333c26563bf2630345025d33ad3728a787c845f08094b90da9f50c683c07077c0a4abac94719f6f4ad71e68523821254a11e3da2b27013fc52540de316c627cefa6be9b1cf38fe643cc657dd5659e9a8edc7a05b206bd4c0ed6a573fedef4ab8112707c5f9295299380d77d322d279de73dcd797e9333761dcf67f8b7a6bad4f17e4fdd8667f5cf7962601c3f262870a1b43b1102513404f56b859de6361507f2883612de9c15dc8791daf144b0b23bb413fa7a97102b7531f90545aade2c79519df1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h665a3f8fdb4ce566c36615b145f189a5ca40a58609897f71cdf3ab748cc15ad66895b20f08d6346003122972b4a812682ad34dfafceb91c8a0682de3217bd67cea8fe34a2c7e5eae42b1f0d5c5a4d4e00a8ddfabfa69911cfb668baefaaa3614d52badd9f74638c3e17cc6dcbaeefafe4e079b14a0ec1d9a665b81e0f07d05372bb33b085c4d71d9b41442a56fbb046fddf53dae5d45c0c206dc51d3454145ea6bf1bcc71dba5732b7ab09bde6d4015127edd645d1a005af9224db17f37d3ed732a12b0b6fb2281273c1f76fb9eff8230486791be1c3d28315e34d4603127c8f7b901e850919db02f7ad929e81ea6cbe158b01baefb218843bbd22fd7e5bfb36bf8a673bab3c2a728f4de459948225def11daea4ba377af6d7eaebbaa913d53920296ed90c7f2a03be816bf19edf84ade0740750a8d4e96168d43b28a5ad146a1212252c66fc898defa909d7c44fb426c053a1caadc0d375506fba313a8872606761d6c73fe8d772f8a1507081bfbc4d8559b2f55468da7888107de239d8e011a753d0765c07c79fd3f4d57e2d401041febf49173ee1687bf033f744241bca0c39632b6c3c17f939751f5eda0c49c17c2b3bae54f5951cb16ba67be25b7e51719726b33dc2d00e25fd41c7a3fd003797cdde022fd743cbd53e580e873d68f4233ceb878a1ac2ea27f5035bdff931b516c6daf9188c049a6df8193bfd76c6442a8d90b2339b59b38e76b12d757327350227dd7a85dcb5ad598151804d750a0d605d581d8c24e1f6e390ba5c262a7cb584162bc07ec3d74b7106e8fe0790c3e8e4555d9ac4336f17885dd52463d654acd9727e8d9c2bf7583bd810de2812817c109c5883048663d7e18e8dd9c2131cdc5c2de684006d7c9e77c3a6ab7a519f61972e1fded49d473c81247e6724f101ebfb614a4ffb0eed199c14317d22ae7f4107bbc2070fba4c1802bd6c3f29352cca53a418dc9bd63ebbc8b543f8d7fc72a8f4ea7fecfe4c60cbf62911f8e413ab2240844b81efdeb97ac80c6f5e7edbdbce52a202796c63e227754392d5041ee508f3ad55503bc7ec166dbbd90b68ad617fe09dd6f1bac1898e19d2d85cc188146552ecbc9508dc0663560f202614fb31bc6f9c42a5c5382cfe9594ec21cb88a747aa58ce4a36c8c5dfbdcefb144434f709897236e12d2a8e1c7b5034a1c97b5e1fca5da239efc8360bffaa404da4b4b5517b68172b30467fb5c1f908cf1b3c7f8c843eb8c2089d277c490ee3174f05da232d6db7f65e5af7e243cfa8f2b02825d30e37647aff20c5df014fecd41d4c0e235412c5e35e9a9f497219e52820c6f90d2c674e998a4225ec59152369cc0a9a2207f58806cd9c6c8566d81b8829;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h46493edda1bab07828cea50364442cba4716b16871db8da0038f5b65ce95ee907249054c42eb2e4fb06a1160a0802f820c34e107a9194c265f00a515c97cdb8f38bd0fb6d85e41772d5dd25d9d74eb6f0b644afe5edd4d6bb0088192d6e7489dcfd2e39f0689ecfd987314366e1fa1d53fdbb8afcdab5972c07c453b27384b0ae411a5809e5e1f1efe66370a8b1ddc3056beaf061be453ee9177293fe7b0ae443100efb57308efad83382c347b21c302f333fedb4a04cffeac297bfc2901436ff7904a0005fac565745d1eac4c314b2e7d45e99aa7aa746ac8d436cb6df30e9218b8cd95d7eb4a3a75273d03855d2b3ca850b84622767765868b080dd0f9873b2bac8da6620cdd934031b83f92ff5cb5b7af27a0cb74288840be7ff19ca48fdd2a2b821715a8818ef850a0a1e5805ab7e73b2b452234e2b0a629c5f5d695abba15434f3750efe8d495410cbcf2171f4e24758cf5d797deda1f3a2cad22a686c591599444dff5262adc9b930a23befb2224f82a8f6304537ec2e1e6116183216fb9383de262b5d88ad6653ecf3ce0aed9ad47b7fe4b4158960aec84af779246b5285afa619b222f5ec4870a9f5ec4450d46837d5908337938a6ea6dbd071f3c46f43fbffad664e1300f3c92086d70e45ee3ee055bd8da770b408961e369845f193c04d8776d2e99c8af1d3966ee8928e0325901ee64efb78875bde17533749a89409492fe3f7d3ac38c15f7cd5a587aec1bd81ab900cdc886ace9d17d4f51640321b35bf37f238f40ec7428b5961b34f41b0307175eff682896613e6b9f8492de0f10a3c167b260d9255fb388309deafd9322bc4353a79466595d01e4132d427aa5b4488cfefd17763ef021160e91c6c125442f86c6a4d21c7f038ece2adac689b430f3ce6bcdc3333a39141f6d7796ca973495b0a8476bf3c9d9dc208babd54d5191b2ed495f17b8e95bbc0204833d2abb5d0908f5460896d4718569da11290560e0ee7ff4802142759f3c1948e62f603b10af43ec45ad17fbaaf11c5f0d6aa06947473c4cfbfdd7c9103342db22532aebd46f4658cc2a5c0b74c617cfa8f0f0b2d6822ca8a9d3107ebd07a70ead2c30067433760f7160677b3084a53de3c99c739d28a49b0f4f080e55624adb986322586d00419a5eb195638dc3ed829556dbce63b0c86abe3175f13768b4a493f5ca05075c9c3215d4ed87980191ddc71e92f28d470fd590a79cf9d4115192abfef3fa2accbe722f001837ffe3eb0e64fcde0a7442613d6e75eadc872175ac1b789fd013d12e6e09593520e3f916dd31355c7b8b1e7ab44b94ea458c0e56ff37b01a45dff7dad4608d0ef81c22217de9a37167b775c827ea23f3c663d603;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h532afbf92be632047c876f51d0245951a721d9791e2a1ba06630ef18d1d205d302ca0aba2f2a1b24fdfc3f861ac34fbc2d56d53a79c339426278384720bc943a90b973342a96a62a212f5721b9a24428500b9c6dd2c47aa909da4c7da805adc77969d0de243d5bf15e6105cc530ce72d3b5cae68b5b679ba02a3175277d4cffe797ab38b81b368ca30c3b111d0382cf437d6e64b32757b343b3922f1e6efea61c1467e8171451f4a026d6d7a3a6c38a844a5c5e7c0ec9f15a133682e965f52086bc9582da22e30b08504474e8fb8e4c4b925079ba14776cf916f070721eef2566624087d5fa55bf297b2357e1784d5a9faf9605689169e81075d160ae613dbd5c2d9b00849abe4ed2d3647d0b11f11842592a3476b3e360f005c1f184c5df894f23d863b8921ff23e287ad44d0b3eacd0c6f6cbee1fd69e7f49b22a78121a234246bc4fdcead9475eb41ed26f5064cd7d2931cea4db0167489e200e4b7bd00c34f959efc201e1ac36a16599e66f0b32447f9ff6aab4f9f026ffd83133896f82949d074c954ef20228388ebeeb03273c56482556b4b6ee35fb2830df798089a233f4b99aeaf691a9607fe7c563a655c62316e0b25103b40a2d3c391c8e9c552089184fd91b747891a467eb75c19c26d566c45170d8257a0ebb01aead45475bef913f90895360d348774b4d8cca8a27c2920bc2508565f6de5cd0eb80b6242acc24be343748d32c8e147b9163215b5a697a72a36c2ef6d0183a467dbe8b8492446e79945437989e749abe1a0624479fe106e8279e07357b459bf5cba6be8cc1f7132be930737706531fafae6d31d3d1c23d184b386ae710d2e916ea5dd6bba8b3133768f7760cab6507d183644eb6e24a26bd919b689bed6d11e9dcbb7d00df6d1a425e9dc3d7e7dd6b313cad4225d8ce2d395869ca8a9798a850219e398296d8d1d7fa998e85b7c0dcdac653ad9cbc2c9a0be7f6ef54ad561b0a897f4386f02402e4ffc089922eb420ac7d19ff86756c9be252e2a522f5b1c073e9332583339be4b8b0671060cb79106199af5d6e669d563e8b9fc676baa0303f2bc18a6eb1bfd1ad58d70a316c5cbf9c3aa21f9a9db70ea082831347bfa4e4a244363fff81b7ac92371b27203b3472119339245ff592bb06e5cb43548df82dd86b7ff0e5ee96e2cb807198c62b82ae47fe7e4482c52b0b89fc0377d01f6e6aea205faaecc5e734fc89450e4b76d34e5354db59e26925bcdaa785d677580e03dcd478981c36035daa3a1122af6512219b6f279ef6fd479f3abe0b39ea9fcf7fa7cba8a37f61348812576d043e7efe66eb918976bb316c7e1caab95600a34db33f34cb27957dd9c310c0330a86a922028103e4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h260d88d2bd0d57420975ec513dbdf4963c1f43e3b5c9c9fd1371e1eb1d5f52883975468e619d61b311d6f6bafa0224f7f524eb3b96e1ed5d6b947ca807494d6e0c80ac6066c89e3193ba9837971abf2a93d207170879214d146d25abba5051073ccfa0029390710d1c595e51cd516fec8ab7e8aa9e6649c1d200cbc303e3c28a0fb82de865719d421c4fa5e233b050e54bb6336157578edcf111ec36b5df86060cb09e230f7887b969a08b6e466bcef1bc7e63541e9db61b6a6a518714b908af2e181ffc1ac5a9dbb3548b47f40ac120a1deafb58fd77b1bb7dfa8e066c3676a304ffac457ab0836a3f04eb306ae3507fecb0fc57d601f6ac0b7b757549120325227b964edc8060532c425e64acc44daf0ca75b3f5c85e44e717b9132f4d51c1f6f9612cc526605c5b043bb7e19d9ec9c90e35fcab525adbf3b9a157f853d17b2e1a25e6d0bc604786e877082fd719fae2ecdc14843aff373a507d945714f8c0539b244fab228d024b28feb901490b9d61022b2d1b9ed357d08cc920738c673ca9b52d19f68d81418e81f1cbe9988f4a0ac53445d67a328ffeef63284d38e308afa42d4966cd0bf8d3eec63208642346964832c5ed48e28a0963465a0259078716602bb8260ab47dab65c58933db0bfefdae7098a1356dda9e98f8480afd5ab3dd811129bd649e4b6c5d14eb4271e6c02922bf22d52c53c88d27d434dd288b472707533c1f6fa5e69fbfe02e083883b6b6686f632f891a3eb4a73e1758feaf6c00a3f0ae58ea0e1237c4b32c9e7633c7ef96b9703f4b164eaa11d113792ecad35aaab8316b77daf8ec53aaf9b159cff1a4790c398faec33eba2529ff05f0812f718fe60cbbb7055ea33098c40fb493385150af1709babb3f0de41ac3b8eb0b8900180f2111b47e11d647b4c5b4dc5cc5ca762714dccb5deced59750f488f395f4a7341689a98c629709bfbf0d61f5b454cc3d719c23dd6aa8e0dda232f7344893d26252d87e3309c043e303211549d65c07b369547f5042dd311b6ea3ed1743655351e8ea0c93d5ae9939d9c03db2369630712ba6c90e1f8e9cf439030fed6f6edfd98fe23bb421aba7e6b9e7b12127fe4495f23d56d63fe634ece4913efe063e099044c95f865b5c14ab9716f72d6dc35fecaa9b714cddbf33297936dc742dd7fca913417b1cc3c3289d7c483f7d4411c5c4308f4a32548b0c52d7f501ea1638a3a2bf4fffd5f8145638e3cd2958a7d18a904295ef7c4215906df99f4785d39152e2b504244854312ff94864b47a8e28c21b7069febf4fb6bbf80c25fde8f2a42ad210f02f91f82b909aaa46255b250d4b3e8f3dd809475af6af90297b9e138772d4ce2d68e9269701442e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hf7d69e190d49eb093b8de89238c56354782c2852e8c37755e7bfca267cf7830463ed3f33425002fb2b2c7053089a5b427491da2e8c817389214a733efb5b635df56fa9e71d6eaf5fdc8a0092e62c56cf2f03160c096c4a56874447c8f29eeed1c28a65dda07295e5590d83dad6eb307d3419e80ba04dce545a02cafc0e60a40d52b1695ac4fc58dc57291584d4f743c55cbcae17049aac6c03a5ae2aba6e2644452e097c6fa3de9d556cb3fe47543dccd9533fcd62c51aa72911535e0912a93912043daab8998ea96913c1d3b63d3e0711586f69bebcca69bdf1ec904be470b036730e0e6dd112d9d99f504e49fd7d1187cb489459165f979c83ec7d5987d840e17c069c1df21b32ac98d72650e75b41da6a7b925d8f747f8f77265b755e28c6327a1b786144c55de2742458cc19a6f424cc110200a5161fecaba64beabf6b3576d76243159b83da31806a123ced75594e9cbeeea1d829ac4bda05571c08ca606325d3b996e30b3e21aa31708e6271e4d07fd8a92a7dd74cde21df695fb2ed1fe50fd436aab4abc1623f03e1ec3f55289cdc9bed425f31425e0e1edf14ef12d56db89286e54b728223f9ffa99860c0ce5d457af64ae212fbf63374fefa45d80a5759e95510bf5a4de0bd39a62fa515c13cfd39c9a7013312b2a0a983d2142a2b51975a3bb5ce5a56e25181efe86b84f9a64bdd6cba32fd571c6068397ebff7a888954fadaf0edd79ecd4cbed0e77de05303bfc94d3af2bed521ed27ff5f6a64f8583658c75d894d3b9b0fb3bd9e59f5ee55b0a214c314924d3a94e6df4facacae666b266ed45e1f1b3d8c180adce3283b0675b3c4af57cfedbfbf21cab4d03100f2c24fd5140f554828f2bf45322eaa778bdc7228ee036963c5250454cc4f0f2b4f3887c08c79246dd08b9a7c44c9f012e591b4630e4d54aeb66c0a5447696cea49bc1c98354525ae3b585eba20990d49bf90ee9142859e64d808cb92082e943b84eb7255415afc79686b2fe53ffd7c46a99022ef57b3c907091d8c1d27e38dc9c3a68592c06d170d2a58c78b1e80053782a9a07b736a05e39990ff49c01e61f229886d6c504a1d115cf8c486e7947d2b1333e0368241542fffd224d30f55505cb9f61c3d7f2b6ee0aabaa94676c887e59c1c8a8363db26bf43cdb49b8ba87e6b2192bb63a956ab34f48ed8594b2f36e7d554a06f4891ee82f033c2e3afa287b2aa8ea6cf9f17d6354e1702090feaedf2ac0cc7910641ff572a94be9cded8107b40d4bae5e103adb5c59931832f53f7b0f2989ca79236c6c55fc4c9e34638d46cf1a5f83ad10f882874c9a341e5cb737ec9d0e9c62a74f0741dbc92d6b9bdc13df0a7d587e06db34943559c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hc100b1975603b6f32c9b31dde7f658d2d321f27222fab4781120a75a14c08bd4a3df160780a0b7ec4a82d4fd23cebe3f48bd0b91239939fd7fc786bb0ef779f53fedcf6dd8fa512596e3c1b3a13d963a261a39c99d69e92b0ba8676778ac58f6f4f1aa5502ba4935270aeeda41352a36239015f949954aa20894072a21773514460451fd2ef34bfa1b7bdf5dfa9d5a350fc9eb574ec2c4280bcc45e52a40f859743fc8da600d9407a59d9065cd10064aec6f3e44a9539995ae8b330d30e318d350fdbba2fad6432b91074a5fa8eb50c1c668462420e908ffb2ddc993c1b87a9c3b837b1ba247746fb5d1707bebd3de9154a4e6e4657b8f9fa1d55d38ca72244bdc614a291a956c72138a418106db233920363d05f66a40ceff4baf9b229feb24f6334f5afcd29f0cc907ab04013f071c568bad92c9a05cc110520cbf863feebcd621f81b3430bebbdece530b338a66502cbbaf3a6af9233e8271cf4e0872177687230d8a353b29656932f929bfbfd7760ddbb21421bddbd92ff0940a5ec76e864adf1a0392277fe4e4e87d18cbca7a3a49c4ac317285df8edbb2d6b547eb5b372106c781142cdbe6f5e3e5d2508b3b4ee4f37f6c0604f66ebc29f3e773f650247a29539c7883074dd9fc64cf27bd998216a8efd7cb338b1230a4c942d44bf53bfd15cd2d0867084f5bf1577c29762c6fca09bf1ea245aa3bb8f5acb067e172f6cd91259637a70c9d7ec362de1c0dd406bc61561ae9d51f88c7ed6a9f7b02d2882744c241bce3e9b062e85034e66ba2d515e9f25c7b79e98af9006048c3243c714eddcb4dd02694977093cc433b1f45c047c45104b0a11a93d959cc1d6712318cf194908e570f5f816ccd8c8133f1611a52a896cb775d4f4658f06cc973fda1f68656fd748c8248b6d296b1833575f1cc080d9aec46dfc6217269f0147e4122f27abf4f4896ed40b0c750bfb2959325d48818cc485e84237322ece71653e1bdee9e3edf242dc8d3e3afe29def12e2315398383d1d0f50e35ecc1e7c01a7a44027df2a92601a1f10fac5868f2212c5a37e2fbc6f8770178b2179bc31a5826d2939cd7b5a3feb53f30c91c9d83c9dc284615bbddf0b6a6da0df065aed73cdc1679191878c27985e6e4360b299bc14df9dd9771a4be9bb604182e7dd4aa8b0f1dc61103d6ffd481b8a935d329e1e54ccac2aad47014d09ac1353f00e2fa743b87bc80d243a85d772ed8ee0d1e5396479faf5ec1ff7977f05d1e113c1acf8aa5c5a399b80f33bd73cb1f15dc47b91e11644b2a20c877ad66c0b7479133545fe4132ce82bcd86312a59b3c9600c626635bbd23cbac23ebb8982129c2f9c28d12df705349f4d835f98dc203baa88ad9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'h30209234275e53f767ef48584acf00e93b9e5aee1f52b3eeb0c06794e8a4b830248081609c22a39a5683ac5e109c1d62f74083c996717e753eb860a8b06f5a73d69e59796dd3c4b86c055cb9c103fad0da8c117b1e5c4ceb6e5c310f9c100ab7bd6d55d7779974ffdf3e55f087926cc2dd8ed22691ad81bdaf12dfefc9c3cb04f99f864f97ecdd933dbe85baf7cd93b209c9a0e5c82666c49d56fe522ff1a094609283c1d839a07c7aeabac0fa2b32b44a26a5af86ee90e21cd1ae947ecde18e6c0dc5e2f1de2e60a65638ab1cb0c3ce80e4afb60af25c161d000798ddeb416c69b2b8a390ca7f96e9040f44a213ec92323f86a705b8699f7413d9a04b943d5a4b87e69682a36fa75954bb8ba0224ac006c3af908c195a9d8dec854c9fb2a06b2b7764cb4083aa432058e363af8de94eff72a018c7421c7492d086597d3a5d3d6b31db7075ebf4e185288fd26c717dba3ca1859ed6d9a6d3adfcf79404c09f512adbf842e404f1c1758dde340ed58c3e3b3ce1ff2caaa353e9a8e4d1449e6d3c3d74c088e227f278766e6306fb235e43b3bc360de6994baf85d40febf6ed9f4d7722f698a840079f0fad48dae40a540380c258a0497ec29c633957382679606e9b902b269c7bb0d8690567e20535da34c10752ef4b001c29a46c23de3f175272b135567bc4e08941004f23cceeb734283b9f7f9cfd0eabfaa9b70bca99ed65f3e2e00017abbffb8148ebee3e98fec8d747e3fa9c8ceea7d7efcbf0986d54d6149a52b1a868ad2c8080c2094a419b5e87deec3979f80970547d0f8f2fcfc9a90e2c3b6e44aa6c98e6d5214cb1583f9fd84ecbbc069c42715572184288155457324c4a9d66cc2e3b37752fbb5449cdcf7ae58ab1e40fa1e2734579693fcffe5abe184ca97331eae7e1b4b9cd0e5a89618e220f1d2072a967bde1c3f52549e8ead6846bef4d5e241e998764b24b2072009335fcbf92b2a7f437ca71d63fcd5afd815c93b9590d81bb01a2a4ea6d845f8493e48d6c3b9e80e0cfab5e65c2413b62b2ac4139ececd524cd4c856fed341dd4b4b5ce76fda0001c37ecc23dd671f4f40992d32565898e74167b738511e24d224dc54b137bea55b192118612c7faec3b444d63aeb134a51d3c08cbc7de15aaa568b6eb3713526bae48590367951d0b2c34d9882c564f24dcd230faa22e784048d76f2fd179a1c01f8d815b23f785aa71e23bae3f6524fedf122e638e69de4cc1cb21ef775d672850f5623da1a39051f4e3a40bcf92fe8bfa207ffc6061f835a12810a11037bc08733394edfd43178039f359224609785525ec7294f776aa70a42602d69c188ebc8a48ee0f09fdf386274967c390cba51f14e9055aadcf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hcb2978c92cf20f95c24faa9b65dedf3cd1f11163ca6c822eaa46ada9baee54a2fa842e2d8af5dc03cf6bb7d2c0723c7b4b84699eeca0b86100869f697f1b42304fdc8144126bacc1440d69c521a845fcb675c3b1a8d5504d80c3645e8379fc75bfdcaf13b96e04dfdf6c20f942bae1da4a962f2209f8f16c1e28b8c06ba024c2db3970b5da3915ea56bc85ae0e72141da407da7c7ca38237f8f90fc1cca8d089b0f53508bc012ceabccb353217485420b5972c4a56621859dc2446d04d645178f8f7028227180de123fbb3a62d8c898c1001685b747a3791d6ae430f666593b67ef4628917ddb8ae20e2105be159a5e150fc656d2aa169a60d02fe4668e018b1a8dde720fd4905f5f0951312d50d35ead9b283d9b9ae52509e73939f1db83c9b8127835963765ffe49c6936068529acbeab39e9b7b2feee4c6a98889bd614efa738d077c21333d060a648ec4b04444dd0d8959b859b7042213e415b791b659352041e455e0a0815120d8348863d1d015cac56406be467c84b411357a222ad4dbc7ac7a1de50a728ea52a71678167e39f1e794e5b59314feeb9c09a62e8f4fd40145f12f06d75f019a2978fc9e3539f2416697c693dab2e1e928f1da2572b6a2d9ef929c42e16804dc15d062710d5a764e512f1fdae0061e478a933b76cbd6d2a119267308f27df850314ae11b46e4a87d4d3e0f7a4ab8495e7f7a97652667b81097424ade82ba00446e42a782db7b8a1514af545af39cfa47b46529330d9794478a08807c673585fec341bb271bc27fae4252d23124abaa85fdfecd36505308101eaae9d031c27ce244ff4fbbb75da565c0cc18130051c69efa2c93bb9846b7c7327c3870afeae0d223968dea89e00632260caccbc6c71d34fbb2fe886c1befe49e903c77f6b8d713bc5b7e07f4f730ac85ec502b21b35fcd5f8b977bf31fb9d01ab8f2927340b2f94ff7ce682f68c32c9c0edac1a0c670d8b162db0349e1dcee4dd91d7e0e3c4cd6ce598cf8ef9bf8d0a47529fb8a6ff386e5cd83f46b1379d6f1c29f4cc8d8a22ba01a79a848875e2f03881a6c1755544b10bbf7e2e58ebf622b3c25d10e341cfb132cc21eb5173e1159d817889d18d71bc1127489d9fae4db404d23367bdd70b778077b45f0b7f7be1b8191ed019599e76776cb49dd33b2583352afa67b63daba953ffd3f0f361156230f8b7b1bf75736c2c819d3631b8f5dd8beeccb172ddb6037d3e862d2d8ce5bc5d588ed4516e15653c3ccde2a110712ff1285b82531e4d703a0b14af3ea265e8e9ed4428710381d171ba2a42195fe011ff56623182ecba8ec0889f6be82f41ab3836558e60c3ee324b3500e5c3066d5acdfa698426a4236cdbbd0e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 7776'hd289876360b2deb06810d8b87f576a31b0568d31313c881758e787a3867eca2d28c56032557cd906e7a82c90a6784229f6947c1a933f98482526bb8a2d509c1494d801410e1dcda697f4e68cb2daa80329564b8147fd776621da550115594c8f9a7e6391a7885616f56122c89e5ca4743173117c152cb6ada403473ec71be2ee132f75f4d48e6db8661cf1bf3638396b1ffb1819fb2438c0178b55c94b2e71f2ce05cebe27505d0ed18b565d69ab678215170d40c9903d9c35b93994ec80aa628a28485b9835c8b89aa79ca7b078ee53a7fbf44efad350858582ee1931ced9414aa05006989d532153f4d71b2a6722d67e7e41237eeb04eb9088b81e1867bcf270290b43163b3034265bcf4f132d393b82b9cddb3705a7fbb9a7a49574b1bd086b8ea249df1d7860efcf319985596ab7d5a9efc86b0f97854ad33edd3f2a89d65cfb1dd80c882abfa6efdba8bfbdf8ebe3c3e917934e6185679c9fc8673d4959c33ea7d2685c381bcc6b6ed739cf889b6afaa6aef6bb259132cd2a7f8ea414946f99444e7e93a3e778386c3c6550f5c0912913320382da7ecb2a8cf481c01c2b2db009dd17927298883129ff8c5e40cdb36e03666e6dda7beb7b4cdb4e813e86a716bd70b474b9e6cfd0fbecf0f6fd8b499661a6fb8cf64fff6bd5f8245e1c7a08a9b8b589569bb79e77396df8073a270763d0557cc9652e0b5e680cfa361d19b02492a67d14a39a4a27e1ffc1dae2031d242b48d810b7b229ca90da3364e8d2a630e5d3726ba9654c339d6237e224b0f338fae8d921e2d62867c3921f381226c52d6c7a7f4238e24281b188d033d7c78c651d61e21718690f4130032b40dd66f19417c174529928b3b069c333d145d2796a22d8a6ae1ff879708cad00ae6b595f82b19824d3a1d42818ff93cb642e14a1cab73b791c8862b55caca40aa65ef1be708d0a910de350b18b7da160266642caa497bbead1ea52c9f6aaf2fad1f494a9ef6118912aeae7ed8e848c6646de5b00576ecfd73a705053a8e861d86467a3ace6177eef1e5f2f91b18c152409cda49c38433127ca8eb99827f78a519c685e1ccf8d092bd24acfb5be6168a141dd13eb3404c78fafb79f86aea4da536896502099a912f623e16a1c66d664b41412cbfd09714fd09dbb25066f48f3958b8c501e39576be51fc647003809f446301667d3729112e72d4935f192c46649c9d3e69410faeed35c06e424456a1ded738b7341866569910a735332fddb4414105775e467b4b413c8435be68bd799354eccf6331067bf1a6283717f6ef3f2b679a66ecf5e95650a1fca1ddb71812a6c47fc5b53fb5294c54e535d7f7ff5e9c8f2e8bc45c3a394abbba5fb48b55782;
        #1
        $finish();
    end
endmodule
