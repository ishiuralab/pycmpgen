module testbench();
    reg [14:0] src0;
    reg [14:0] src1;
    reg [14:0] src2;
    reg [14:0] src3;
    reg [14:0] src4;
    reg [14:0] src5;
    reg [14:0] src6;
    reg [14:0] src7;
    reg [14:0] src8;
    reg [14:0] src9;
    reg [14:0] src10;
    reg [14:0] src11;
    reg [14:0] src12;
    reg [14:0] src13;
    reg [14:0] src14;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [18:0] srcsum;
    wire [18:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h51a2554b0018cd31d7202b5a22fc1f6b8ce776ed4f7eed38b6438b79;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb73e01405af17d4b5d744656c83d6083ca1878f76c35ea6726014706;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h138c179b24bcf0873ba68754016c03663c87c04463725e5c8df149fa3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9f728ed888420f4f72ff9478ffb6febbb946a5eb18684162fdf3a34f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d7a6ed611d5977d561acf0161112d508158a356192784962081fed1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h410aed329dd973e05cbe5343d1f2a97b222f2fcb2b8905b4b6cc8158;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13c0db122100b15726aa4cc177728c8b03db3f3d141b79905689f5399;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc1cebb4b6065ceb7a44ff4e09050b07460cd97d2d0777039e5887311;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18bbbf47b0d4d9b91b0aa542f8363cf66b9d2b495537beab8239950fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d7fb85804c7d47ac2d20dec6c52bd78ea76f915e8def884b965a09bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h181353c1c2edf0600aeaac7e1d200ad1a459cd51a87063f76b266165f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h39f4f8baa1722d55a1255121bc3c2f2ea57e92633f44906877936c78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17a2392dd52e5b5ef67dfe6eacbbdf5f6c067361c036e80812a8c1a82;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h467efa5727c0476b7ac40bbff9c49dbf0ab59af3e0cbbc2d6d3b0976;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h170d9ce7df4f81765b35e954cf82ed66bf2ddeaf2878d91af2d44683f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1737a21040d369359df93810be06579edaed4a6ac4ee2dc638f5fe9ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a1cf20344327a8c9862dda9a3b6317f822520b5545718373d5db3a7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5f076a070e1f71c1579938c5199deb81d1cf5f88945c3f7557ae63a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h65dec348cffd8e7e190560586863e622b58db7049d6a2d22e0a0e03b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1453d1478fb4b371abb6e408a013ceb36c8bed09791e4f4a9dc61288d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heb4542d7cbda71e1bd8f79b6da692aeec5bf74353a501291138b8591;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13c76f8298e33077298ad50176a09b61c8f795d60832c0e33855f53b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4e1d40a96fe8915bf1a77bbffdb5ac27553f31f1187c61af35a4d8a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1708cd28b6aee334901e9ec7f83851b6ef7b5e70d12a803a06e2bb03a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2d2351f11596b88000935d1eee1e1c17ee8d64d0816edbe9a9e1834;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1204294c286fe69b2154bdeeaeab9ddf7ee0e27315b2fd3bca3440cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b3cbae5cb71bd04b41e4252c75ec5f0f1fbef0938169d707e05e0640;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10bb4cc9e7bc9f0533332f0a95bf9c7b5df2fe110471e5681fe6c3145;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h41b31fb3e3aa545d7c841f6d292fd1083725628c82b49cef5a7f4bb9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha12d248994876daa90505cf9e49fab446d31bf6c71dbf983bd08030e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13db7860296c923469cad414d39a4766fac0cb151fb5310d1805bd6a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5c53c7da3fbc61cccdb52afde1fd0a852964f034daa958472dc10cce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h65fbf3c5b4a00b6d50d66faf3de54ab74d50ac5507a49da6b1c6ffe0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'had0f8fe00c5abe38897de407f112d450ba2c29b810d65dd1ec6929ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h65dd27d9b9bb3870c3c507267009c4ab13b2118692976db84b7d33d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h64b097180bab1150e9fdf94f40eea731d3a5e5ac3550c3c29019fd49;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13159dbf192e7e26023e72cfd0989af7a50b585de4eda170aed97db6b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3395c94528bbdb1633a7dcee6b251bc0ca0649418f6a57518a28e8fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1972c6a02aca5c98c36ae0cfa8cbad920f35402bf8382f7159f87e958;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf516fc5939611aadf8a13bc9b0fbd2b21788650f6c2c06dc18918a5b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h424d6da3dcfc6d5af8fa145c16d3880b54b84190170f266d13379806;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16ad2225d168f80c678aab3e1b97502f2dffe556124cdbac5db005ece;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hde64abea5e169855f33aa4ed77ef3ee706b298eda3f08026340c07ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aca118c2dd9beb7d52dd9e6b667573fd31f133d6aac439df79a07729;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1277e16c23b7ea2a94093c118d72c21e3703ddd13ca2df524a4c8f6ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f4839bf09e19911b23d7566d9f374665aa84610062749e2177d149c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h153b3b5f2781a79dae70977f7b8583dc75c2c65663633742df00b18b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5d5d6741a6e6aa1de03f88dd018ad4f3256412e8dc5548a1a4303a7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a3d20af3e9736ae011e4ad88ea56bf9173a016057367746b28a8634;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ecac7f5c611cfe47721705fae9a254e3060ba407f98f8731685f53c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h170fbcff17c020a09ded1a37d488b5ce86e8793d03db8f4334c6884e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9ff095965b40059cd244a37a258934e4d4ad4f08ec864ae52d9aef34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h456d12c5d288b5ec80b4bad2a18f246d5705dc7cb8cbe968e070c25f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12e58e674bca903589b1d3438604d6f7cff9cca191562c3e843cff71f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd2bc738f530a797b589150207c7620530d448f92c2ebd4f31a1643fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b21f2fbcb9e68d2a0a708beb57a2c9619adbf9b2ae5bb10895a0105f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b928ba14da2c382308c15ce55ed790afac22cd4c0675a476eba6e75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h152211e18c17c86f1cced1b731a6cbf19fdd80881423a48056dd69c7f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ce363e20fbe6abede5dc0b861c6e5ecfc210391ba6a932e5e92c8c30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d8066be72f2dc38733475426131d40d6f9f5f009ab855d27d71f06c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd2ba219e558c8322a3144947b2fb457c980b1979147f5b2cb9d8e439;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ce24b571f75e1dd33f76c368c1a79197664f27fc7728a1400e050014;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ddaf620c2b75b9835efe4f380dcc9d483ba8555293c64638068d694d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ca1b787194d800f2a7f5f345b5715f95911dfbbed60b24a61d16bbf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef1aba95e2ca4dde0cd5cdb1564589a9a5f6d03bdf6a22f7c1a5be88;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h505d56e886b0b8119d509690f10115c9eaa82ea65a4cad0c16ffed60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1935c7fd52e48cea960796e0f51970413f3776a9e75269e070642300f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h110c254601a9154698c7ca5da7957ffd0b32fa96e317ecb03f08976f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdd58782016a91f98ea12f8dc4e711b074aeac0ecb9fb6f675027c2bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h874c144d7ca44a0d8577dac548f2bf8b7b9d78f3455e6d8aab517dd9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e84022f2c67c87b6358240ff2499c23c8fb57f23ccefd437e3efb313;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h255486b67ab0828916afd5fde1eba0b3c25f1594e3afea8bd3426d12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6c768d332f02a254e8d7e16beba969d9f99512406df9741dad43e16;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h185aaca7b9b387694f17e6a80e2720eb02267bd19f984403198efb163;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ce5fd7a771bdf75e66dcf884004182dcbcc312be09eceb547f82e571;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f9f46936655b32605719859058422a62fc27db327af7dca0767bec1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h41ebd89041127a453db99aae973488d4cd53d150f638652b7fb8688e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18fa27ff8a677f229140e466bd02ca3eabc4299c1265a48904c9e11b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h35e0300143419c106a234b4d42e0a36b3921aecd2e96e6421622ea52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h126f5d9df99dd43cb0750ef48d25d472017534add9a51ce51d7a13c13;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1585c022eb5ff59483ddf2c6a99ccfcf425fc7252ae4438fe41cc8ab9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h167a023f1d38eafc59682423043b4df5afc2e8c180462dd2ccff91286;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c218dd007d70db0cf8700a394344fc771042b4b7909e88dc69ea4928;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h30e4a9bcc5e03e5684d36a27f1ff7b25df93cc4e2041ab0a7619ad60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h132f8ee04a4b077b049ab91266c6883acf088f2e6f9de2aecd68088e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h33769c29bf415c1ddd2cf676803acb218760b87d533791667e0469dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4f9546d0be1758b82f940d82193e412c64c85c5002f2892867a1f1cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15968335c1502e60987bf8d58b01b0270df463180eab80ea79b8931bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7e96aff93ac650d9dfc9434c95f6afb37651cac2b30912402869e6cf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dfec3ff5a45b0999dab3db5b7864031b56dc62dd67e3439539b9e742;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf29a256053a4ba8b0e663dc1899426233576b8d76ea4010756d6cf01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16615976033a20ca678be7294a788ec702cfeb220ec751e73c2be06c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h53c8a594d529a5f1dbc2a08bd789816a0d6c0ae7dacdcd31c5e6e619;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d6c2089dec60197f7d5f481f095604c36b9876bf0a1dc786afb2afc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h51f0ab3f79ad011efeb0ca67e844aa4b52ac0d26b950676a6eded17d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19439cc4991e636869d0c6442dfa0b173957b51e09562efd87ada1f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h175ef6ce9c496b2d6162f0c2fae966f2d93f78c719ea6fcea256da0e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cbaac9647479da0a1d432d02a5e6c1bdb0eafff4403ed8cd5e2d7497;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h62d66f8c3e4b0cc7d3edcf8c8a836a6f87294cd4bcdd29466225fb94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2cc5edd2b8e56d2dacb4b24e9f3b559c6641ec6c739f98c24368fec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d4c3eec0ce67ed464fcfad06effc72ab838c1b489f65095193f26c80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfa5ffc8e6b0279470875b2abfc29c80455f2a7ae6b7cfd62e8ffc9c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d82f50cb3a82ef3d6d90a6af7535eef638dd486ef97688298a7a381b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee20e69b8d106def99b9e0f86bfd248b5bbf6a31d48cf35365282de1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6ba86e62795c59b0567a0e56b646ccd9277945ae6dfd222256d28087;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19585607db8afdd3933c5b87654ab4a9632468c41ef2e4c5e17c9062e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f7da088e2ae06ec69ec927304ac10ffcb05835592cf96146306adcbd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf33317edbd17e64240805a7233d66b13f8d5c60bbe719be0d4e7f61;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bccc05f5ec85989e86fc9ccd2a83547f6db56524b95a96d63c893d15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ab85e201da882d0dd459b31112f03c2304eb498a7830d426bdf15a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16fccc0832d54fbe029fc52698cbf52a90eb083a4c5c2061646798fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h80778e3ba127893ae90984595cc0a9cd404138bd619d925108fb5159;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h782d61a6cbcad65c968ef3af5ea2fbd572531c4e3e337a44a372d288;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16ae86503ec52afe8560824e9bdcb69090f4161a9fef4b05ee101074;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11c083722af3797bbab77ceecee64739c50d8ca51425899078543c319;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5b2f117003f6997e2984740430f5e39bbda04fe3decec64ddd652198;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h49bc7657ee6726a5f414536aab93edca44cc6971623fd10294dc82fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdaffba80191f73256987c9517d73445e7a7a5eec48a851a1f83a2fc8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1725fd7ef2e6075341266bd81133fb4378be2e5d80a1245f68673db7d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h995257c27108e787bfd03580c9725ecdc3e8ebe7cc9a426bffc87c8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf5e4360318b422fe10e21ab03a43f2e46c98f7e6de8e513a1949655;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h829cf87ace749511781cfe4975b3ea7e49a33eb889889f3853a8ded7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcce683b1da6e73bca299f2df2736d63590a6a14966c34429e58f29d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f9f74cccf469a852af545285567e7dad6c7340be33c61d1ee1aeaa04;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc2f14dacab850975eb25880733fdae6ec58de4544c59766bf92785b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h91819bdcb1310d5250fdb21871bbb4a8155c3b0ddaeb12d5657e93c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d042f5e41e0a5e6ba0473579d25d72d0b9e5a4072a1be97005d9704f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdc90fd6425ffc1a64fb8d3292950f4e6eae9d63cc551bb36193fa6a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1237e451597719a939488870435e426ca7e4021ffbd6e6c9d7fa5d415;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13c2089803b2c9df5c208b75a324ae7ad060d9c8489a53ced631208ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10cf9b0b13c96bb489a519ec70d972647e2c5e764efa767abf864169f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b966192690031d7562686e65b1356ded9a7407e0ac6d5deac638f08d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff137bada4c60343beeeab1a92332fd3b7f074e7d64451718ad56faf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd94cdc4ffb8e9bf1b3ca6afcbdceed598f75f4fafa9adb6eed2c6fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1494ec909924eb66cb38026b8cd73182397c43a9da6ced7e3017daa71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3fb0b2cc07a353fb3107fb14669bd7f064b3a476b4c272d65dfa423;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17a7ad461e493bcec73a333f134c5952c269fb1138cf945aa8fd099a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15a2f9c6c3d7957929e7d6969cdc7bf59fc0d0f74fc904cdefdb99322;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc74750d48700d2068c92c451c50b9abe8d5c74121d1b716a78292b71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf8eb4f39a9ea3acd1445424c8aadc49a605e0ac05f09ba5009aac0d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16abff6ac1c620dc91997c726ce868f8d0885d034b58c92f0af24c23a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1484ae8be5463c56737509f572257bb572b431257dd1b4de897d4bba8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ecb6cf5d27f7f93c65c7e0d0c45010519347a3e6b5fef4ecf4d7303d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h29160cab7e08f1eceb74e0f80372d1abc4007841cc25f652894741c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12b7bebe5883889be08e41ee5cb0f2cfa09215cb20d84f98d9500bbe7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'haa6f7b4d9f4e3d4a72df30f63303d19dbe40d9a154bd3e9aab36bca0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a471d79dc021c349200a8ad703ece8e6d9f14a37621ee6be70c7df3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19187d3c04c9b7e93f6c8c45115733a33d99eba5481370e840bf3cd0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h311fa158da429ff9215e34db1b7e909cd431e7ffe7b1c7bddfb02139;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15494a5607e9cc3fcc8efb2cc4deba0e4e40d10ab1bf9a9cc8a6cceee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h64dcf6374628eb6bcc909c900017617d3b61af865b94c2f08d0e730;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h48ef57906fba09d2ffed5a68c1ccebf007960144f97f6b68f97c89a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2492092bd2bf8992f7ee225cb33eebebf4e74cf68857762e13e894ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2f525c880fee14ce0ee26a89c231a03808ae366e5e906af95077b034;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16defd719597f2d93a623455feb755aeedb0184a4f8ec99615a926098;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha930455182f11be4e53718348c22d75377a7607c18625ef65a4c03ef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e1e4fdf779a3c69ae8405c2eb0c0daed92dc643296f0ee60729fc75c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc65bc81ea2aa2a5d23379330ae6aa4d6ed2357abacb7d1f07be677ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1971ea733c2c6f82495be88cdad728a07d4b0e6c252b4684a119126c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5873ba64a039ea551b6f5591f0dab1e0598ef2118bea491cfa5d662e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h72a3df96cb1b4ccda96156898781db59b5a00ef3f1dc25d7a43a0ce8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hba344b13de88b2c6482d6c67da6fb2b3a6bef74d9b238ed10ece73d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h23a8dc0c65332060338c2b57ebffaae039d0da3e239ff46b674afe5b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a6a39c448b0f174cb0b3c1fa7b6ec9a7978c82c61791f4d565df4d7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h181e09c127f3cebcb369df4733403d16fffd3765b2b7bee28e6da57d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9473726439a4a407ace757286f8efafaa9980d6d0d190260b6af3d88;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3387c442f173e4a9cb9b74926157a15900bac712568d4726bdc360a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dfdb4809ca6e7cdf583a0ca2fb6cb377d8da89e63f8a335113783465;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb25ca8da7541af2f4ea2939088736f39f011f4d8095c0d0ae5bda7c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3409e7b6765e7605f36340dd8697bf5ff0dcfb388897d0df3036025;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15e30e6126f7241114950bad43fb4983d829e15c6d0ca46166ef22b0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3a54b09710a907fff5309b6be19db9d677a8bb0e9830402c0bde2db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17d9e6ae27073c36f4856648004636b3f56109b43e5054240827c0d91;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcc4490862fca806b98f2a7201ef5d84f6df30421575e093770491ee3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha1ded01bb4986d73177ba907c9141395dbbed11c44aa518543ce0f7f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha69311b143524cac8c544d93b05a56d1ef1d83ee3f19a698adccd856;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13776cde0086f658a9505c920335fea82734705446297d13e4d132713;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2ff5de34e48142b2f790b14e0c7954483ade344f490e5216b78fb77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15d40108de2d40e64d09af77cd4b4182863d5d29811c6af4fc3b35956;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13d796338248298ef848098faa54c933618789d042b9fcc9974054c28;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4de7999d1701b8a87147e5d763ca63cf8dec50ca89b62f3be0a482e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13bc8461cf2308baa04e771d03f275f83cba09f0ab90cd71eb0683b93;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h179551f0d49ab8826b536262015af46d74a30219f5942d0d9501e7240;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he7671da789c60c62ac9901a9d1cdcbcc8c0126ad40db206ddace9af3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd54f8c0cc7723014e4b63ba6f220e9e4b467ab9f1fceab801a242335;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h758b2ee13c01e6c21b4a662a24514c6ce00b6655eb08ab1f5f8993d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h45d5a07e4942f574d50cc577a7626b6d797bd5c05d468a91ac92ae91;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18cc69505480034b0a5e93d0c6684277dd7dc03fd5719e1bc36a7ec3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c9f2a3022366c1f3a2d153734459937ac28a042f123f8198c1a0f276;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf4f8625452b81b728c68b330aba2fd1c5249958a96b459884f8f1855;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17c72b0d8c9f76e91e33905f476fafb6a6de98af4d472e809502e592f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbdca611269cd7c50efb99df71df8fbf30defe10b7aaa3d3eb167003a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1416a1c3b8937275cbefe118b9d9668c36d124b274f3b7c05f3dabb84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha490c20cd5aef985f59cefd0109512734748db3619daff52dd444aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8037ae82321a02db12fdbca35dad4b38f64415e61ae23a2ebb9e0552;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d95959fa6a2e501d8e3fceb9c1c7fe1acee83261b447c15e4ed34603;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9f091893dbbb7c010874808357c150340ab3538c643f85275655121d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h30a0249f688cda2cac571bd5a6b0d1e35477d471b6b623d66a7c7dfc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfa5db7104371e58f51c5a8f4a82479d484671d9ed260b73323b40aca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ad7c4048d06100077bf57877dc74eb702127d11103e7a30b21ba079;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd2c2097549fbe0666425ac8f0e09700cecd09dfa2d060af9c62026e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h28d7ae87d0ff6eb1d4dfe0e2bd16890eaceca6f0d3f3d3c64f6829a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc086f2e7ae8362be7fb65fee98a28c97af65930a91b202abbf0503b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c7a9e5cc611137aec6e22cc2d7f443183da063acb17e4d8ee33ac75d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5dd4f576d658fcabfed993ab49ba8571f1903115b3c5afaba055425;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13cb78044e441178ed3e0044bfe1049c19946a8d846959cfd85d2207a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h193223c80c026b17123df9bf8de851b953644f17e64e379cf8785b833;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h40f5c5d6dcd2faf4f2c472e60cf73015ca0f7b68e76d766dc7e5b6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc45c7d2efe6fe38988db32eb1cfbea85a6f5f8e587fc49bca59be75b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8f89219b5b2620592b0f51a94f204ef7b34da66986b6a12942d668cf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9729f9ce7be7b3960941caf3be4606c74a8418cd369bbc31d836d152;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9100bdfd2e784d6b8e65c2bcc9f46aa7d8d33470bc7cace5c2a3152d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb31ed9457b7da1bf58b94fe4b6051a8ba92edc33d33424d68e354ae7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4b402e658dac0628fb587b3ef354ad84d15f0e78670e52656797aebe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dd52448b2158d9b5312f51c8a001d18ded73a16fb0cd708101f5c093;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h168b77a8d1502b2e60719629aa69b8f78a36a0837f6873bce297146df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10f65862a8281112899833c79d01a74f2f415c1bcc9048d8072b51698;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h209577bb6f058400c737d84ced008fec05c4b3db912bde1dcab014a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1429579da041a83027bd5aad9a43380d32ba921aff9118ecc9afef284;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heb52756e9f9f98bcf61fa4791bbe1f10551f7c44b0f4998b9ed41fcb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9cb2ba75ef80985b7e193d85eace035288d47ba8e35d557dc7c7a0df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12f7ca3aacbb1bf191e3c14fd87fa48f03222168179e4907a6ed855fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1383f918ada698bea1e504922e7ab834e3c8c3367396c5924e588e45b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h133aacbef9bb42132deca51f19a6396c01028057527ec647a513f9813;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2f3ed23ebf7f6d4bdc0d231118fb3ac09957dd26068275696cb7f610;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190ffe0c99d7c6929b9b0c58a13449ec28c48664c1325ae9e4baa012a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e745d46f3868de1caa3a1ccf0e8d57955214fb3062f0ea2c4f9e372b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h60eef38bab4d13e413ec8246635ff63c061dfdfad30ed8e7f7846669;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h78baef0fc5b911b448e9a2795981ac0935ede01bfaac35776a610ec1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h78c55a5b2a288aa54d4b4cb65c47fb98880f9ae6320033ebd07295ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he52330757a2b5ed2d15526c3b552c7cd84d44760b34f0639050b19ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'headb973824c6fd1f298e06348522a2fc6146701c0a0b0db6c08601b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c9251b9b751663c26fd1a8c28d43087883b4fa99d03c4e46a430952;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h274cd542081fc43af25981fbd3ed3ad1d94dc1b8e7a40e1fff5e6e7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h106036d8d6208a245ff32ecea7fa0ea2c1e5ee6d07af7525d2c947c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc206fa5a4f0513d8cdbe9e0965f0b2f1fd67e17fec3ccfccd5ece4cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcf9be56cbb86696ff9fe51b89384b500811bbaf1a61d47c3e0614c68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4517241a2540d8fdc204063a23b7ca0634bde39530addabafd9018cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdc4fff6ec07eee57214633c0eb2350b42868b51ccb0cf157cee0cc2f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he959d530d0d85940534d16891c2f80b5b557cd001002a83ffa02349d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1214fbe43db714ea94396d1bdb4383c079952aabd34a4773c83f1fba0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12d8ad5109814e00ed98a58cb6de317a7f758179d04fca1b784c5c501;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1844ccd404ff29395cb1a9b7e4845b0a1c40e3278d5aa50a0e5e7ec04;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h527daae31aa7481b43abadb2f4c9a32b6b7295e729c7a6c519be78bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc7773ef9c3e7dc5a69868097f10d424401d0c51f5c450ca530d7608c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6f3ccc82cb45dff4695877507327625f4d794438b6c3bb261da25f40;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc90322cd93b0431ccbc9e710612df19d82562a6f53fa80828ee8071a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h88dff381130904ba44bbf41b544404ffa6a5d8ab814c15fa5676e1ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2e3b10b9ab7ff66330753722592eb4d011ec8809d93b741ac11c6d9f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8c30448fac0b7cee299c93fd7db9e03d53244b8978baa66194c3a99c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd860dfaafccc748ff9063add4bfecadcc6c852722dc950c24fa59f22;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2fb9202969414111ebe829ed2e6f4509f29ca1d86b7679305a314f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd145c55964d81adfb9cd4f63f1ffca64367d21fd44bd708cd192358;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h198cdd33fe022fe85b6db4d8d711a914a7ddfbb4f2acfcb361a82e70b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h190345534895f67c17408271598adfb28215afe234be29f68212d319f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha241b563cc88877decc530d4061554ca5bead684f5025f11ec56743b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h513d57ec7b839311fcb9f5692d74f268f00e38142c1cd826c23b4e39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2dc2d17bfe7539f9996d4572ce0d40042b5361b29a6eb5eaebbcfe72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h67d20bbb6337e74ad2c132193b1406f42e187df4a328ff38e8f47f93;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16b6ad40cd05435112af58510197213c9f50289d46e89df7b8d1e938f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9bb4780e9b4954039a648c3dbc3aa7b2bfc1c161afc9f9faee4a2d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15dffdf7203e7d7408121e0a4a5c4ab3bad87d93b280501dc27f25ffb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h41112c6a2b03b8443b8d4b74bb4d2022de41cefdf5b41c57f84f336;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6309b6036b9c98ff61525d8d6a966fd1d907ef9595e6eacc81cf011f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5ac202ff67e50a2d8a90ec296b41c35200548602caaaa2d0a7e21c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hec11a2bd78388ee4432dbc81af02bf62fcf848f0134cd9c6ab93cdce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h26bddd6237158115f6996376a203c6b7f15e2dfc3fa55911c01d2654;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ebdf8acf77dcff85808aa338e0b5f476f792529facfdeadd182fbe30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b7e1410bcd748e1898e10abb15ac8d468c2bcd75eae9ebb86856fa73;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1270acbf06dd4e29abc79aa6dd4591f6248d67d3a742852be7c78db30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9a37beb9dacd7e13eaef78df5be827a19d7c4dbcbb88e1a697208c89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b76b11031d3834a286d5dd811521d47d19f1635c2209533ea4439f73;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1995a17cd1b5fdb66f4861ce9c6e916501627bbd120c72e6523489919;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc1a7d3f4bcab44c182ee4f04e1a24564bb11eb03df3031c239d02890;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5369a19f1761fbb90dba40eae4f5f429b45a1d3f086a5404314b20c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c0b33cd161f427f4cdf79c8bbed376cc5eb215681c0355b4fd42d06b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b77299691a684370d9e5132b081d13fcb3b9ba604149c09f90f85f57;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1841e691e823ccd5b12d3c18d5854a555dae15973113f3ae819865f98;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha7fbd581c0397de64a6a3b5094fdd5888849839fb05991d0a5cecdae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4697dd8a8c316fcd4c538fab2274bc084483c5cc657d6adbe390a9c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e0c761b2add85bc324e67de0b33e709a412d8074860370af8a06bce9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11d9b276ed307a10f64fd8f27000753257c1ea459e82b9de26d4c1e36;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a38963f60298d0d4f6c57db868b913ac1c688138959e7b05fb319e9a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf5ae84e2f5355b84aeb90631c74df2cae0e5644abe7e30332bc79977;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d648fb97ec3ae0192cdd522c56ebd03bba9ec7bfcd6b922e3a68292a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7dae1f2cff82bc8257df3576d82ab39d0e3208e0aaff4a851f7df13f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heaaec471c505c8a329741ffc059b97814f023936fab10893c80287f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc45f1690484eec4489a9c38ec90ba286ddee58255f70c1bb1eb16319;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16cab736cb89e65470caa77cbb720c4f8bd255213fe6bb752d5cde7e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h257998c5406e8d9e11cb43172f7066b4414a8f6d25537b926d3f7319;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hffb729037b72f308427663c06f8915cabc375994bd79a9e9f44ab03f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf62e294fcfa4439391121f0311863708857ac211a4210efb384b9f7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h140b4d1e56868ba0d9ea59836aaa5a5ec8f85363a3de22a573655488;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heaa4177027dcc1abf7bb24844132c9ddaf4b44959f75ab3a1265bd54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5c4493ff660a69d94e2e4db3e9a02acb14540539d40e105ce3f17747;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b403721b39332be1889afd6ded7bf65a7a6a0b4ef1aa1c090b514e87;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha6eec2387149ace823442732040e82c76aebd0f4f827ed2304e0cc3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h114ee52ba2fdcf6eb11b71d1d51d68856db96747b37efd70e622b1377;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h171a7aefd785c80f790afea95f825d0af12564817690707349477653d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8d77bf0d23e73fda4dd0b7068c0ab5912b77a368178beb8fc6298978;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2397605675d16386b37b738e20a3db4f4d0bca6f558009c89a839384;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf46905617e2b9cdffbe19828c02de2e7f9a3ae5610ade95363dd9be8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b5bd47e3aa3bbcb9029b7bfd84a9a5096d65fe114a04d2d80ef1b193;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h478e6779eb4115f1513ea53724f0098aaf293b79d07a5f5f5ad94c6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10b3bd1ec32e0c556d4ae4e8f27d4e9e0ffc6166154381d94eac0c66a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6d160d70fa8a4ac687c34a1bdba45d2a2cfb5d43529d972756bc18ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d76d28632f67f1d41605b7fb9d483f9a17507842ac81725a1970c45;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d6a84ef09e24ced1cb6e57bcf75f82027bdb0d71137c0d6dab2aede8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e685846d9624a7a40e2d7e4009c3285409037fbb4c8c099dee09a33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9a950e489c7223900c7b31ef64c6650f1eda579bfcb2c8bab8c21ccf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12779eaff715376829332f8e8fa8aadde8d6ea078ab21f64658a3743;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h21898b55fff7bd82a052573e82d87c6d8da501bf8bc232cd8c899960;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h155544733544556390950959b1286e86f4860f11f1f90e0a5de7f9585;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15b27683be02122ba4a6301282c69a8d21198f874d474e0eee8ca1344;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12b2065973255f2d17c15db1b31884cdb88c0cc443aca486010cf96ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h79b05549855d1ba07328e847dfeb75fb2733efa5d15a798f32d89627;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a3820e18348eafbb12feaf234bc8b24b6ef7f7f826a14f44f2d04d50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1be4f7d59f927b283970f76f276644f670f4b10342ebc04c1c686d681;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dbff32bd4796dfbc99aca23cb1717331549b5dac54b17a0d98e3107c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10e0c091aa35f5501f6288f361c8eee51c3bab9d76341c9b95f959641;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eba08c75e8eca08cc7711a5332836981bfd87faa6f042d50c3fe7ddf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcdb6e5d9d9cad44672ac6a6b302f9a29628d09f34779d97762f92425;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbe01fda644bef0930a0a5fac08a8a472fcc354790d9b1ec741433425;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h533f3bb1208b056f53ad8ae5157a4da6169b70948c68cae70abad81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15cd7e9a0f0fdb4ec6ec409feda6596465742e192a4502f37f90c8ed5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcf1555c8ff91d6da669dc0d74a8ddc8735033ca9c8c9568bfdd8af07;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h971a0dfefffcd8b46b283629b05cf38fb5564987a041aab98ff39a0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heeb8d9d4e80ad7d2600dc674ab5dc4c7e8347636e4d91a8e1c4e1f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee24c2e3f1119886916afdc602623e32421a9e1bf2d9252affbebc5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h272c4f7b50b12ae0f8c13294e366c80c29b0e87aa386ac11e74437;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d874317dbf42733900d44a03c87e39752a6aeec908281fcbd6f2b72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h546d968012ea5d8e6514b5b91b3f8ae3a6c3b74640eb7ab38c386199;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19748671821ca165b0d67d4c50e21b3de84aac0105588f6439278e5bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10ae9d73e883d0542e4bd684b1e394cefe2b357a38bc2e8719280226;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h25581450402b8b979ccb9330f8ff36dc9298fbd89950c2460d81b975;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd32695e7d958736790b09e51ee183023b7e4c021946a04296f937e2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfa00ae2469492a02f56417e7819b1f8832e30f5a2529bc0eb94e4124;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2888bdbd2c7a66066646dbd6d190c9b540a58fee9cbd295634fb5ea4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h105b098cf45d4712870069c3221c4bb2bbde62a2c122d73d24134e25b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf28cd37c529e49299b3671634be1820c398eab4339a906c533b615a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3620e78b479ad0445ec3f129fe24d1edf82b15be6c2544e1cae81869;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12ba8afc1d6a169919bd814ff0bfb69275765a397235b60d90166201b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h168713f2b25ab180c8976c157f01f629f4e189c98f4219e9afa66a852;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6ef056755f9d6e81ce8e813ed9dc728506f45712bafdd556b48b83f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15272517513c295525e33b915323e8b628c596092daa635b65b193c14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd183f02ec73d4a1cd7342e210a6de839d15f409470f9c85a1803db76;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ec288bc6ce004ae2ff6a9796095e7b95369b53ef733598dfbdd47811;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a2b73b911f140db928cde47d00fc30081e0960030a2b8b4965e9647b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h174ad29092d3ec934f717d1de63b840b12f53e2589e2e37752ab32179;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86d8bd94de51d0dbe6b0df211bc1f836166b62a100e7f3a0c05547a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7b96fe911d9809ad8fa78c41c710322b7294825d8c22d2ea02852f83;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h131172335fd0803324b5d6098884cc077e363191b856245b3fbcf19c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcc71068fccf3b45e98ed54a23bbf45b1fa07b554cf05fd7567d8741f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h76770fef9cfd5bcecc74de80d0ff9e65fb4796fde26a46153741ffae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16874fad5dd35d362b41f8e136db9161d0a309369e6a5a0fe8ad4362f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h189273dbde0708d7c973252a0d63e333408f8c701acee7dc25ec8ec19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h768664fc0001e2a75a1abf330ccdad892cef63b6c1b69300312944e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4b63ed996d2586ce93098316044cd4e05351f595ffd0ca1b7bfab8a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfe7867e947aa360add8cfb9a4113783cec304e1ef579918adf641674;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hae824aebded1b9ea09b57d51aeef44c88e4c27514adae7f6319fe0e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1da9ac7b7004366f19bc0d42987d7e7c970bff07cbc6dda8272e4de13;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7de4766278747e76ae93bedda0fc5f43d97228c7f7e14c312fd26e34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd1bba7f8137724e9f9cfa1bcb1ba3e2b8bd1805aca573f1a79acd6a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1499eb251c90061edd1b4c6ead8e4c2e314e3c51bcf9fa92c73eee7e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15a68936f6fd73b30950a47b59d169b79a9d7db62f1b2b5f0035f3288;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b8f04c2df9ce758972d76883f6af46ef0f8111558bb45bce70fd161;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e66c7cbc31d882458629773689cdb6c83e3eb73bc1dafb5eb5efb982;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h118e5a48aba0707fc462fddf31c4a4f6101f6ed0dad1118cb84ce2218;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb489668ac51888634234109d3649e2061aaef7d94d10246e5177bfd9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f12cf598013275c016d586ae3c06ca697a9a2731a1b11eaa3d6fdab2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf97deccc4dda6a77f0f1c327e23867cba3074ea216d4aebf620c896f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a64e191f15c30d7c4fefd9b29081a8eca4c50b7c41bd6c1f5d6fcf78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19a81c0e2d8a6d183d0b35404c3ad34a145d2a72ec667e335fcec7451;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdf5eb256a0dc4b758521041e6eff7dddfb1c4cd527d00e4aa5766eb2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he08cc8d1f97049aa7a1d1c95cb68872624f2fa1b927f589b84fa76e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16767d461c911aec8a9a0680c2bfd57ba3a831a6b0c84c79bb19ae6f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1856a1fbb9898e7258f3cc5110608e85d88a3a5a2cf80489ed958bb57;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h40677eda0a314986ef75a4981976c55859132099418ad3b504812cfa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17c667375ebd7bc3865449da93d9a93cfc7b0b868d2d5e98ea35ca937;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1083458d1ab346e5cc84cfc8e2ab390a231c657692be4a81118c0759b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14b31c92d2905765876968405941a99def6c964a7b45933e620b4d09b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h174cfd9288bb20b5d4da958d181b5bbb39500d2c59f1134839163a2a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5acec5944ab489790e1b007339045164f2d0efafcbf880079bbc0d68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ca030cf50e42029a976d57510c40099aa9089280fad3d9c9acb22ca6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h142d1c07b830ee958f338020e123ca496a1a0cdf8970e2a573a1f7b34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h223221144cc2a5bc9bcaec3bb26b8dd2e2cb5637ffbd2a2d58e6b0fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he82a24208315164583374fda719677c766289b9a02ac4616849f8d04;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h604d1cb48f9da5bd7e60539651ff0c233d1f0bc6b5319d31900db343;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b35fe61ee9b76a0acec93b3270e53e9f5448d72b98f3884b5ff8ba71;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he8acf51e192d513a73af2d43cfa900a8e747c3c119d954778a67edf4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19f9b7cdba2e44bec5685910311e9174ca365b2c36ac1d19975f2b646;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f0c779184e6ae6bdb44d4aa5e1448f0e817ce0c5b1bbea939c247fd5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h189b320b86a2553180b630a8f765a102bbf6da3921e634d1205ef557d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1743c355ae143e5d60824706dac59956e4a772b5e55f96f170367618;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h508e5d6244abdda33c84d4df3129eb528da6b8010a04ba59f484775b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dcc6fdc6a1f708c8b284d00884567605bbf1b78da2211d02aeb871cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha70887617a0310222b05811f55feb22b0e2f817ed0207fc5944ea023;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bb14400b2b39caacb1dcd95ce8fdf3bcdc564e9ab1175e65454641d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcfda9961877cb9a4bd57f61df87d83820c40dc84f97e446945779c31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h138d7dc309b50074e5bb89d4d370c9979b93f2e6feec626110b590b52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1344df1991f8c1089ad89f30f441f06027456a9424e5327bdaa5ad333;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc303d0e0f3193d91f4eb885e5b3165970a3274f84f1d760e3bfb3ada;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb082b7dca805a87e82afbbf3c9fe4fa2e7ab0576491bfc242eec4faf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11d1de1209e4f13bf05fb4ef65be0c399b43fa5de3e1dc8635cb1271b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15dd60db2eecc7d116f5ee3d39fd024a25cc8629ea87e7d8e8dfea3d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hae7407fbcc288b2235a3406f35732293d47c9239785e93ef8ef0de77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e9a2932bf2e63eb2521081a52ad36f43c0bc418e5e7cf7032588cc12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1beb52b8f31869032b524aa07bde8a7bb7b3cc914b5d7309e20c3d084;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hecdc5ecff4a958e1bf749d651915f76fa8e148f725dca93246ef0617;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17febdac3cf8fe40a2367a1112f8cc54c4be6371f29089d5c71e1ea5c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ba2faa183163feb51b87fee32b621017923321e9024fc2c59efcb927;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ff7984a4b25638d8bae922a06b7a62fb64b6a62bf5ba550f0849e3d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1679f76c2aba2cdd2fca9566366155d09ca7822ca4b152dc05e570623;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb52f65b08e53dfe7d591a915d905dda742fc206f4f076608eefd0413;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16d1ae8a58d5159603ea233525879f42ceef0f2bc10c98ed2b127156d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17bf2de869e1734eecb0c29cefd9b1b51e781e8390c2cf5bb0a602d68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12066a46d42a44562d8e507054eadd0ea2b2dcd50ed522d841be5021;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3cce79236d85c27574ba27f11e3ecb54d700ff3abd1727292bc5bf5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h131e9449253b4e32e8f38fda47fabfe76b2335b6627689b5f8fe41d5c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e886e4a220415d3a80f8cd66229e8ba77b803d3b87045271ad49384f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b58391a27b40f482f7877b74fe8d201e64a7ca2bf3083a515659d74c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fde970f78ae116ef08ab0c7165c51944756c130daa03a3cd2430f3d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6a5be093dbf66d35737462e1c6df8e666d2424eea4bdcb1a2ed60716;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1693ac9062f492bb2d89dc0f686d4398f5c2df6c2afe5e1fab7fd0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd224f043c22d6bd016aac4c5c71afd19e81918445880a61476fbdac8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2a7a8b9fc7cb9f53ac7b3689f1bebe3c5766732646a2f3b8f023be5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5516ccca75b2e4ddeaee9c791f0a88a1cd55f5be0ffda1ebc323d54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14db033e4e4321d82078f3e5e1524ffadf2ac3b90e0c9b0341a4f928c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14f232110cb0ce96d08035aac908fb8cf1349a00ad39d7e268765e040;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h166dbd31eedcca1e30f97fa23de2a61d77d5102783df5eb81820d7d94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hed85be6f9e169235ba2441974bd1c9e4b85acc88576dee3ac2d410ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16f70100713254a89ede4cee0b13c8f4eab848a3ccfe41b2899122b3c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc2b46d1f09359b7f089642b823177d2a356ba0a72572a993aa44836e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bb9b663ec64353a7a902644353261b7407007dc69a15ec9313a0b0ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17670275429b36c447274f1a8f5558493c624edc04ca3bfe3d0b551d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h69b36aaedef00bdd283d3fe0678918722909cf794de75ef05b24aeb1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h445ba9489440b0adaedda057b7f8a90be6e8efc1b9cba327fd55d0be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he8a59db48ff3a892900f6a00e3903135d075e5b388c20a41cf86dacb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d8b9e6f7b694364f381e95a087817e8ebd88ef714a40907a3743fabf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb2392a711c37882fb57349dba1275a39c44a37c14deb93f491c0317a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15285b8add3ef4e7dfbda85c12aac7893d3b3b41613939e44890b9c86;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7c3efb0abd81bf01c78daaf6badb34aa3c6b58a59ae954023f9bc62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h98fa9ebe824d620d6b09d9174784642e30f77fe9c9a25546df0d19f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h279e4ab1b13bdb19b6588a74c9f5f68764b2549c54b72aafc5bda260;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h47064bef314d5276deea3e1cd7ca76db67d78078e43c9589f37020a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11dc3d8854b533c9dc3a800c2b596fedbcd69570f732cbc8aab4d4d5d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1650aaf22f91b6d96a0d12eed17a32da33c8f162a74bd5a194adba87a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8b6d271a361799a16c58f125ee942ba6d6e987056a6551aaa22ffd2c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1255f93e5a907a95e0c07a56e905f7181767059683ea85220a20e3ab0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2440545ec59707feceb31c020c956232c2e8cf98ab57dbee1c79c1f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd0662123dc26e78f63522cba23d01b65b5262da15bab65e33f70b70c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17e10a898ff162bc5e68f0b9d4c9ae82b42b185b9499718739f18432;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19a76f2ed11623972569c186bd219033fb7c89cb7c106447e91e8219c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7aeee534e2374ec3052b552e85330ce0a916dd66fa39d9e1e6a4343a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he209e10d32d2ee286d83d378e4e04e8f587a5b66bd8e83efa969a76c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18d21234a9b3929b220ef1f5783d80d3814355e2585f551401fd96c89;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h38c143f52fc65daf7e6c61e821cb1e97a8f886ecd80241180bfba3ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13c6728babc4dc21d6dc396602cf54781c464060754733f8bdd0452c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h70055cad68b2d1bbe6a816062f9ed3cf69079f999d1775a99e559482;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h529b503555d2f14d1d30c6b36610a4212bb6a7fd385771214c647569;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18d979383bf1bd1991ff2206eace0eb9630a39c5a97efb2f2cd631b83;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d73eb1f59cb3e278d58d9addcf2d26f8db24b6c66a49739331efe9d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h72348f24d0b85e49bdb4ee45537941ec9f195aa63593b520b1b55cb0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h38aa6ffda2f066515b80949d89b139c40a582bd236efdd7d894956b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h187193dd1c76174ec2539f802c6de41932e7b6a6d2d672f80b58b7b60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3f3e00b478a9a835e5dde36dff085bd4f8228b2a0ba994b2deeba553;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h133939b7a12692329315153109474d4720a8c1968eee423dad7ae83e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d258dfd2ae10e9ee0488c622d3f469bb36f277e787b5caf81d7654;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3cd6bae1b52a103da425194b75b527b634990313582c10de89c39a0e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h444964aca87d02845ca52ffa577fd3266c91f28ee3c1a15930fd5b0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h152c2447f0d0746f642cb2eceebd62895f39ee76699fabbc91f4a2f5f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf08f7585e1bdc592dbda604ddaff00fe5535813b3064ff0e2af0d69f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h74fca1ec7d153152325f903254bed4194c123126f2a92d1d90d3e034;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf43cfda72bd6a09ee4fd14984520836f1e0593ffc1d377e897f35114;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7a09be56cc0eea5ef3775856bc26c63a020ca57bda7696af99a0a911;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15bbbb4a76794b6584d2ee43b90e9b5a9863be6f4a85155ed9078ba03;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hac4e78a88fef1464d34eff78604a3094c6fca5371ccdd7ab22ffa1f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f03a853d1b3bbfe6dd0b7b5f8c0a50200b44838b3537e93eac22af2a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1170da00709b1405fa38a83df70d60eb97d1edb5a8c2e7cd1d4611ed9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fee39eda1ec5c14b115e0594274eb54d3ccc3721bb216cbb0b655401;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef75c1940c2e69e007ca66da255302eff7e327c9fc0a25cb4a02a2a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h146b2498739474c5431e9da0984ca0fab4ce65fb370841f9eddc80562;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c7d8621aa3c0454d093efed3e2826836b9bda3188b4853cd8ef5e2af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h185b8d2a022e2c591f5507d0ca148c4f6935d1541cf53b8c34d5e248a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc4e3dccdcf3282fdff29e41cfd87172b660ba1b9ac54255660674477;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h70549415bc5ee56222cb41c71b4be2e45ec7762e82aafde325423b24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h184cd68bac85d58eb2f526339a1d5c9d0bbe82f2545376472f522222f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h153500103a4291507cacc72f69c3fba368b4911865729ca1850e8f014;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b1d57ac6c37f4c67c28a08baace807468d8ad43815edc006bbce640b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he8f244d948a7fbc18cad911b688ddb99f296134a1c685f7272870d92;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ec50120f8a85a3326d64b7caa1eef11e8f8c7ebf58c05510b6b5dfa2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12810f824ad0141aee84e420e075d08536dd48792d136bccd1a1402e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a7d38e16d6c1fb56018bfeaaf7e4de504dd4a3cc34b7cc5feb952ed8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3964c74ddcaef7568b6fb6f6574461844a3b41ad329a5e36c77600f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d16a27f871289109057c8385957d2c31e43a199f8cbc0c1e44582c52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1765d09857ac54c9e1239cca82d8b0be145fbe37c88eff2fa9407bc55;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h120e23efa59839575a81b8fe004d70b66dd48b6f9558109744e94942e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb3fdeb668fb23d5e8b1172db87a240b9d448292e37669699dd768b39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbda056f6fad3fdab14246c2db98ab98d07f7390072df17e5e23aa486;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heaf3042a43063be60a2c771f001cab638b4e307b1bc7ba2f8c492dfb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h56857a0210fb8efd41c745be567cb72842fb7a342ae525d5870510a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dc5b07997482ee39778e3a9b80766e1858d2f7d9b2d46c6e378bd670;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a6e770436f3a0934332e5589b85db1d7382af236ee21ee6c271833e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc2e415e51f098b9e8c22ec25c875864752b2db8aea2e4bd8aff77218;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13e4140277745a2b4c0b3fdb1e533e6f470ee2c29027f06909284ee5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15eb6ee39fbb6a4e633ce653152af8ee94d025e27094fa1b72f972bad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h192fccc661b977f2cb6576c141c590833f0910b96acaf413a415e142e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h191c3c345d999e20bbf0a6c22983aa96083295ac6a2047dc19137ffdc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h139fe23f4a83de6706fcadbd831b2b3163a3bf170ff96d1ca9bc3a6c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf5d1466083872049602dcd1ebe368247948a17f66fd3080a4a1b0b72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19f83beffed5e3add59346720de119df8ba21026f7dc41119a57e746d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb6fe2b956c784d8b07bb286586d25ac259a0be39cc2b1c5954b25322;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7557b0c13988af2eead8bb462e68ce7c4708ff23729a0c805cfecf43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6f96e662ff4be5690a497911e2c6a026a8e2f3e4742d9f20709b56e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h194242e2b6cee7aca97b0a37443885555d5313c9911ca5ea5322464d4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h942f8db81ab7dc73b9680a709b703aa92e84f659cfc68ecede7db5e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb1f6388348dce077fac3fb5c3eef76d89c2c7231ae1f6f4e0d01b214;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a32423310709fd4bfb6b457e0277008e7ec19fb47d329f8059bb978a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h53d2793c6ffe886f054aaa35dbee52fc717516a6f0a70c66f31cf94d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1249ab33cb76421d55e4ed6d89209d5344b69429b10efad1e1c030a95;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cb10aba8ded5c0cb1f940c185a856c3de596d46336d220c39ccf6305;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c79b9dc84da818237acf2cd2fc64dd14a20f9e36b72bca203789dcf0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h263aac4bc8259f4c5c4afbc4e6606de8d81ac7e16ff087211cad6e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hfc5379a9365c07f23b0443d0d9e4c3334424afb978f098700ab1562f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1374c93dc029bed691937c213d2c5833f1885acafbc699b6d395a3473;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18455a44e456ca4f68bea0aa0f81ca149d19e4bfa5ac1aa43b33d49ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fdec0128960223a44b5316a3a14a041c7fbfe797e3478659b9880d02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdc02bb7a43110248c5960ce9d3014428f31e03b8859c8a82d9428e79;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd534370ae438420b134c1911e7789cc6b50770ea8c7123c1286ea91c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h928c01f7466971fbba2e30137270692748f6c104086ffc405f7d6870;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hea7f6a135e0e5fb5d0051632ae696ff1bda3692264182acb1a91e84e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17387060ada11ec51a8e7012f8302814635c0fac76f49dd4c874f8108;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5677387cf399fbb88cea4503d1147a2c124448ca638f8d48af7365a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a1ca74db844c809df357342e0eb5611f534bb01df5dc8c049f4c78ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19721ede04e1d098a07b6db13f9370e5a3b75c83606de8e982684b49d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h134ceea1f833cdd2754df7ff24c29057224bda7b54f0256ffdf5f1c29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d726ac1c4a053ae8a854d1e07840dd9a1068a4df1fe8d75d7d8a3cf3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11b0c8bcb812411598701be8416e97dc2769fa3cae0a5ac7ace750ed2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h122921c309c741f5b9d2198941f659e1584cfbed5dfc79e2bde5f8ab2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e5fed99d336bba1c4bf9bf5e7a3f62633601d0d81576ae6f9615889b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1acc10af4c0c56c3fd5ef35c2e43b9cf9674b8cdbdb0805c68b10cc5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1247103727a45f4aed151a95c14c386bfc89f160ec51296df8e1319c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14f8667c446df41645b5b089a84a273c20488bac388124bf7c7137071;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h95c645cee6ec8d0dda35408020cb64ee1fd617ed253a70ea3ced5b72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ceafc2fb211c320c556a5e0b429801e770723505c7d9a9f2f3847c7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8d7e61189ce7e875b14d2ae998dc8be64a943cdf3837792dff55b479;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6a3cb2c93a77511d5a3148848b035d02c64a2c404bce68d46757d146;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h139a78606efef287ef47476ea0f83f222a6f554346bcca4eaea773ea5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fe8a2e9e2534beea42206a77a41c1b09744841117c3d4bd0446a0ddb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf66991619d4ae96a59b388707a713c192c91663a534a32f55ee03bc8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10f796bdb0923c2951778add0999701b8517fd43a2121ed292e673abf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18c53788a0582e908afd4645946ff912cae71abb6eafc21152a257c37;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc2edc61d533073a07623c94f63fbff58ef55bd2db96b5a711938c321;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8102be88f7c143d495d0b0e70dac70eeaa887aba65fcd9c507856d78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h74becee36b18d4a5aa696c9c3645cad23a05c899be36fc092ced2daf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18ff3618b97eef0e78574d8543af557a448129d9015d22c31fa778672;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h137dfe0612376b0e9ca93b8b8b0ea79a052566ed8b457c151f878c514;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8daec5778f58fe96d8df1499f9f76c2786b5c60a7b2ba20e7937b89d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h176c2287ba274367b18102269b164f730d4a614b56f841d437b531846;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6e29aac9babcffe91205991448a19eb176e2564f55bcfbe8dcc17b7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10867bb0af267a9f26aefef61eaafe6aa7cf37f21ee722b70dcd76f37;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5e175ffeeedfc02ec118eedd59237544ed8495722b1a5e8b45dc81bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h90cea953a0337a6f9489fefebb775fb912dd0a5e86a07bfb2ddc5412;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h118606afcc17cc71492c5c0a60cfccf61620a839582ce6e024d6b6350;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6dd7f18853a67a0b2a7e2194706899a2db6ba7967e9fc9b5769311c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h177e92ef9c2d1ec89414eaf71d4db45c3b504fe7e1a256e68d85017ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc5dc206777fdd57c3a303268ad5f7e51a0f0cadc21503758627cd3c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5ada3446ad85922c7f675a87d80c3098ea8378f9d58ba5907c92dbc7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h137a0aa5e087c2eafc21ca9fa6e4a26acb88dd61ef231e24650fcec6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd3ae5f9dd133b813d8f6c8946ef5863456ca555702ddcfb02f0136dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h177ecbc85687ace6ec9c1e7208beb9821a3d180dc76fa5b90e376ab81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11f695b8e184e63c589c23e47655676584849a3dc32aa78f346f2e6bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12e3f1903ff7bba99d5056de995387658fdf2ca9fce39c1e1257395af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8b7531b97d772cb6f0df5b7c353dfe912b37285cfad29919f126c976;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8a86b050e8668e3be96cb938eaa02fdb17e937944bd28cb608d9ca96;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf9b1f3ceb78447e80c9a2e65e57a67de0c4fead59270a35606bd866d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hff626672a7606e905c4e570517f1f0305d3d0db9d4bf4af64b4d4b8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5dcfa929a7c55346fbfb73132d1d070eb5ca456cc9c85f12dd01a5ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6b67f9d623b505341e6396fa623ab3efe8f063adc725aa86bf6d0a7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbddb521af5f3d5a211f96c12ca2665070d35bbba462a65abafa52dc0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e30e3ff666040afe433c3d09c13461cdd78503a1fac5811fc3d457a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d6c257c65d148a8cb37c665ec29184c2811ec779d41ddcc488338ffc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h48961417564dfdbfb6c9e103a3cfc28bff3b94acbcbf1be5ca078d15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h139331b53af139248d85172151c9a46c8d70499b6ef987065b441c68b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h171b877cd25850fbe9411d50489f709f1db7747a4e8f4531de868fc0a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1584e2d79693174725df8f1a13fb7daab4dd052ba7864c52ae84bd166;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb06c1ab029bd36f763e2aa3ab967e9834732d0ef549c4ce5b07d423b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bfc865208e0608d7bc409560b994714d6f141835aca99b79b421fe6b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h20f9e020b30c434aeff1776fc9e566dbe0a569594320a8c51f82dcc5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hafc2f032a7cbbc1d06f434ef4aa5186e9755ff592fb89500bdbc9e84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee42d379f4d77cd5da8d484abace072c9833ec2355e326cb904bbc68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h115809a3c245164f4f0966c2b9452966c69e0ee77bf97bad5747fa471;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11efeff72da2d5c5aee57e96b9d646550aceaed5f811663cdfd90cc25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc20b72501a9d89d9c2d1d6fcb0e3e46ea934773d3f2a2599cab2f074;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5d0e7be34de55c8682d5d87ce56198cf731a87b39cb79867366a8279;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7f36e0962892763c906c0f2ddd579080b2b881eb93f6ba30e82a0abd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f9875c33be228be05c2535177ba8e93a7528c7d8097cae8f46504c77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he730146b92482a8a065431a88a2035d80dede5fe26d16c40ce7c534a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6a35e146f3a2f2deb8c2ddc99520cc82346c905ec400ff364b27665;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1afaeafc8a84f72f1f938830d785e5741ac59c6ecd65b80b6622224ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6222cb2056b8c4db12ff4409df1cbfa48a18f3c5203e7e8165330464;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h731beef63dcf1effd3a263bc7810c4041082ae93ed7fdbf5ff1fbc7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bcbb8cfb5df21221639add0a743340a60149022145913f7486abe476;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17f01555cc52110752174d4ff9c728e9840b474452eab0136d0997e2c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1929245a8b3637a69fe0cd45d85e54609c51cc389622ea9ad9735bad2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h125ff4500d0d96ac91665410d775ebca8bac936fdade93e4150ee67d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11ce3968aa9115c9b833f7a88629efe92e133b071b26a1c7b6d043567;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb4f856dafafa975125a229dc9b13adc9c8cf060ee40342510c77b5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb68f53bb2b10524f1bee38d4901525b8aad083c6d350e312ccb1392c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11822dc6b02ad69a3983463085adbc5473e69dce5b44ec29cba242d9c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1142866cb0ebdeb80754a54dc35a00ed2a08d0b361838c38a0a284208;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h705873e2077c3d8653c92cd27d47df24f38073d2afe7f7a2be9b5ebc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hea4b00da73704491524378a6835e3ea7fe4885ddef0f304bbb56d13f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hed562e6254de0dd81d3ddb7a81cf126b5c217bcf8aab0cf33db0864f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1302433b3ceb90a2b6364ebf60157b30de18e8cd20d8db9a2696b653e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3cc8c51ee4ceaea1b13580c52d69baa8c48991c4855d18b22dee2802;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f15971b8675ca6b869cf192b28e0e48f8a95efde8d2fbb49fd47d465;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h417948d8ae68106b96182db072bc3f51911e1fd58f000dfdf1dd9b02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ffcf225e906d9cbf4611b08173558b93a4e89b3f6d3f0f049b3fea30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha3357cb67052808624cd14f430b8b4a2771f2710047323d8a6994d75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f24e9d8b4dfe4798fa7696995e099456ae526bf409e84ebcab64b559;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hccacb6d385ea1ad680fb9fbcd91cf15fd2eae13f16a8ca20068f9f4b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ed646171bcba661c6865b9baf33b87864e3de3496cd0170ab95d9b85;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'had610010d6087ed5ecdf741a90f49b2f87c5396affc6510312ed75d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10911cca55f7892f03fbc48ffb3b3624ec2960fa7079919565948fb28;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1873b493134e8a721014394454e99f364744d32d501a5e739715c187b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha45b55b6f5659c166577b30eabf9c84552d75447cefeeb6d8e4531b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h61928b555b6915d3ecbf6a1846f903525893b7b189b15f1fb467ef24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9f01add67d44b84a2f84ca142c5430abd49777bf8681d2cc734eb6c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c0f8ac685b51bea10bff3cd3267c3a585d733ab722502c54922fd913;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h195730a81017cc5d6663e38765bf5eb9d25c44213ab2f7856d1c2ec50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1aaad8d901c9fd9cfa4e809f5b4feebcc465d97eb0c2185f20f860920;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c874aab281aa98e06d84eace242485cbf4333bb9988ba82f8a8df77a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcf5815b0dce0c197b527128ccb7fc3eff239b984d8e8c7906de443a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16c5f7130f044195bf664828840d52f7e72733440bc106452892164ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13444362bd16a756b111782fc94d27af0a90f2e88194ca7fad671edf9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14c0442f4c3baa493ae95f6955d7078b066c6d1b74e1c6ee45bff9037;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ca67fc968aefde86171cb4720a6be1fc5fec7c5d9796b4e01fd8ba05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18be52c63fcca53eedab99f0023b1244b64392a60aed4894d9fc382ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1db8fca49e5036c455fd9bd6caf36e28c91f107094dff13dcf62a4f64;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15d83e713ee2a6abb49c32dea0e3a4227906777983b0f8cecaaa597d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h141557dc6354ab8aabc5c8d88c9b584b28fe64c81797a784a19677bfa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bb0b6b98816835d41fb6cbdb95ef9ed6bab97287d6b73bf3d5fe267d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h56ba6db3f3c1253fe61e4058f968a08ba580498573b1f602e8f56ba9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a979d3fb5b63f49b350697f66f26d3f2f057946b5afcb701de3e2803;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16e51358ec736db9d53228ce9a0be04caf4f8cabac295b3967bddedd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b22fab40b8998a361faf55c19e7757119611d23d8817fbb2bbfc791d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf949db1754ac2607258cd9deed045a603dfed1ac8d3012c692c41624;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h153339e5a0dea0a331d8797fc1e0476e1a37480d580ddba79bcdf84c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11c9b592e911aee3bfd68a9cd199775ac950460265a3be8ddb7209dc1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha751e80face8124dfeb712f68b77db41b5a033f509ad28ef6bac49ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6c2146e0818ed48ad5ac94544766e6b152f49ebacdcdf192d7a5a55d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h479ad0f74e4742f400f79cee4aa2dbf1a30798380d4f8173a8f1589a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h82d9804bbe2f98c5555413757004092095949ba0dca681ac06eb1e25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13218e03b9fdf32fb3024cc0745b6b31813a3f1e7221d8300253627d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6054518ece8f4ac40193784483800ffb6c4b38f8fbd17ac14f5833da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8e4fb942c4bd20a73dd30bf94d3de38c10fd760813ba926fa0c607d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11db8ab96f2fb3b8ab564c600fb2cae18372519ae2ea258b99bfa7d34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7c0626bcfb5fb5d8fb5bef278cf8d526d271683c74abce66f378c09;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a75be599237c587adee5fea78df7aece17f64b2e450bcb503f9ba619;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h655e9520a9b1bb63f7fa3b34d2d5f71b854f2a8b62a2041a1cb4bbfb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he34e165315f1a9ee63951cb831e6120da189b96c9afa49908cfdaff5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19791589bfeea7713c1f40551d61ee98f9342b4dce3e211dc6e6a902c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e33de2334676e4f39148dab7326a4f2b58f2c567c266797617cbfe2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f1fa14e7d8f26ddd25bba339ebf609c144510c03e826ccb25c162f4a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hef8bab02ee91acef1992d6f451cdce3311d0770ead041246d07a0335;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11f1fc0868eb24215a5f5b9eb96451feb5c754da08956e2d4dc6ab2f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha8b9f63dc12b338a3358424417dd160677ef5157d29616fb4e4403ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dfbfa3e908ae1d0e749c8bde3f3a98b9778d852558c4cd180284a8f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf7ca159f2fe841facaee0f8b10c62172a947a727f3510d988b05b094;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha78bd89d87fd3b979fa4aacaea34a85f7863c989e647c91700956d1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d97ef5317d07f964e273d82f31078c9c138fed2ff8a0f47c78226da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15d5d0f779a1e7c64ab8cfa92de58ad1d0336bd3c98c7dd1a64e91675;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h37a3bc588deacd2a491df71065596d341c227a100f54c34ddca24f00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8bf02db8b3554a1caf3fa3c1e5185748a416aa216c6c7a31779b1e35;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h185c63835a0aac69f870b66262b6a92d28cf296c4f8e97907695d74ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19f422776c51c5a177efb9d96a7c939e32bbc5703f7488f024649bf14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h61df1a33eb9b1f33daa839a7da6b948f1650380843546365c9e312bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd8a572176996bc4f7d8775425acdfa2f100c8efd0b75312740cf6845;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h121500d91ebb37622ebeac0caf6de5e3db1fdef838bae1031cd4cab60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f53478b37dbbbc6c4b62a9ec20052dacc3b1669ee28be71d859e050c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h179b8486cd337faea54793dd37c97c2924a9dd3b9ec60c94751416f56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eab8b410f5f180a02c8601b0f4499524101246f26f68d1e6f53ce5b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e5dec810e6e623a4dec70300e7e3c8726f4baee109e8e7cbc3b4b091;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ed8c9e19f28414f28b5d12c310784b7c6ac4cf957b42103a84cc87c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h114ad2f41d195327528ed2b4f0c20b49a0df98d79b0c5c060027856c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha9ed1b9d905263917bcbdeaf2595f37725e9761abca4d843486f4430;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h174ca02d7af33301df51d53e269d1cd2de63b903ee86eebfa6855232c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18a943c72b95e87723ad5c1ae58738794745158c1dbc14dada20a08e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15abdd0e3b542fac26874a43d500e7f3d0ccb4e0d27e33c9468ce4561;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bdee3d63bb2d3ba233e062d644cd4ade3f7ac3d0bf81d7a3df791f12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he6c991bf37b6e405dea172712c740b8065835171428e0d696df949ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc7f02c8aca95735dd48aa0c8ad9dddf62a8e13e45213e4b5594777be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf1530e0661d9d435bb199b16796e12cf5f47cd033255dda6a8c1581;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc8a7a2da53d05ca047d48f16b5867a59c173b470f4f91fbab0d4129e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13ae9c24d9dd6b3b63656b35d34b7354c72de551f6a29968fe782912c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86b69f721f9d113368a41056fafa7f03b1b9d839b84a174b443b0bfe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb6998efac6db81a4cec06644c425607c379ca4dd25132bc03777dfe5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcb9fbf5b1211e63688bc204b57996654e7a718b432d1acd3833de572;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h29d1fb39de0e13e6a99f9fc118765f5b556c4ca272cd02f604f76b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4ea022e281e4d96831df06df3c6ab7f61f4a12d3fd92e55cd9cd3690;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1abdf081f756843234990084b1dc7371ad3e921c8df4de4e941e80bc8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14c0ac632114d22b5f8bd65eac10a93bd98ccad5372594433b355763b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h640776dcf944022ff4b4a3306f95e30b65ed67f073e20481cb6fa670;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1eaacd1087329338d7224be85bd2926aaad33e9c5286c5f495ef8329d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15c453e7454e94dc64b297c444171c79f0a0fbfa571c41e08c812ffc3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hda529efc9203937b729cdcdb582aa970c4ed473d9a6c924064d9f6c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1224530ac19a264d1c7d775a39535a049b73d4e8ca5236a74a84aec5b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h45b1ed35d46de72afe278162bbe6576c3c8003e301fd7165bfc5cdd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h587efde5a78a32c3e7a791c18109b4a9db4d7815ebac80653b3ed065;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e3ef9b740514ffffeb5ba2c127e4da7d42a8242c27d31f73e22fc6d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h72d6afea6c5e43aa6ca45bdf29e11ced9613d27efa965e6560787640;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bf702fc2d57db4370f90f670a9df0b250415f43c9825fd5d910ea8df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6179fcd2809854b6bed196a476b14f6d90352320bef745983c8337f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee89b65be181f4d3ac1d6d80b88f96912e5fe7995e505c51b37c273e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e5601f8914f104d974148ff73e26fdf6777c7c960203cca4acb48353;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h149fef9417ad4ae61c8abdb7579bce1809741277499ced91ba63f4502;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h137d2ad33d736bd53d7f9d58ad53bb91b2e55bf9780405d1df4b6d8fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10cd740a9a683bf070ebccf05640d51e24de1c90cfb9f704bc07c53b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf35d546fb3b88dfc2ace9e93fab310934fd75df11b519654cf278840;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ee03d571741a093c64f1258f957c796524d451d8f7b7d91f7e21e627;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e701f3695f2d2d204b92328b90f6fd7c7536ec7bbcf21877921c60b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdc8d33471bdd97ead1b0d5e242890bc7279d7028e17225236b7ec496;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11c090d502798a6e01158e39e399c78ca082723be48f7823865c7f0ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16ff9a4dd6530ef0eeac71f411bd4c958a23c969b9ed4c7bc110e7610;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h131695af47ca5c0d2181d55a6ed735ceaf78c1301d17be9a2545d73d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17a672abd18b33267934148a864d72c435270a4fbc604d09e7c410468;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb64713bef3b987f2bc4bb623d75e2db934a1c6f7e9e01047a2e63f46;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ecdaf59688e397c820fcf531831cdf0899a59ebe22dd8d5c508e809e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1143c27a72cffc9366d2b71f1fdf543e496586791d77a76d7bd4be53a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a965246a87e65a67ff4ed1892907b59db84970cbfac5d488cf374aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9e8697eae2a210e217e2cf8f013601281a50d9f483f49a98c31205ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h685f325acac559c01372b7ecc90415e9c2c0e230d91eef9481c9c8e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1688f8915b1218e7b99e5ce3eec3513dd3b00c42927067afae9924530;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h128abb7d9673d550fd44e0fa49d436920a805ba3dd2296d3dca258669;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h484e2278562c2677ece9880b25250b22c36dd4b927ee5c3e74285c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13ae1da5bad0b42d65a28073817cb5ddd1d1649463b8764a093d2707;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h258eb2e731a958c3c24c2867043f0e134455f770ac512fbad4f2040e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h889bb3a9bc1c9e629ae2f0bafead79ae6aa4b19151ef9316ae525626;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1278ff1cc8c38ac9a9e93511d004d4a99be57d7d9db348d88598501;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h322b418c51e1ca8b4ad664abe137577c86edbe79f0feded3e931e530;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16a96817c73204d7c8c6dbadbd1653a8b0c0aabd76546c67ab24c3cef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h106a99f88893c817c844621bb9ac3b43addd31c4028a2cf0c9c6cce9f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15fb744691f638c0bfc96b585af593d999f66f41511eaefdf5ef05589;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1361e9a5889a0c126b274a16604f444ce09e7a49b6f3566715ebeea56;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h173c8b49d102d28aabdd440fa3427a8af51d17ec0046c84a056929b06;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a20134a12a5ebd7f60ad670f75908b1bda6bc572e8eee930219e7ede;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8d79f8f99e5c21173e7f833eb6105b138194acd2f1fa82bd3f63c956;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hccb115e9b6aface30c4740e9aad3e1f91e941ba05530069ae241b26b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc6564f1e1c561fe7b717501105a2fa9530d0a8221bd7758b4ea7347a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f2ba3dbc94f877bac633fbdcd3795340740e52ecd821f84c63978d30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h53fab14e20a771700f29885c359bd064aa2ddc2da8010181fece8f46;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha71c710ad6b67c0ae1a457f898eb0042ba6b6b27c102099d9741b301;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d0a9310b8d5a18a10938c70b22c188624f9c66e676f537242e8bd0fb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hea1a1b719e56f22f61448aa442679646d0a30d5883514b370b4cdd31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14c9ac16f6485273085652287f80f7f15ceb3b6266a2dbeb83956f243;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9b5f8e3dbf073841b0e6bedfabf051d7f5c14399d4d2fbe54f68d2d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a5971fc55b23db51de01e46594c31560eb2632a9a7bddcb98cc3925;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h33bef7e1e422d96351a4ae436cdc9c8e46996a7c4221bd471ad67ee5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1672e4cd8a09266a84b1571f4b826536b041004adfb7fc3aa79b812fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb98cf70fd13de5bfab13b252e406d39de4402e1949b3d02f0c2d72db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15cf3f5555885be684666d5d7732f01355ce95979db9a5096eb6baba1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h43ba098312daad1611d5fcecd5b5cf689b1528845e9fb2d46c9223b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb34c771354ce0792d473def08c44176a203ec9affcd76e4e061879b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h143fd5460bcb0e781b9f9d50b1202526b1ba02400d9d390ee480ca810;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2b65709c8aa3acd52e1b59d4a242a53f2809e5750465b95a58777e9d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6c8a2c4c1d2de96a2c20a50a57622e1e4410a4eec317b94f0d8e56cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13bb6bbbea60d69643e84a1664a9cb5310b194bf99d55ca04fef5a6fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h128b37ac584a829cc1541afa4faf9bb095b0a3cc6d5d65241714d4cca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he14207425d78af5002341e9c6d181e936acd747ab8a7c7da9431eb1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10bdf79657fac3a602e1615e0220cf0de52d41ee59b6cae1231f47737;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1308383b13afadf33c693b3d5892a1858cbd0d0a0f3ca40925a2c1e50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he68b53601e8d91af18dd5369c09645d041a9299d883dba5513ccaa0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3a29b1a097fba9e7ad91111b71669193faacf7a73a4eb97ca588d33d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4fe1bfc31a2912aab7caeed339fc45adb8de40c0266cd13e435894f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1060da94bfd224e1e8d6b9c5cc0112e545c4b0ac8e107692b9f22a0a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5035f1e4700444e98aaae50992ebc4c33c9f96dadf53c30eeb231894;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h65c8e5731eecf547241a206cb0ae29fb1382462ad5577accb16a0052;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b6d0af26d36b7ee05a165468b3d93fa4033f369de00f0f8f67e669dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1227212f950348083aa23ae0d25b5ceec7943c28f6ba9c67585981c99;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'heebab1f0b94d8c872ae4ae61d5bfd80496800ae953d66327b2f37509;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1dd8aa9e8439066c460b9d8b9dfb7d63462142dd2abc8a33d34f729ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc7a1352944f7bf52c0473c555979bc9acf684e147582ed00c1146aa1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc6168c500f188f9222694c5a819753278f71c5c625033de7729a5504;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h139832fb01b0195cd8ca6acb514cbc054aefaf566c6a1df93f9977922;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4eb5856a7215cea1b5e153b431fe76459a1e96757a96938dd58f070a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'habeabb5e23c2008988e81b047343730def5fd6e25de83395b14edeb5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd98bc001c67cb4df982022f485b0e5de0d4685a8062801113c7e30f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1500c70480af79711e831c5e6d6e41fb79c57bb6ef22db1070611b831;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e52b3b611c2563eadd0c0db66943951ec2ada8447f746b9e011c53a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h169180ea6d9c0cde77ebac2fb33b8c7a328eb6ef49fef683c7da5c45b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c03c96bce02ce4ded1008254d31038bc73fefc136265b149d887e325;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd9e49721dba366091ce0500fda1a309e0bb647d403bd497ca78bef3e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h168f1c2ce685b9b81c2aadea08e2d10c94f685a9daec51a2253ea17f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h127f1f84fb6d22dacd1da431c4f5b847759d7bedb5e923c0854e6c235;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19f7facfc6a9c3e55fb489e637672ae584bc6d0e20cbaf481b47878bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcab4dd785cf71e16ed2867e0c84857dd2f4d0ef0db957831e948c525;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h78acd4f491dbb0f62eec66675e33cdb4185e76431ca850cd28542e5b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3b42784601ce54fd9e0f9d550faee7ec90dbde917c3846432caf86e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h153d74f1a977909b2d824141a628b3518e2a7b8c9340e33fa8dc3676d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2547e09274af93f04f4f189c219fe00be255ce2653e3c50d679e16a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h96dff93dc0aad0506852991b71148dd7c3e51945add665fc3a7728c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h795687e03ae7e1ee9a8a7e4d7dd42b61b99e9b0e75db82df02295719;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d743c88cbcb0ba36bc0d6f4acd7b1e56bf9a4a482c80a8a0efe4bb5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ff077a26b631e6fcbcab51097e9493769c908e10cb3449e770831488;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c38430bbe69025b60a5bb17baa5251e19e3095296b8ef06625cdccb5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h79f7eebc9a2946f197b73ea11f36139a7803549ab0237a6ccff2c758;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h33b2df68911dac08578d49ede4cd14d35d9a4f88fa1bf161035492fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6f664be5114a490b983708122b44b9818829064a37ef8e5125a81b14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd5275089a47c5659b757be9ef00b9baf382816a7e80602c041398792;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17e2449436f4ed9ef55da1c8a595cf2b5f65f26bf8fb8a5b7c0bfb3df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d4496b7a0cec05c3f9c1b2514f888d588e5ccf2a21c4aef6127c24f5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6c4e7f3a2f95d515da994e2bc928f0c129faab4bbf2a66f94465425d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcd2baf97b3b1c944237d1851cd39f7b871fa7037a72f239cb0e4e10c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdff8fbe86d8a4a6f7b97ec67b97fe7cfcb2f825dd1d71d1b10995e00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17893833e89805e633999c8a2ea508f2f26ef32a3c2cc0f650cb9f6fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf072fc92beffcbce7817dae0c834d2d246f5ffe549c9a3a3bdf8f306;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h112e76844649a3d6b6e63cb866d49d0f162810cbb87b2293b2bc8d4af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb12fd296ac7bbb4b5ba96211212078adadda34f14066cdaf510f044f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10dfe6613a537061e9f40d8296840d6825b66df9045df9e8490b917b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbb2f52332e853689c31c33ae0da4ef65379f905fcbff6e71a8abd307;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd2ca2a132360e1facb4bcd637f6c85dcd84002ed932b9d6da2833b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b13afa1c3641bc96d9ff0728f95629a63bf44f228fea34471743a45b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h19af1b269799bb86079f383ae02bb008ff373ae39593216931804fe6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c8672b58fc9231310a87fd89ae8b5649e086d9e2e52a8320b7a57cb4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c5358f43f68ef127ae520e1b50ed10be6c9dfd993a6d4cef6a71c21c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a781be44c78ea1c2eca6371f124af18be93e07c2bea6799d57b4dd30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb29d9e9379d9587a2a957b9d0497498b331ef94317ddd8783de0ffa3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c0cce361cea8007a63b9bcda9049b72d81693d7c81380d110626aad8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he9356ec7b507e0c170cd3f1767903a54b76c01911602ecf1b2a600bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c7811f39304baccc7ad0f3a8793f1e1d9b3c1230a17802dcb4552e8a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18cf09152ac9ec224452ecff29a69c71dde1ac09cba2362b8beba99ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h125db7cdb2244a2d5c8e1c44ab4bbc720c6ee93c705375f394e189cc6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h763795a1233fde4b196d39d1a31c0584c25aedd15999bf05006c7b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h184aba4efd01038f62ff3d1d7229fe0666431c2efd45178e674c54eb4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3eac0194f66881bab78daf0ecba17a6263c078bce483ee662a2f7113;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb4fef7a8e3673f59978d7e9eadecb46b5957aef8bb1055cad9bcee17;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h122d4ccf276db9ec51bf951b735731c9a1e7f64a12cf7b04af43c9bce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1351c903867554854b96fd08050e236b3d8f5b7b26b7740adc40fbc0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h88b94de6998dc39d52ec05e231a88ccfeceb88aa99c5a54b1bc56490;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7abe7f70d341bdb9aa9346c65ddccf5bb6f43f660360fa1d75108b46;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h253f1569d7cad630b7bf8e028a6a48cbe658478e044f3d25c1308b06;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c33b04028a6eebc1868640058ed8a3ecbf56cf450b8afc1637219178;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ea318bbc0da4a075495d3d9f5d39e5e2e97806c8f5f6b56c9b511a5f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9106d3c109ea6225926c4fea500cbd7f172861d845f571278805e33f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18d0afeac39ff01d7541e99236163ac0c56eb2198c17fcafd291c5a7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e1e98952f7fbbbfe946903300578151415e53be29c4d22e21136153b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h171e61d16a2db27dbb14f03e3fe12b037471a3e67b6154e20c08a9b99;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1986dcebed0f44af96c50fdb73b8e8a0fb7ef85f9c5f55c479206dcfe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15bd4e0c860c607775286d7615a6bce16ee772a7bef2ecf4237e7664b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1fee11ec01c1e585cb3aec549ff92c95333972309c83797bdfeb75be9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h193e03201a0dc781c50deb1d1ef52047ffc621cb307fa1264a8ca36ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15e928677efdb4f615e92c2f0d5672afd8e0c0866c4563bddbb59f03f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h28b1a8b2cbbff84d7ff951a71e16c24be935db87b64b9d923684e204;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13e46afe8a2990eca190b48b46a86618c7d630f6fa696d5fbcc6b6375;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hee1a7e8d6ad3757ba4fc6f79fa371c081bbd4298388d1f7b48ece5d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc085a7ab5acb8107d623231c4df8440ce8553d2d2b3bb968afde746a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hadece281040bbfdd9b4b349a94adbda990fe17c674552f6e43717cc0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he17094b4ec1e554834f8b5fd6ccd9dea07437200fcb54ae6b23689bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h20c08dd2487d37907e1368b751071f25e3cc831f1473f65a53b21e05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1db0ca6abaa3228c03d8027e2fd3783797dbb1cc8027b3646ea34fa5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a1c097f52cf0ce2453b5527c46f3b6a4af65426a9806bc44036f1d3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14f8e30c4f135378d33d887142f96b3703b2375ad19935e885404bc15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf2b453a83a9de958d01d78f68b36712795937b23ff83bac38ade36f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h2a2fed4a0852908c15781f12ae4c26aa6dabbcaddcebd693e01a0b0f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'habc592531882f3a530dc72de170a30a2289935d94b25e3807fc7b1a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hccda32b144a3e028f9de5408de69fc5c242d8e2b8fd7649b57f2be9b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a181b4586ea02d40e397809990f046a36fb094d33e37e033523f37b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10e1dcf4f11b47d352675d7dd71d157e951eba1e39444325e52f05153;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7977c83c6c9b927dbd18ebe695db708a9b303bd139cc37252a3ca95;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h23409eedcb4e5ec93866e4a7187ad58f61904bde30148cc53055be3c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h57b79d76fef8cd7bf05ccb7df96e2218d9bd2c37cf7f1a4a3713a98a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc4b992a6844fe958b914adb8537844e1c3a3cf182b644d047bd9d14f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1383044ef5ef775192e4ee427811534123a918be6f84d762e9c4a661;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3d980fa4a94641a66dc978554a937ebb8f1726ec9a37e1cf1c602a19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1061f97b846929f964ca4f2324ec59c3390df6aea972030ed568677f2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h18bab5a8bd6d8ee17ae3f6c19c58852afd4641fe94f1d42bb51f4fadc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d0b7ce174760e4c5c5c6d1b94b44a96ef9762ad08f8e77eaa4755d79;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1313087d1bf9f396d450bb1dcc52904e43f411ba92a00b9090818d2e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a0c3387c2df4ed394ddfb2ff44f5447fde158ee3ea46794674e5507a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ca4f3a5f08c2784d2c8cf826f340a5f4b4627754d8efc665279509f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h191e9243cbf9f5f3697b1422eea56bbf59e55468b6418721b4996a2a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cd485340f9ad9c85139e293502cbdf06943472fa91e2868d0c1cbb91;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hdcfbb854779d4c3aa82c940369458f4ace087a7626554b2944ea873d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ea3cc1ca449abbd3e1b63511c584552b97191d03b3f04e467cb30b80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h117ece16d9d5a71e02a6c429f801e5fbfc132d1554a98e29da193da8a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ca5cb6572601d61a921adfbcf4d7e01a8b51bf6bf9c66bf34cfd545c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h99093972549b9e2d76313db381754b6609e2b9d371dceddeff788c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h769cf2f9dbf37070df50ec9ed29640ffdb84ceb52a733978beb91f7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10a6de1d8f42e6f3e27b17ef630d1391c4d50270f8aec96d0397d8cda;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h29c935e2540a27b2194268a0a0af8a0bdbab9ed28408a907f1559913;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h86abc8c678150e7fa6eb3fbc1cd401e4363f0c9bb4f7be68650df9ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8cec90661852d2133116ba737ac511c38f452c61d6c412c86ae09c51;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h451fd94c26c4bdad80a28170329485d782c996af6f17d67dbb8ae35d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf7c27760df2cb433163461d0678541ec81e46944d97491f7a8fd8f27;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h177ea8fbe6807a8b54d4bcc04335591d9efde989402560a6f96c5f22e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7024b61c66e58a6e6e711250f003ca87f2db64a2de03d9d9d82ec815;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17442ad047fc88cd33278f985cce3e049542125c40de607181837eda;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8b41b6391228cdcd499877c9c5edc99108e8caec9c89863b79f72305;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16c7e0b658ced7b7b19a877f4fac500d61ae2cac749f6cd31568b24c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a1d991de5106d56e4f15f131ee9f3f795e28cf8e9729be3965eb37dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h93f7731db3f5c3fcb68ce87af64a193108c2931a9e379c21579d3f08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15529e3a8cd191ccb957cccb3f5778342b9a495018706fe140a38850b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf590b62c322d9ebd290b6687f9ea615cdc660cfef7839566845d0945;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1360fdc170577fb0ebaa8e309b34ee0bff247c429334e0f2d4d04aa95;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hae75be50672655a8e81c248703f4419ebbcd9e0d74213779f8d92a0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1412ac9adbe7c886fed6f3f21b872c7ddfccd06ad2d55c56dcaecedcf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c73c015ba54dc494e9d2e60be0d35680be7dc7b49a9faa07146a5921;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10dd4ba95b788e183660bde2e88b713a5ed3497b951abeb52d34a315f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h111cdc233287139caf6525681c32a7afab78f2f7dd2d027804b036093;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hcae7d8f4aad06b8ec1bf453423b08ecedc967ba502a846a248d2f783;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3732a1f93df8033093ef3bd930a80b570d5765a5334b8f43efff0967;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hffa004d848f0af80fa57b8f7468b37eff4da2be03f8594366aeb0cfa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3e4297ba31d5f1333f2797f7537809191b82733c720e88b06ad0e8c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h764bd0f8949fb0389ef53ff4b29135f7642347a02cf275bc1a5173f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef8921e5748aed4801db5d65a00235bb3d92c37fbc01fda861d32e6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14ed0381186b52213564e08e4a67f204b4b873b36b406c49e71fd6d88;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h95a4a37aea5a9c3d78a62dbfa9477f685d0d8f5a0c02cf4acd9ada08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11116140fc5b28e66e61764a285ddfcb48fca0d8cb3252d0678b7f0cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h166c716766c36bc0dc3b393dcf0b255c9dbac6b5895c586a27b0a9449;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h120d0da97e00b7fae44d15636b22c33b49fce56ece1d1d1cf399c9604;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hee3d22a35dd642078c74055af7c37e669f73d78a96aba96b73379b65;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h35098038ca98cd73d032531beb667d7e138b245b730ef59a4a6135f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hec3d65a529ead6d2f18bebc94d021463f785d5fbda216fcaa20dc162;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ca2e6db027611d48040509dd2093dee893bb4ea11065fde8fd92bc29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1490ad455588c12be932ae65858e45270f92c50b6dbfeeaa91cfe09bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd2bd818f9ea18b3a372aae7043918088a1b96e618aede410b065209e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h93499e6c5d4b5ce23147ec27e0f3682b111e58cea44156df3bc65965;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1719af891d54348141ac99d07117ced18fbdb2afffdbf732f4db13d3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hddec8c25d77d291ff9dc0f4ac19748b12eaf367fddc9c6b63c5f1265;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8265bf6094fd08e3cb060b93e53de8594f6a5b3ed10dbc30c689b39b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1963f3aca2b27135ad1a0150308f3e9f6456fa58448f6a072cd7f1e87;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h617446b2d3c675b678432bb2cfe56e60c2a2a02f9b02b39d583632e7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hea2be3139b3ee825b89e522fbbcac00abb19157d11073cf1feba5df7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b681c47c3519af5fbe8ee4b9e894da400809491c728a38342ffc9469;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14dddfa0e292b7d02a33f643ed991c8b6161fcfb4d081e1cb50b09d4e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4520c14492aa03607bfbfb6af95f6d687dee51480a748e4043589489;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc0a552389c4da6261b3217203aff24967a6812a4bfed4c3b09020a3d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1312806def615f4cbaca5acbebf719bb5dfa6111eed40d002d5e14414;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1420a2a8f1442ea5063d0cabd7222dac5ee907ed2897eee2dbf35582;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8b1fcdcc69c0ff3b3afaa16d5c95e6c934b7e9c59207e88473f784ef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h14d7352b8793f098a302f7da79faa9c0ffb66807a64fc054a514eda2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hb407d3a39558e34d713a01612a93487b13544ee44d1ed9df7741e176;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h172c3950ca99028d51f8f486c089bf4ca7804a04514266f4a8cc08763;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1316f0d6182d2dd8d85b2143351fe7b66ea4a18c93f4aaf1633518453;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1478387724ec0c87129251d01685e33bade3d952e0afa7057405aba4d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1de0c7c27ca359190127787282f6d12fbd66da9e6bb5f5113b86e4943;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d63f99d149c138c05510b966c49a7c13c6b0f9a8e8ddac7c4fae3c14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16d91049d9fef95301561a2a1a39e861d0740b989a0bf61216a8462f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ef8b4bb1f4ff77c765cae695d09969d0cee4e46bcb3f3ce1b1f5220c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8de32c76f3945609e777ff406f930be3d00a3b1e0a742a0916a8895f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e4dc564420271518f54ee7c7a5863a3803d221f02fc1ddbc84e625f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he6e339781c334d09b77b2d55738f40d980921e562643744e62ee22d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9ed14570f5a6971afb217d08dde7904fbd227624727391132fa4e8b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b89f66b3c5f2d30ee43f6fbebc25b7ef5b40e87e36cd5602d1054bd0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15072a1d51675569a380fff099b2d9ab041d274182c90b1cb652bdde7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hf2c47d4f1838bf7918561d6ad76c9071606394d809667e1a3031a087;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1d2f8c99a69b4a9e99b9f22bd3e3e264f22ad59cad41518cd974dc80c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha42ab6f1c5731c39b5f2847d0c8225dd1ad3515072111721935b507c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f425ba5e250401b1ef5bf2947e9f9c2651b101d7c09530cdc9278d48;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h155ebd70c4e930123f99b34901574be0e5e2a622af4ad2e7040d28b50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1f99d3e45190defb53c526db99b0ae88035452a5b4d4b83538713af7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'he7a276309d30396bb366a91242dba2d17fb0f4bd8c9492bc9b02369d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h994258cabdef23fa8f84757012234a90d30ff7b2371dfcd6457783f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c98ea9856466de14709fb179a29e0435e52a33841c42200bb5a79ccb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17e76c9ca154355ac420830cd84d58258b17ee5ad6346f4aafd213811;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10aeb4f6d3cf1bebafe129db8797601c09ed7b7cec874b514a59842d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3e407bcf0b3d7a60a10da1f85ff9ba48a5cacb40bb05440aea193460;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h111bfbdb3c36d605dfe90912a5a7b8c28cf7feadaccf3ad5a0ce1e8c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1e2ce4a356d7d9b6dda8c8a63f93b46fd07836086725996dd65ae5b80;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h125378fe56f0b410914a383b8ebcfc9a81e21b8cf917090b7bfef9be3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h9c5d7e9db4c6f5f30f6a594f8868c7eadb0c5899a7c067e9336b8992;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1a87d9e6e2b9b78e41506ffd746d5076e455d18d52dc88990e5700105;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h17ca85c50121afcb4bff2277225a58759f88f858ab4b46e1f81d5c29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h286e9aef33126d97f233664a878aa71961f6bf0e6560adfff71f64e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7f72a4a6d28972c4528ee7a1158672f17a5fabdc5b27e1f9d5b4c568;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h16ee6028b7002d5c5fc277bd09eda76836628e0371f5f8065414deb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd37eeaedea67010b1490cb8115a19db29f6b01403a7ad632f31acd69;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc6e8267bcadcfcf630882cba72769e8076b33e85e97e853cf7f04979;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h388ee4229d980a8e808ae5495cfd9f495f290f62d68bc7914caaeeae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h155e30f7fef9395b342c9c844676efa5bcd61d52870ab3c5dc973f18b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6f6eccdad36f342c49cd56b7c4c8de526dd719aacb3111029bc3b86c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1bdab81b67cdc400c7435c774d0984f516f321b8d866e77da7eb4cbf5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h15f3f18b3dbf9f342dd055f12f4fb34c38d6115b0e749ecae39669c12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ac7fb45c9cd8bf86c0812d6a92dc8546e3cf8cef184805de0ad8f9b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h828673a3b92f3db66287adbbd11cb79c93990396b6a7d796d35b2298;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10fc241a18c92879aeb485190f2e622133411472f044871d3115f99b2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h183e6a2e12d5e90bc56a226b946c02209a785308dd7df504bae86ff4a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h109e197d6b3c7c144ac837788893ed8e76d9cb1d29af87c7d46d64384;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h787f86da1c04ba18ddf362d7254fe0d523aa519890817ed98c2937f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'ha97d37543e00db6792da74d5292ee88208199e9a9d5cd7be240e80b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h11b4172e6599b0ec4b64e9e6f2a5d0d3375e2db24080ce67b93071b68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h186b3ece23caf158441cc63e2e83ae9fc94e975da95da1237adfed46c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c849e08841e719f286bcd26c3f98b123d1abbf8d7f65990fd1d55259;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ba0b5973d21bacf1f2c8a0d0f00b09639740dd98b767d026e31a417f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1190aa1c94f2e12b192151c72b8652aff0ccd5713a962813da7ec9024;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hba385f6efe781aab9a31a00bfd796967f30e78416affc7316f4dc7b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ff6de0ba3b262e75f684cad4302178f522753e8c57b0ab70d28d7fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h13bd490df0d060dc3430f627fb06182ad10f253cdfd9c942551b5a903;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1c9f2248e258727c2c6f466e45095cb42294f950943ed403d2c0545f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h8aa338229f6856387de794ba2453c0056b4c52a721012b5c85a83ef6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h26ea48f65c91147775b4468556c73882d135bf22d1abad8ee9b33e94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hc37df9cbfdc769ec64f3231b557e5cf6e42eaa5ba82fb92b4b3682bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1cc5609b6bdb64dcb7ffeb113b17febf37750185901f4c033a79e424d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h973f819494e24d49828f59f6fa382128fa249e8091867eddcdcaf58f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h39ebf0d580635f18f7aec6f74d6d994d28d1772e1d3b26e8333393a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ad2fdda9eaac0b53fb25726799bf66eb974180eb18058ef38f40a470;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1b4a5d12fe205268b05de733a3ef43618a43184c550dbd8eec18a103f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h936dcd627f8c5c52d68dbe5d8f06dd0ea5c9ffa1aa4c8ed6b9a419a9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1ca44402470dc3edfb5dc1fbd875c722ab00ad656a2d61f5209d6d6bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h10d34d61c7c7cf7e972f1a9581a7fb93c256b6e9748e2bf7fea41db6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h1430783d17c5cc47353e2398fe2c8b4e143d806bfb990a656f422b88d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h56e236c895eed3d1ac5d952fd3e7132893fc212c100337fc69e4a126;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h5f2c114f7d9037e812a183d9e25ca6d359200802c01851e74d82320d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hbb4534b57996b86eb101304c9456dc82c79e62407c0829e955d59752;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd0034d6072e3f0d894a23bff39d9b13b98a0d3bfdf4263e3bbd522e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h115ef141fccbffa27f1b4b26f506d4cebd31a4bd114405d80dc8df10b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'hd6a0571e65b4711f3838853ee5cdc33b7b0decdadb751f5378698b02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h7a2fcb485902ffa75a76a2b976183d1768f25b9340ed88ff4b3d4c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h12b98c26ce59e7ec0f878b00daa42c679f071aae3b40aa15a4df10088;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h3c134bcfb705abf45fcc9af31957ec0cacf59dd4a87e7dcbcb03e097;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h4a54ff6c614b60ae8d64df625b8e18eeca31e273151c7d199a7d4886;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h6ca6b8dddfa428a0abd257f10d48e402a4d6cdf17520f9f911a8fccc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 225'h836dd7b4c3a21a7580fdbb620e8320db5a2737c3a111da18cbf30262;
        #1
        $finish();
    end
endmodule
