module testbench();
    reg [29:0] src0;
    reg [29:0] src1;
    reg [29:0] src2;
    reg [29:0] src3;
    reg [29:0] src4;
    reg [29:0] src5;
    reg [29:0] src6;
    reg [29:0] src7;
    reg [29:0] src8;
    reg [29:0] src9;
    reg [29:0] src10;
    reg [29:0] src11;
    reg [29:0] src12;
    reg [29:0] src13;
    reg [29:0] src14;
    reg [29:0] src15;
    reg [29:0] src16;
    reg [29:0] src17;
    reg [29:0] src18;
    reg [29:0] src19;
    reg [29:0] src20;
    reg [29:0] src21;
    reg [29:0] src22;
    reg [29:0] src23;
    reg [29:0] src24;
    reg [29:0] src25;
    reg [29:0] src26;
    reg [29:0] src27;
    reg [29:0] src28;
    reg [29:0] src29;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [34:0] srcsum;
    wire [34:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71a5eb86fb8cc17678d634ffc6d041886ccdd27220d9e15b402d65da0152fc8b5e54d8e2169d61fa8e3ebd08216ca846dea58ee9773896bac7c3cc80ebdcbd689ae42f1f6264e202e31a8dd3733db01bcda6bdba64863d7ca2996287691f9998c6b6aa28128b843a54de1068a058b317b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23d0752040c3f87290e63a6a459cb014b71a8abafe0c32e3b351b5fd96f53d26014ffc9e255b0f155e7a895b690c9264e9723f0bacbbbb40a1bcc60cfbbd0b0af88a38f217d40011f81fa1ac42ce6d8052c2a5fa0b1886d6bb5c3a56e0cc15d573f0a6e526865528d709107178919fdc5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c2ea928c96bdf4a8a780e2d253b7d69294c2b3cf181dec093571c813e95b9ca5f0dac6509f50e30b905ad7553e8ff9d44311fc3546fec08de2d7a5501a42515dde56d51a557ee1f7fe0b834a68682ae795059bac4e22ad556cdd964fa1f11c6a3a3df9263ee78ff7bf4b177289d4a351;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4875f4d672398b4eb2a8ea0d54746141542b3155a7711366c9e5bb1ec9fae5eddce36cedeb590eac22495f1f12c912401b7b7c7372c07ca2acaa45e791f4c65ab24877fdf7614b805468a031c13678f072a3fcdd301306d2c5d3272d1fa25fb06fda697dde5c6ae340cb9a4fee4f03266;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe780b7426f569df681b8ea7b6d9b0fd9af286df1fe6156b2222791fb920e61296a55e79ce84207794042f87c39c4e1f1e036165055b1cb3e48f11e024729be2864a87336925883772ef94e71413d6b71297f70efa340141213451df5080b9b7386f6eebe714d4189fe856216d01e6639;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he266bc382ac35a781212624350fc61430b2c22fa2e9c53cb4aabfa125679fd014564c00ba7bc220cfb1083dcde5f8c4eaf49c5eeebe6a7315d85ca738019ce0bcdec5bb8f9e5f29eaafd2216eea5760a6d06d20591b8f0408d03e24d420e3c7a5b3aa2ce99c414e06664a04ff5ac3df67;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcf7d7100329439a7c8e618236601d7cf9dd81f464e4c2b8421738bac23691be3945d019c12f7d85e2d16646623ee87ea6850b1f53d4be96862a6e82b1cd5a1f8671f07f5dd3f0d37f1003f544190f42aa8f8ab6cc33535a86ad7ba7d283d8a26e64eba39206e607cda4d0b9d86dc9213;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc289e78be7c4a2afdf45babf9002bd3afa0ce252c897c417d39390a796734989af761d9297d3426c14e22133e378efd6a8910cf6992814be73f8837b9bc73fed3130104dfd5af749c50ced93afb6e3f6179e4376f525224490abe4086e83514d5ddcb83320ece49ce3fabe5f2eb49cb4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47a9d173c93c14818ea7b075720e4db011e68218a118c2eac950b053295675630170646aaf3ed230f68ee0262a4e6a2e4ac9897396763869cb5190e4cf410cdce88a3827b0e188fab509c789eca26b9e87c58c9a5f665abc4144a2efe602b492c6843c580b4e60c5156defaf40ed684e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdedc61e0a2b19295bc415cbec22f4c7c0a5c49ef19855dd3d1a48c90812b2fb9337f99f160ce7d4b50425c632972bb75625ca07475b822ad82629db3fd5be5a0f90c3bad9085d2a617042dabc3a90d96c1f7408fc0cc85349ce33636702958c0eb231b11f4faadc91dac22df966a54f0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f2defa43b54542b85692f618dc7c6ccac12415b19e5f3ce3acd210c779c0f29b0db4a924492264e9a5f3210d5f4c75757142787358c538ff0617944104dcc4a62693c98fb4f00d98e4d334d546efd169fdf6bc2fbdffd87161fbf3b358122ecbed8763878fe89f02fe7a6399f0ddcce2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h521853ccadfbe2f344315e106283659cad2b5bd32e2fcb29136136c2e391d3c6a616e02c608156b80f82036e883c8c76d34a33506ee7347b218a684cda0f78c3758eab2cb40475b86ee2e1e0f5247c7cafdccf8ed2ebb6f9d6695048a2d2107d05e3af4751ee428eefe580aca8698ede3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c85711a483d7487737957be72ee79d5a2b9706db62667424ba63f4dee36ebeebe5c09dc6c723b4df77c84e6718511c869db026a45b30048a53781c036de98af1604ecfc4b4b96d6168c28cc28a2282749df2f678bb7a1dea86e6b7642b0202cae04c1194d095ebf742589579ca43260d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f8dedb91fd862b70ae0d9f3f0621f101d5ac287fd875157ba0426e8166dd20216d131f371045893d2256a22ac77161ced8365824c4bee074b946b12973d41b97f48df34c4f6336c93faa43cb61598f4f3ce1281ad552324edd1a659380f1023f01b7e20b57baac76f99f75b2c0fee0dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had9b0e515dd2e24c2aaa693e9236e26f7fa671db812d65fed4a90cee2cd766761c9c575bbeb5f71517ca8cc2edd1118a0e61214d18d587e73af911b90016029b666c9d7da09c33e83517e0a1e7b3e037728c6163ae7000f7899036aa038b2de56ad66feea05631ddfd8a388646487c502;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4806de2b75e765c67445defd42cbfa85dc3376c837fa48d8dbaa40ea807b57be46e875cd967ca9e843bcde00f4da5d991cee97deedf0a2ca0e752e33fc16157f8fb1f37b0e0b91c47ffe596a8fc587046d5b60ce9a7f1aca7a388975a404c567fb8c35d5fdb6cd8bfe7800c679677ec3e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8b8c048911b9f222d0a26f8c7ea60d9c2e92be6b9fc88e2b2d9f3b780523653af8ee0114a1a0fb73e0744c913358cc33ac61b49d94b6a7db990d80b53e38ecddf6e4f1c288e2273da8e4ebe4b892229a4ff6fc5cea3b5c880fc4763cb91b002138154523d6c2196aabf123c8a5415fc6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h138b329296cf10d60ddda9cd90a9e82bc70b7e633359e0588b292852b063aa5c5a64414026d30af9dcaaa203062c294329bdac03d405c0ecd2cdbc71e829e5bfd5ee8aad875b9047cdbcf9a4bd49fa90db355b5dd2acc5eff0e8ffdded41ebcf11ac219b92cd2d0022b933bcacf25d37a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1159b49c09aaeced2af4197895b121eae1752b41d54987e25891d408acaa9c18b500c48d2d837e8efb8f5740c3a480e22b114cb16ad1591065f1955e11ad5d84cee3e5bee183ce73cc7428b3685bb52956faefd727a99b7c30ac207c1f47bd96dcf91a331618414d742479c513eb6c6a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h988826fde244764491683bb7ed59fc2e3747443d09d0ded274ba39a01499fdfdc26c91a146796ad4c2a4aa65cbbb2e9ec3072effe8da4d52442eace70e672ff550b2d05c761a369232fe01cb6902af051da916684a08d67f2dd2435beec148825acb62908c2394db656844579623888b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc1842dcfafacb67110788be6b4e9a89604108890fa0675bafed7c20d2942a58ddafec9ccfd901d0435253604208bc0ddf53958085864dd27d7afe83266701bd2618ad691334b39e9d9d045d1aff588e133bcaa4d98fd78cb47cad9cbaead2fd04f1c692b6a4571192fe6c50445344f90;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e77581d0a0dafeed7f0697cf628bb28bbebb998e8db2c28d675e021449a3dfb666f3e0993e09e495cf8c9d82f5d1f6b37c338f9af813f4f94b5427842e8107d1b9ac53b5789328b89f2b4fe2c6e3842cec32810fdbab1efdf0552b770e0ef9657cf338e3ec2d6fb383cd446bb9eb94b6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51d26da112ecef206b74e4b49b74f0aa7bf8a96e9712886a79a4a74eccdf8a9db1a94debda55ed013dc1adcf5042b9dfaef711ddde7379a41ed34f65bb28dc85455b4e168a2bf84a5ffe24bf339eba8746e8901c73d19b4101018cd12ec410db31773d7f1224c2fbd805af861efcefd1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf25f06b4f7a36220e6aaa4606c7d51b38bbce5d367ca3be6c7c27c4d88649b5ed717a7623cc97a8ea49b425cd52f046f0997256fdb79cbda90f85f23889c850cea676b377a85277e5c86dbe2c16354576746f04535e37c1caee45fbd8a656cc0771fbcd434548f3665dc97bc81bcf8aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5ff6239e1410dfc4a0e0925760ce54376f6006169e0e745aeb88ea3e720911d6ac0e0d191a0eeb38e3eae0d4f7ed778263525dd0f8b195afa4b3f76daaed4f1f0226f1eccacd47d34eb09f0772e987a3fa4f644500cf6748257ac22e62da154ecf512561ac44a06fcd2c0f88abae4bb7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4343f777089d7e95b9a6d87de9f4377138d8bdf322b54d00419fc2b28a925405265a02d317d16ddd8564a0723e204acc15dc6c1c0445a2ee26f18a5020e2ab6b874112dc209bfb0ee701b2effb91a85d44f6d02d041a69ff69b1d3c591fe90462fdea057830d6eea986d07063c7cc39c5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1610775d3e1bd3b4c7c3d96ca504a2c8e14bacf681be8f23a6b8d05d8413896f1240e454756850f71440a0247893db53da41e9c7cb57ab11b6ab23932782e71eacf2f324ab1d7c9fdcdc5fabf515147804ce2e6ffaf06607d0d5a382c1690ec6e294c12b2500654c9af8ea91da60a7ce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h615c433eb9fd670eacf6c389d02e0d732b21397c30fa8cb1f4a62455b08a3f84363746e2542933198ca2441cdfbae65c2a2b2ed76a6b934c84d0cfaf4e578612d680ff0d5dad2e19b17148f2972d3455aaac88cc44e084e486ce9558a0e263158cf06f79c9bc2eb1aee9dbc0725e68bb5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a94f770c6b5a03858a0a601392dbefc77be78a232e58d0f6839fde57bd88dd46c9fe70e3e9f7e0e7d3578f6bfd17d99dc1ad227ba3394a7c1e99434ca58c64a4ed322bf6b5e6c1303fd191166b82938e2a58a8b42ebbb3aecceb1abd4bce94cb8652987d592afc10555660a08cfe9906;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f23fd51033abfbe408d955f55f26b2e4f94f6599775573b4fc031aa7d87c35a943296019d502fdb171bc872107fa252b4b11b0fd2cc86428457123e22d28e44c5324e0d2c2ff1459a173eab02e689f38b65eb2008c9962e91c4d22548f4bdddde8816c9cfdc746683ee422504195f64a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7cbbfaa8b7e57de52122faa4a9858215086a32f686693cfa0c58bd272beebe898acc9a56e3d7aff6d993be9a059e9c6d62b3b9a2cba14d9d779831fb39eb58c7b881d83e917dccbcda9d6ecc62ddbf7f03f4616e2790e0e3ed972bb00f33edd4202a73391ed130223d70856dbf24accd4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfed304d504dcab20d01da1a8be00cf16b36b2b94ec10fe181b593b6a293aea28c6b23a26f5e14e289489ca52c72376a54d2fffc78089de7464ee6779c471d121bc704931dcfbd5329f74b4e537c3ba25bb00d857b48c6be4cb0257e2d0972fc199cb0cc6f054f88377207b1a929ce55d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5a4ba82dbbb2f99716daa7f804f8ed1e538bd000faba91d48ecfd309a78e6fa78f82d9eb57d3b6ca036735feb0df41b60da33e2d3d0189a27ad8d90d4c71de91424e1a0152a16ae631b709e57776b9769ee67a2fe3f8159d78efa68cfeb74b8c999a6ee49e05df6b88cb8765286057bf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8b3f8a3dfd2a29f6602f41620df36c8d006a3e9bd612400222c04b9d6df545b88fd422d59cf20b508d1bce0a0757161d584a87416ce5d15f8b104def1334fbde8de1583cf3f093fbb1a2d74f50f30764a39f2e61d79a01e60037c6d4b693caf98723736f01404dc6ad4b25abe883478b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3bac1c5b0da75d7ccfecd0c71a3837a2b9f2468b26dc4929a9589312330fc7e3ef2ede4f09349828e8dbc7c05f65afed0cc135eb7dd78876631ba4edebdefe30091d60c6b49c0be649c71790e0ed43b97302f62a0a645bdcdc5abd79ea4595c0d571a160dfb1d7252c2a7371b3021588;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h690cce07225ba902735c1a6cc3fd1f7fac79fe57ce259d49b419577f7f7933cd1a40a38baf5ff0757be3dc1c88d9905b86bb1ab1443ccbb56311d07ca22c3dbfd1613c95a947cc3b0b720263635346144c02269ed43e4693640fe1ca250abcb0265bb094a9f2747dff501435ee60643b0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h492af300a4c160c7a86a7b8eebcbe89b849221f4e1cc1d36bff09df5ac0f3a282c4e2f3a889be9d68cd05f5a1b3ec458004e89f08922d87f4ab87c4e1ea5f9cbae1beae44410380b1ce4816f2478634ebed74b0922be956b09cead5071f90b06984e00ce24d5b93b9f31f11d68be6065e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb11e7f16136ede1c1317e8728fe41bf28bd2933ad5f022bc00021fc3ca91bb46ad9fe28d6d676c77e6e6bb74837f3dd0519d2d25fbda96cef315c0324174de4f43a16256fd84d803c7c67582c1fcaaecaac523ed591314b0307523da96fbab5a5a6360cf2e570b7830265874dc5ad0ec3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd7d891fe5e1937f71c5bf9e77260321f8b3ea91c88b69f151e05f4599a46a9f1207f84877a1e1ba6306a35f92f2bd9ab40e574bca01abe2223596c853ae51d3e06eccd8cdc916aec046e74a1ab3b6c898f5d33a7c762e5c8cd254ff60acd5502d16315098cb6552ca016429a2fe535f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6259f65d9c12f5d1b15990c27272811f667866748d5f784fa7b646bde3d7de243f67867d9624212cc49a64fc04991bec1b759c1647b9fb9182eab902825d8a5e93b500f6d7c90fbfd38afd3158e7725e386caff028245cf829a24e8b69af1c85a59c5f9b9670c33bdebbe3111ab5e94e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a796ede8a62ae9f7ffc93dd2ea9e2b0b4ce824a204cc542505ddde4973ebda61db56d1225f9147cf4af894b87a7fcd2821aeb610e1646971b8826dc11f598049d7ad7279abdfb813b1da41efc600f21dff86bf3afac954b4e5dacfebc9e2e41ee8fc0f9d6e383a21c14f12947eb2b5d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h723796e80299e5535d147925311a0cb9f8bd88f7cd9cf65eae2c370e6ad2ff93da4109263eb781515108e4279ac5297d763609d0e5bb8934697d80a6fd74b95dc944a9494801dba34d56fce5af518df96d958f95dfd94bc44ea660ff9a464e58e5fd13bbff13121f26f8208f15d7ee67e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c2f6416010fc20c924221e24d8d02d881501c0929ac51ea2c98bb3cd14b0f46de4dc3d6d60752b2b9ebd2146133260e9593a6d6e2a6b612c285cbedc07834553cb0866b65a86dce052fa33384fda9f94041ff1dc8b739c99ec9123d4b6322c98208266c122ef02d80323440deb9301df;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe6764f6973335165684d206765aab38568a58c4e8e2e54295a30e6fbffdac4ee499b1cc262262401bb94ef16c7a18db5c6bece03f77f940db40af3ee2b125e5d62dd093443b53b782a2a25b2e310749d3a7d5774cc06a04ea7818926e8f90a62ea9bb06dc7e442719c14bb8344980859;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3601b6b1884cd27c48e61dc2b67620bf3853d108a8e2d52c6d72162f17b548b5ea7c016e6c6fa9d191a58e07d51ccfa31eae6cf16b8ce1d980641652f891279f935e726cbd6d1d21ce1c53b3ce92eb88d9ee876ff2d4f369506432a96c5ff6a064fb402facd156828ee7d83d7b4548b07;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7cec055dc7b6c953ea2cd88c55d3d6d819383f7baad174fb4bda1dd5b4c7fd7a0660731397aecdb5527133ba27a29fb614bb6c306f72d023aee4b1a607c7af52fded70afacf57a1f28ff642fda4f060a2c342509a22bd1daecd41f24df1a511e2deae69cd7f1881850876ce43cb70624;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed3fd68bc196198bb6732d34c62f9b685b4d9509ff0fc2e117392c9741111063eba54795442f185ab4d85c93b5ed2d98ccebc4dc33b0288fce1af718dc7f8c72044d8a4b75c6b94fcbda8111500cb9ac41f5187f0781fe9dbcb6f475d301d908a751abf16cab2a998fc7177845fc16466;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4e7e3fa80aa3aaf27e248c59c178a41cf2e7f599b2afce75351da665363fda7190a6cdb8062a35713e2681794be8daf58f580cd696e6ba74d33932926482befe0a560521247af7f5586546f1be628e4bd573fcdeff1e1d2a77813d7f3f45108467514c895cd948fab5baa6db6d05999a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h799758edfaa7aa34010a42e33fa9df3e05e1670a29350b927a7eabbf407a7690b7cfe9afa5162624770e2487e91dfdbdb7ab15e1de31d3fba83b298e8d99ed1410b438fc6c18d1783c6a0f17bb1f47e0b67bb784629b089b6dad8f2a9d512cad3bac8979c9b750189b36ce2a7fa72044a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92ee4fdd1db44520eb87cc1c805fc5a7feac8ce5c549fae802e0d1c7d41c1af2059470db06da93701aa58b7ab88fb853450e76e78a3eef0f06bf7dc32831f61463f4b84e40eb41f23df7c46340eab32db0790be55128257ae84d2125281fac0f5f0afa592e8508fb952c99f3558988ed2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h717950af49419edbdbe62fed5a69d3c1de2467eb8c7868d686a5102ab48ba2d867091e8571f1dc6d4d551f93efeedd322cb40824fb4e60a388c7f42f9c0deef868a62ef28db7f7787e14f90cf8c4a7f1dac7f30574e94f3dfe1d58ec3b9f6bd754bd3f982376f7563ca52d0fa7c12e40a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d432f389a729748058bbd40881ab8f34896c31c37c0a7403afe96ec77fc2e50bc508f4bb8d4fa7d2dfb4a812b06b8071e8a6e092442b85495560f9e387d3390b3dc74f49de2344d1ab8f01b11e717e0cbf2e32576dcfbed876c4d19eba8c8539ba7ddad09cf979768d6b70e566a05aca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf28fe2ba963b34bf0aadd1d8f30e30ebe418711821d623ffb9a237d5af3c1ea7384b17b925e7313301275eac2ad0d5a12ea6deaf8fde9aa6f640b4d1f27705c075a73f5a97c640de4324ce373e857e8d82816d21f8b84569ea689bdcbb9a72e4826398f2d6a92edbaf3f7829d2a550354;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6aeca74102a52fd3007a7a60ea81eda3681c7ff1b8bcdbbb4ec567fd0aa97a34280dff3dd6d47e47e0f99fdc61dd70a40b1911cd4f0e19dc05df53c05dc4678aefea98b42fcd322c0a1bd5ac22a0a85ed01af7b4db0c353b92074be69c396ebcf9c112c87bc8592f83f2151efbbf4d6dc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e084575c0b727cf0dd9f11d30b8883826caac47efb682d2bfd505f64ef5bc43534598ceb472742f0d01928db4947affc8b3b8a0925540686b194a64643d24a20053542f1cff540f6f72557d41d5a9df0eebcb84a040bfc226c2c79f20e01a31c98572e5aa4a75342bfcc0ecf976810bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48e9a40ff1537802c0a11b2a3591106732b4005732a4aba1af5e08e5ecfeccd19a44e2914f67ced39e2f801d7e2db48f777acb4763b7ced2a6491beccc1e9f4b8be410de26fa630f8a9d1fa55a7fd01629a32c941d4bceb3ba0dc737f2e8b66a3afd468dfcf9e2d51feea56a71b46dd26;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73e92f9b093f8004c16aab8a7442db33591b4191e7dac9579fc7660244b82a773d5ca505a5730086daca83918b0b2433708555ceae20187674a3ad7847cc6de892557a70757db96252782107b1103ec3ae90e8426f64ddb607dcbea0a528750a474d3f834dbb2a21e419db6ff33613876;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32efba9874ccc6377a7fa6709c3c27651d4741140be2e110aaae3d207f3fa48650a75449e0abe3fb146f8699fa5bcbae50d541295ff0d4bc0f8d32d88628f37ee98c194aac53e69757ff10c4a5f350d155df32a818322f438c7110b7d4402bb316981144a1bcb620c017e1fad1dcc7aa9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1608bae2735a46f21836f795f7241d1e960653efcb5ea45a9c73da19876e15761999d12a95539c68844c3f3a9ee5f12fe63a6b6017b78a0a473df5c0059a504395a912c07d20357fadf808320d3b4a952aaf063c8bc78debe9911ebf5dceb82d186e1ace6cafd545965100a9a11b4765a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc7dd15f4f492947a2f43b04b1cc18e0b6fbe74d67fa673e242ee5210a26c6685f1f8091fdc3f48e127dfddb0419ef59feecd9b8713876265b8da5c44afacc178f5cb61982179bd64a981034efc7665bfb9f22a6dd0013af06c50de05c36aaebb0abd39262c417f6ceeff1a99a869b828;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c16d06860e9023551cb072d74a03dc74ab4ce29fb30725422b93bf85e502591fb44346dbd39007a06bde3106c98f2bd96e2bad8b75907222f5eeb3db33039a12ef2eace1938a2a6dbe05f3097fcb6345efdb88884e2c847639e7a638d10d87df11706ecad0d433f2b6c9f5deba94d982;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12cef33486b03c0dd356e640a718590bc3fe1350779b75886b621b4b26e0cf0030147cb25d8d223d89463d0b8898944975d65bcbef3c3e0bc3b997bbfd36a8bccba3d4510bba186e8bc866fcb65c48ec478a251005f560199888f800b8492e0c56b9cb5dbb45f53a4cbd9e3ab0f09c4f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc596c903a8ef57d507738813772ad5fc80ec19e2fcfe89a6db9a1e81f87d35d73aa15c81a0a0d0dbbaa997f74f768db99398b5a351c92324d9c5d1ebef0f2d99284f199b9cc13e9d29c2d245e15b290c93a90d8ec173725e93f4f601f8dd0913bf7e1a57915070bb0121206783cafdd59;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4788bd7071d660a84ed689a0ee76ed3855eb997b18760d97ba8f7d70a306a6b2ef52b1987bf85a28401ec0377423bb7581fb4c88b9f4230f5d3f5209fbc8f768aa6c15e1cb0dff9337820fd68128e980500693d6ea4420644840ff5c81498d07bfe493b8511c4d766ced9a4d97e7d893e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e22e38961ed9af226cc94a7e9373dd430af5eb7c11bf09d4c8b2f58a273cd0a5a6189ccc63c6ba471c0b958a4fff03c0d3e291da2406d4b4b98a52d22036c5759f97af53f1d1b7847efe58863932ab82b248037b800f917a98100c85c27fc9796e5bcbc6c8b986a5d88c4bed89e77d7b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf86c56cc9f6e3daff1e8b57d52ab5d24d1abb10555a83031272cb733d91dbf7ea90fe387e4a0cd87648e82be4e150bc20a84be00f44ab5531a2f12717dd5875095b543f30a477be4994bacf26cb5a9e14ef14b9e25bc1d1382711e387c1c3921ac4d7f0ff238d97c76ab4db9be38b13aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a7d3954bc546425252a2b1eb1ea4b0a1e1f3f6db3409ac6c67a9eef4fdb191dce96763f9edc3fa6c5b84742f14d259b28d7a77ddfc8219962a366ff1f9b728057f4c44f2edfd897e2e66e4c1cc3a4d0391bc103427d516fce54ee687a83d795521b1ced9987097817d36fb0d1af52c53;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb010fe25f9809b94c32fa7717d8adfcfc561775d5be2c891e61a0f3a496779e9df316cd0fa9a2635260aff4b8307ac68034538979ed8875e270afaef6216187db630fea9016983935239adc3e3cb08acb2a4c7e2f6684d5ac8e8ea7dda79ee72a4f32acf2be5e360efab18cfc825b7130;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a15e7647c19748160f4d086674f54aebf2bd67908941895eb59fce4e1e2849c5d04e504d2b15ea43ccbc5129f515c53d2a82b117171d33f88b8f6a57441926d66631d4a34127ac8d46377382bed77bd0757dad3130087b59e124832211bd3986ae02a96c1092151ae56f22c37655c68d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10f40d5b2fc1bb3c19180cbb41a231abb7251633d51cfa5f4108eb405abe9186fa751fd77a87fe3d9bad043a14b23509bb8407fad5bf5c0c473384a2a021b0016265f0b7aa3f007ed173a596ad093ffa1e73c9c9dca925c79e4cefab9c459e75a5cedf1eb102109b8c0ecbfd1247b428e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bb1891b199396b8b1f4f9e15bec67531e886863669dfd48416f660670ec104c3d26b23286e67b2f06b8914ad98d0c1f237aa000f061ddeeaf5b72a6368013acfcda2e2c366ef2bbfdcea2cda28904e21ae8b5f6e1037e6ade8036a96cb0af4d5a23bbd4ce2d7ab534ab20ed26165c10e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ba8e6ad3eb8469bcb6320c0d0378405e6378ed9e42d498704df8002cc66599ecf7b98cb98e666c9b2cd5ec87f51d3ebd79ec47e403fbf998d33e5b9c0be99547ee4f4745ba5f86e54e921b3d43b75b4c5ed0b606752f56b2b5c0f3b9144ef9aa32dc5dad6e506232e2c44239f570951;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf10e65fd9a88ad55dff8d707ecf8d979102aad5d75577108e4918a2fb27282fb81d95f4380a44b56e3c14f4b779a9668b6f6f135bae70ed18925a5c91997c8caa182212b2a15c3a45baac0eb56d37c7c5d4c912787ae457487ee282cd59d50d8824d991f211ee2df71290601443493eb4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5354bc2504013d9f16e59a6550c33a05d3dc70c4156d02721b180b0d4b23b4aab822eda7695d812ef9869d6651c59b548a6c371dbfe9f6a188c4efcbd686e0bd429923c913c51b1c2a44e99ca0c8096935c4352daeca938e64e06c4d667e04ee1ecb7308c3ca5ba8cfa9d0ea6e314c45b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77acb08927536b43d5a7cdac9373c050b9b0f7b8725e9c00e1d00ff9cbf69de5176aa62d3fc04e648039eff78365f5367ff9a6d6ca42140f55c4a739b04fec6dff7eebe0db53ad42235f5e71c7042ddb8f7656b37540b76f86d0f67dc21eac132709c9d5e78be73523e1498fd87b9a556;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h762c93769dd158e039fcd389880dc2aae57097d4e6d5a7eafc08ced924e9beacc68fd37251e5d11b97c8f6b26af121c88bebee80cfded2cc206dc0d3b8266ff4da91abc738327e8799f748cf0ff6132e0a4023f55a947d46037990078ddd609211d6f0aa9bd3251fd764ea8fb3212c75d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1698a45a192273ed572305a41e1dd4ff028f9b14c42ef9cb30dd58cbaad55d7642e64f86f7c5c2f7a2935e05025c5414486f78144ae3df710db6dd7e6cafb35759e7f23eed73851f6d9659fa8d4ac7361b2953e6b390db0da86a9daed78fd920c15e33634f354941e21a34aeda7ada034;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3269a45ff3fcf8b8b14d4e7e2a055aa4071e7b48c0f723fefddb10ba91a2b0bbdc55a6f818d543c8ffa069c99e49785d3ff35abc8df34d2c9f1897f978d92a3a6e7e8f72db26aa36f94f1ef803175ff55d7c78e0fe6002688fd4692c0e5fbedeff1a0fe35117e283547301bdc027dd748;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26e7dd9781adb6ce839c7f6ab671b99fc14d4343f2623ac00ff522b3e4e9c4c15b5dee052d291751cfb4a67c3507abf19ff46e3419b7249489a73257fc9396a26a617912fedb06cb7b5e22147e9bffc3b81474f3167379df5a0b74d702e3a43c4c8fa8cb7755687aa1b565bb10a493746;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4706d40e987071a3e4690c3b8c86b4285529303e5c9e4da8bf0aaee1f3ebd5fcc8785c18f51817f6800ad829536cf326cbfd91b7fc6b7cb8789df5780a2412b5331ba9c78b650d4269a9878a6b8fee1dc7f69081b490d7257fd1ddcf5bd161f85e0ce501ba1fc706ddef3749431804852;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c4456919b35b22d42b3572ba56ab4c22d2df21fd5e88c3305cd20569a01264f302a1d173c67c464c2cd7b942c73dce05aa9038605ba41da63ca8c7d21d35d2f670dba7a0a236ad3aabb23fc68535fd88125bc620c55829a3ed6188ca4420b34207b286a53a6e67a2afdc5553fd1447b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4516ef42ab18a59cbf6ab85d930ef88c75c56f5f457483eba4b404bec7d49b51363a9ba2915ee3a8a804ead8297978e4c54eaa2137626305175326b7cc10c9299fad6fa541724aa3d2753f37d6f8ea577c53f51267e786b1ee1b92ced4ab8191f9e1af375fd4013ec61886b1461bd352;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f5c1a3eaf728f0a464759787b0c1e890bcfd87ef8e574a7e9d8752e09b27f9bad23cc91281f11e66d52a325c21d554aaa2a52ead588c74dde6b5c7ed9488cea8fa9d92ccce65d551c7bffb7e5f2e88a8ab602a8d3dca4e98787f96d2175ced1f2489e79ce173856df35c6c916a8edc34;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h384a274e5f5f47a2f4aeeee87ffda733f271205e824f17000080a4a137a2d87fdf7adc519c1ab13767c693d56cee396a2eef55dbd546a7df5ea242bab6156ac9f9ef41dec2dca47603e841fe1cdda4e3154fac98ddbdd8f156c8466052919d1a3f38109ab2b7bff0299bee448d534a7ab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23e25d3bd1e8c2de276de7842166f27ae600933d8e41f86b0c30a796a94862cebb560660c795a9a55c56c9e02357f6eb4ae8e58d57573f4c0eb18446ac89c9a3ae491884ce6876c40bb276c32017e97b3497545e5c73d219398b8db99caaec17abcf90c81185dee9cc4c20172d008fb6e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e34a2f3c350e36507b8390c456bfbbe55b1cfa797ee55223dabe21bd1c8af893f76dc9dccf2534fbadbb8ab5bddbdd8993852f4f3a4e5a353163521f526885bf3912ff27379ba2f53ad85648e4d32818ea2bbed83ba6a3e9c1bdc63493b2c304de4cb5a9d9a3fc0f8ec2755c1161ad8c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd44290b9d4e6c7cce7b7fde038d9c6589e57a43a914e568ede29bd70608235ca9f0a58b191d8c1a6efafcb82325044b3e46d132f34a82ad0a448a163b6ea77ab35c36fb6be4bdf0f71afc3b7e20884244c835837cab5fc9fe23f34a1bddb2f1725bba701c45d97b3592e4d4d6be1c1a62;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he302549af99f796d4af676bcd9773b7d4ea63dd2081ad147ed40d7c2826bf1b44daa7c61121bbf965b782153969a484405f0e7851fb190d95224374468f773bc2fd368de05eb1374ee8ac1e2e5dba5eafefe028475b7a3b6f802da2adcfc522a0290af7f199e63481ad2a6fac1401afe7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb3460cb3655c235a3d04b6edc9dec6a40032e731cd0ba18899b3dc0014f70877832bee0deb3b73a118161594b9c10d56ddd5499072c6e1ff2c26df9f26f07b4dfa2594d759f6e81febbcae34462f22929ff5c00a1aec4df6a6adc0623c1735389aff2bb2db86532258619d7658a276c1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc47d6d21eb898b1c8bcfef381586de1810bf320f27c890f476fc39330f9d441c33958a0332a280c5b74a7d7b226064b1560d4838615b118db2ea4a435fc36714803ab950fb938f32edfadb07670147cc099b80a19569a8af11e8dea264450d7a34f2e9e26f87c51f1b5b38afde2255eea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65bf36a8dc44bee7ca13f6134baca2aa6ab56d432dc0a897d3cd9c11b9d91c56a793778a944ac8d20c0e253b796e06f55f1df90310b413353d560f70bd5641f870769632599568a84c2eb2955b2b21985edf20a48cd14958af37433a5cd5799dc898a78284e311ad268bb09d3d37b486;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b2d3eb30765c1cecc1e1808aa616f2d08b40aaba5db2bfc923b2b086dac86fde5e025f434f17191dc5986e344fb333bd36e77b9b5613839578870d83559c97c4bcc5ec75dd34599f0512244525adfa8b988ae9b216c8862fe1a72ed1fbfca69f778d939ae9c1f0496a6cebcd890a40f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3143f518f020e6ea8c8dc8fd3e0e5c8ccae95a19283e70826dc0d02f982101baabde2c9222cb01abbc3184148c8160d9eeefcf8d33bf9d460d62029503072d06eebabadcc84184f413684082f896ebb532a7ef3066ded893d05fbadfbbcf642eff42df78291ae60f1a4dfec111fb9e3cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h736fadd321c19e9bfb2f43de14c4e931589bd39ae436e31528d383665c3f3b09fa9417b0ee62d8748fd6c1dc02a735e8ca7fcb4de7ce6fec78ac09164e433f8202fff5cf674ac52628fd5f4997dcc36c3a08cd489ca594fe3de3cbbef0b4fd6a5cec5591ae4a9b1cd97df0cf18fa82e40;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb44be8d43eb953dcb398720caec932375b9fa155757f7e832afcf33f20350db93761f4ea49eec1eb279dea21ba928245bddd71920d206497f5997bffeb02fa664d03e77214606cf5a47a29f0c3766c59961fdbacf86bd7a380b780a60d44cb2ba176722a0ed5ca5a8b5a360e0c6d4375b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7bcbe355a82ca113dcd469bf5ee006e2d5bd5880151636075dc87df448533610bd5a3eddd046beb446680a14318ebd0f7fee5c3a8fdcd4601e649cde620e4024279a884a92168df34061b5bfd102cf0a7ed6e099c578c5da771a969da888f0167bb3a866be807986b3107efb4156cab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11e436e2034d887dcde61f39fe9682796439dbfe3437fd4bec099ae27c0bf9bc6fcc3de4b9fbdde701c3bfceb2a56192c7ccb1b126942d13358bedd7901047c19a90eb83762175aee6c82a539c6e4e7b301dca5807d54cf1ce3c2dea2d369a1a07521df8efe9ab7208781c948407d8d46;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5d2f0fb6beea7b8d9e89131f81b373bc7db21541d921236d8616856ea7c992f8f7e19e5cb2b4b603f305ad455891ccfb8ce8c314d9573cca44cc358df976730e3f46994da952e26bd9be64cf3c9ecbded303fe1c4a6d5cc0f78ddc2fa85fb4552885f5589fee27c8ea472575e940193f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f704bba07567696010e4698a2b6333f7097a7f72ae98853c3d03cfb2501ca782770fe3c0bb39384f1c79f387fcb3d3a8096604f698b79ef18457d5e9903ee3c5c2199cf7b117710e3759460cb6025e44084079e141b5530bade8b1d3bc3261113a3612433257fb4ae4b721fe8f854d16;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h584c8ec853976180c9513a912f071fc8a906a7ab6e770714e7f5bbec7dad3c8d8f2a243afcf7f2709e7fc3761775b18e9e0ea045b6006a7c226833e69acc70d2c7b7ce4699b5a1720e0e648ba5b9d162604ce51c70ffba0f511ae90259c5bbae50bb20991f87bd661216ad5499d1b6726;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha730c295ff347f51831e0ad351ee312204ed759ad086caa5a0f9408b6502b0995f81c66920dd8a0f4ef73a82159b2069938b0561d519b76746c672e7bee202d6a9cb161436c98363053f9dac55dc065140ef35393c168bf79712609a5bd2c5f2ecff357ffa26604864be550356edb9c7d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1935b1b3c92f6a1f3a6280796c416d2a0a5fa8c253c4dddcb5cac60da801a9c72b79b66dceeae12b7de60627ef75ae131f8c075d787f8166f2dfeb35726d2ee47805120a22ab2eb8882ce2546ebf3d93e9e003d30d53aa0870d641a4b86d40991713abc2344c375dd806e93e304655dd2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6daede9129e2781dc1d5116c673b0bd2e367f03c1a4c25697c984b39216a354661de0483907170437cfee31605af1aa411e8bde766498f2d4bb66a8ba49fd5186517ec2d69561c2cd5077ff31e62442a0b728bbcdcd61261837a9ba02d5b49a8fa1905008687fd51b3730098b3fac3c32;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4183c909ac5fd33907892e96bf5e37349133df2add3c18d67429cfbae0aadb3bf0d2d3f4be0dbb847185fa17944b2e282e4a801821fb9421e429b6426b450d8657832faad48022283705bb38e493da42be396ed4785912d286a15aa7ef761081bca726e381c31dc501bbdaf80346cd386;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1f8f403c5e8efcbfc37efe4bfac880d524bf2084ce3e921a7d2169738fb674dbd4e8c0577ab2cf5303a6fcb291a78943b5ac5f1e9e1900b0292e3e6107fe0ef5f25828d7b1da3661828061fdca1cf72fe5e2a0f1b40814cbfa2b81e28ff244ad7c3208632039eff20079858be7d3d145;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9110f016d3de1e1cef738f67a5ae238b47455f1ce425de93a73affa8714ced0291e99f23a8dfe2ac89923a7c3a52952786675a58d2e22e5a887ce885da05af3741dbb0e0603b977da1811724e47b0550c128cb2e0da790c22b95701584c93b91bcec11f821bcba4b6eb04b30274ae2ee8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9264ae49ebdc7f9178068cc31ce6a49229e50f972a3a9fa080bf58ee80b9ca9bb1b6cc84f8731bf7faa490652d505c7e1f1d8ce78c575cf40f135a2b5f3f8636d185d7fe91e608f5895261f05d4b9c62b03ee5d60a3b20093d8dcc43adcd1cad85d199de9ea879c0ab07279b742ca0cad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ef3d0eb585792811ea2d82f9ca9f658e10840e3ba177abf9b5954b18529b478380e557f850024c5179bdf39c9a707b3a8063d69ab4235a146b650a7382268d5cc4c4a9bb2cec758304a4f01e4c6d2d99b452ce23fa7c1556584922dac917b9a577626dca116a1265eb1b1e8f19d94043;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dcdbebfdacc77a83db1736c24e839e6aa57ca34dfd41327e58b63336561ff4bf6ace3e71d058b8fc3fd80d4461552293262678360934b463059f067955913f869205461166f678096b75f9dbf1cfe589ecec787ce7340eb3e7c5b09172e56acb4aa2c5fc4e8f40071c3a8834eda3c1cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7e81e95797b145543bc9d96512eda024ff979c74b4b5530358c564d0a226f08768f83fc684a9edc51d7d9b6211805c1e02b64c37422d00cc39a31f9f729dcbe7d488a760ca554602706cfee6492ff57e1dbfdde5f5499ddbdc00cb21c4122e1aa25e52d4a9fc4470f870e88a23534485;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a8e7c2a83a1c0d6df0e3d300fabe677174ecff6cbb0fa0215c869e0b1f0f63e2421ebee5606eabc998b8912fb9a4334107ba2b6e3c55ba956a267f64a80506f6d1c410baf74ee0c19ec28a8ee1139cff8542dca31c457b5b7d72fc6fe03d2a4f38602f9f277e566a734eb9da6eb9d30b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2be99098358f250464161b0c87e2690c8b4fa07a21f0b72abb5cfb7f6210b34394a14133fe9736385d1bbaa868c2a8696b2e219ac31cb366c8662b41252fbf91a2eb354ebcdc8ccf7322e55592586050e67a6c737bc184b235344231f38af447df11c53796eef0ecdfa8592f103bd51d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf124090355f87d898af18e3addba63be9d88fcdefb642020c253b63e2b4348b8edc57206423385f6734cc3e6100e4cff3ab242e327e747357dec1b31eef2d2ad4e64d66f4985bc484ff6ae824a45e4f4e99e20241e5590fd07f084fa40162e020c3e5c0b12be386be94853fc1ec2230c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6189db13ded6132adf1885c31a70bfbe4783e646d8340f42fc9607e71436c37fbd8d3e35592a93f41ed48a9838a92c0271216d38464852de7fbf0a028df0aab004fdbab52f6449d5aca497bd1ddde216abd4b70bf730a30d39eb15b7cca61b35abb1199febd81be4b00e4cfd6478fb246;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f87fbf000bf3c0ac736b42552e46401e56d6d6db303f00a6ab5cdd81da073b97f6d6905b434cb53ccce32872b3cbc839ecc68b7945ed5911ed58bcc39f0a33e0ad266c2762215c1d521d4c4d9090c2c3f4cf61b4630a37029b89738f5520e2b06a5da5e914cf9f75cb0081f868ec4535;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31a61f9c7fc24a5cc2db48329210b25038e3b189d63410843b5773ec46f7092c53484633aa3da52ac9cc5227fa3502bcd9ced2b9d7aa9ba0c9310b93cf38ba737182791a05685e158e099b316448fe6b781ef77c8965ec392322b3d25fb94d02f3435d57817fb32a33ee1f059b7daf2bb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75045386dce454eeff985a8b53fe573374ea6aa27b7fa3b435c314a18ed1e2219049962e27225fe940b62cc14c0c0091addd3edf2f601ca47073122ec7215a567c64a2811e8648e37c4ac5eedfe666cdce33c3595db4d93f8b4e9e839c324f81c68bc58cdb5b1b913f888aa4f01d0780;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd9255448fdff15f466c88ffc4147d936ec3c2ffd377f416b16febc8cfb04e91bba0c28736096855de5ca35a4806ed1dbd16f7979d27b04b49b4035c1b3b2cdafb0b4da2f6a24df02e9dd780fcf5cc4a40fa5b42d93cb8d11656a280708e1305a633cc1668f00ccbf313423b7b7734ab6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88342eac08ce90bd782a8f30df2f2f533c1118068467f307cb70d4f69f0e5e7f2a096ac017c229c6135547bb04c88fe46ded48ebb3fbf9f3a5496030a5455617fb6f986280330ac8f1f2131c8bbbf25b3669ce6bb8c1eefda8e3b3b8b1d0120ff2d4e37b01c5d6eed5f02df271804781c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda980aab9a92727b0bcb4f67fcba0c059d9cd03a7cccce35e29195a5b276c86f621d973daba3eaf852ef63bb3272c960e97077de6306ca1a107f7bad66e0bcdb43d1c2721008882413de7bdaf891de80ac74a8e32be7d3b7d53863f835796a9def27e8342494833badb7f74e908feab3c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64aee426fa63750802bd0a53ebd3fbf62e2990c5469f53e305a7a852263249f104e50c031297a69263bf74773fe762afb9d2c171364073cb818ccdc94525bc469fd4c91b9d0e1cc935e607f0d6ca09a8dd614a47b3389999fa8510f87cf12fb7076f4feee5bb9ee2a778b968b6522410f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9162e4a7c1c3dc76bed741f9cd8f9d01dba92988e109db3a6f8af3cc2fc17f3ad0d32aa9599364330c0eb50b75aec0b09b9c9bd3f28f62cec9bfbe6aab538b706ec7bb583df447f29430607ba9b73484c6bc008bc8319f7421bfde9c5fadceb344c7b419548669e92595152c175a4a366;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c869fafde8a0f3f2b851ee265bc46a38cea86fa46915f14f414b361c4ae4d8879dfdd4835a322566722dad074fbb6feeacf356a7a0171feca9c0628fa435fd481ea20e08c8c55be9a039d9f0fcde383526959726534a06d313f205cd2c2c98b44fb2d3d21e75b39562f92cd5e9f90a38;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12dd4360c767106a06d575e9d7fd4051188f7db407254a64077132fb78d3fed1354d082b6796618f242fa32742f5eddc52fd8f14c88c61ad2f9073f95cabf3371025030e7d58799dddf744079d4aee188db7fa9cfdbdaf6abc218582b81b0b94e3336f36b11082632262729ba41175691;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c21d550b8e93f6db472c9fa6bce4875445e9dc76199b68dfbe34fc89c94caa51a017865e35db68cb75a8ac50abe0b984e85a094682adff461654f9d564e0111683d4189a108ec6de0961f2f341825c2ca892e699f7801a0324408f57503c8e331bfba051f31e015bcc34d3841bda12bf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4684a086b68f7c7c2b36023499280d8a73c98179e0f421e0e3aa7a464bbadc48ff36934ae92bc793167550eec7142a8ebfd8ffc237e76594a7bcf554278af3b1cd560e673f91a8ad46302098e40e58cddcd276e2ffa34d32815c3be20071cee2589cf6b53ba81aba1e9c108082833efb2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2362d6756cae9e794710efa3db3be87b4fcab555a31a63d67e55d2e9b29e7df2662390651af9cccd8b38582c66ec89aa0db1788e4edfa2183b903426a76e1a53cbbedeb48d21217fadc8becb105fd63193fa598a841568f3b5a5a552b695afa255dba38ef8e0d306d45f7d9460e1f87bb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb05b773e749248ee8daf39e643e9ba9408a091b83c3cde34ea9af779545cedfd34a39959ee043f7619efa7e334a5a2e55d005a086fff04219ad245676181fb0f16f5f012871f1c93a787161c497c71c9a05f60eaf417b82af3bfe0b3585ef27637f75f9030fd47794d01619fee13ae65f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h362755ef93b43b357b9874e788374527438bf39b4701bfaaf08b63d41084af06815b2f3cd03c8ec9d5ff96be9c064634b31cdf87a47bb7a80e7e2c8d90d91d8bb91abdf91f539ac5edfb7d51d6bf90bd77c18bcfc64d6cd7b69ec2a1714982f9db92168ec5e687f6a2090628153b2ad1d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92c659f4a8bc3528ff4a75e343684ffd4a7fb1bd15e81615af9ed171729d91dfcd928fdb9b07f9287f26157370b7bde43a35d413bd9096a6f38b1d587d2e8437e1c8847887f8eed1fbd47c95fcd790f2babf70c386fc5971cc09b183c542ae13ace51dd23cd5e67910e57c02cefd09266;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a430ebb5f7766893807afde3253d4e99e74c1041b4ecf86469172210491f3aca6bedf8beb9d40336212f95651adde7997ce9941b9ee580a80b27cfee2660e784f56e274ccc3c8034f5ba04637a971bac2fbb5a00c75c117d2b973d9d8c65c07f16b9604f6026d2da153c476094dad9eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h935044b4c9bd0c9b4fa4bca06fb54bf96226423e26dac7b8801fa3d61bfeb657eb5f84ea47e208aab69012157cfc165bceb999f9bcfefae976934e33eb33ce1f52da116f8dd57e8aed282d7b3e1e1bfa0c7d55146627120a76f8d9ef0c94133c3d6b45a73ccf752351d141d1a51d70c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34ec79d1aaeae99f62e0d10c05d731276b4abe17fc34f75c0a3b4a9253a9cc273a7592cce37587547c5ceac8e4f6cc9fe24d437bc6c620b7f380f3ca0955b22e66028e3d4b977ddefa0da90928417312b66351698f4b306b9d1f61ff79ca4824f716406263a0ccf9c1d9a1f99c97220df;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5cc4572f1ca1f3dfa76e50c657e65750848b0f9226460ef30322a28b672999aaf52d8287a847d7fb7d4f696ac6b9a967a79d20c29b575cf8a8d4d0d6c69ef8ab8afd3dba2c3b44dd31cea093de23a388c1a7569cef625a164f054afbea7a8ea3e789f90ed8926100dd5b889fd9725597e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hefddfea9ff1c7fc6835174b168315268c839d62e498398a9e8e71b3bb439be17ea63ca50d936fe7ff233aa14d2053fe55e3efa45ae01a7708a7eb8e79f476a66f8d5fbb448e7963615fb4bfb57cc08a156db77288480bc15e8db39c5ff32f6782dbd80c0f7585066964f9e35cadc89819;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8fe5f5d9b3c84519af04f641abc95d99f1ce7dc9b5bc51e7a434ad818d1fcde3c4ff80a0cde0fa2d47d40efde7eb8c8da34334ee37fd33d408fe82876b2e5c241a9e51960438e8f8225181477c70a6f5286c9bbeae96e9a288949fd2107eb410995b59587f11deaae864a160a6e3917b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd554ac8c7ea6b3b6c6ff037d03f331d11935df80a82127b26427444c0b1cdbba95e01f1548812be60654f5b0461ea822b3c121206608eafa0bad4b5321908dab6347c0591276f3daa666da47436a19ab2ede7e23aacdaed384bdaf4942db0d784c7b4446cd13287e54451fe9d669b4a61;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h825f9aa63bc3f27651099e1d999a3fe2eb85649524aa1b39c39d0f93d30e8b3086605a76fe2051f5bc44e982074a7e424137d6b8db218c5bb59a9e7b3a65ac68b659d06a2ecaa1c520076dd70255bdba9828bc1b616e326910f4ee4f459d29ffb05224ffbe5bb3bbb12e296f4cb176aed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2ad8beb0dd0b16937921c61fe1f37077b0e21c38d8b1e235f8c32a1fb38531f6adc81fc5e71f2ae19236d03c4821b26a0b07e11bac258886317a154f847597a58dbc683de8855f6b949533986383454aa9c63d7f3d64c337b9c8905871cc6cca68981063244993f2ac2db48827a7812d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57b24bedd2b82ac4bb0c41aaa86082c3598333d0efae19612da8f2b159531dcd3bd7bbfcb8c856990f156658612343e87b0c98aa92e7272d78a8d0074babe627dda6985d117a9e4914a454a9c7e9b256d9b3b687ec9d3a7bdf20e87e7719c7edde995119719bfcabf9ae44879032023ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf624d72b4fa747e67691b33b43ff2bf6c831c3044d2d98a142b195b7af7a9edda67474eff2d96c39c0a4f1e43f1eae4cf3083faaef2cf854535ad609829226a62a030e7c5caa95e5fc7863b990707ee7816ae99fa475b553fee3e5455ac25759ff2b1039f962a8a89255ef318daa8d2f1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf7b350373c52ef2a4d50b8d2a8e59478b12ea39432b9507f3262743bc6bbf48630dee9b42386a7ba498db24dd02865ad2b1c4eac4d2c0507f7fde53672fbfecf930233cde1a303b21132976d018d75097eb83fc6e315fa5c075f9875b4d683f16647f851b6953ad128e3958daabf77b3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b56cfc1c8915115743ef283b0f755f653cd6a56d1a8f167ee960d9e579a7cb894ba33f35089fb353f23cc31607cedcc41e918ed2915d6f6a03cbaf70c44d86438be347691321c0e7c4abfac8f41345a87976c4f99a8915d4ea68a7e858aa89a055dc9f968b5dbb00bfe73309bd22c664;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h573c96cb7b778aeb1565ba9f767fb750996501c182b5e24c2433afe0b3d32a84fb384943d2ae6ac97fcfe952cdd0a36a7b288810e08e26ea8d32c882bbf989f2aa9452cf9a625074904e80db49adf242c2c0fd76e55c6eef82977f258d58698c1c82d5f013a7333f19764b839ead2da3d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa105ea338f8a48b895db0747e19ae3a5ebdbf80c0133392a968fe265b94113ae63752fdc56ee36ac1ce4534eb8eca51e55f958534725bae47989064b54876dff9eb88cf7785ba793a8208d4cd1410dd7376c49f7859a29752140058706f268b26a063df641d8f0dfc2479146662bbc46;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf98b0e05ff0dc15d7d1fcd08132b2996295337a3b50aea33450e9d79f0b52258a2b88c4954a49f05aa1457a0401ab8ee40bf400bdeaab18a694b45617b97c2954908b6975c4f92b269c6a49157a00dd095b7c98da1887434892c1d05bc89ae6232326fc7e96a995d93ed6ea61de295e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c437a0f45d138992b69fc5d595a83d42d0aece2b7f0792b150cc6c13e8b574a350f8d665cc8cfdd5902404b619d05ad838a3d0c19802aace5f38b5babfe06d0ba1ee238ff4704415f4c19e3a9f838abff45dac332cf00e94811fcf0445bd1cdc163ccd7adb148878d91ec96b9a35fef4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e1076ac7ff8c028cb805731a5f5f5e090e682ed89b8583e03aae3444b141b2da7b3abc8ed1fafe472d16b505c2bda3f2417f0d4794d925765e748e6f97e4dedeaf463eadae5c8e4d3921b9efbf6e77387fec3ef689dea2367f095da8546dd570e4cefa7179897949e5ecd87fe895c3aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h425ce82a884cd061d3235a6b173faf68ed4a168b134cea29348c5bd27318152e3e4ebd8239adf7f5e8cc24e6435c7a0bce6f3ae30f705d33ce2d4118eaa75c12dab63945d2e87cd6c0d0ba99f4da8fb37d4e57409fd694d6519812812460c05f89e08ef8e028febc22cc89b6c515ba9f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6619fe6638dbbfd84ba9f1d21fcdcc5c78f804bbe0b5a0e03b05767513e7ae2f353c6d77081729bcfa4a37903ae630d9501e25f3837d3d68ca950b0b76f84a2f0c39229f394cd93ff4dc1b426d2ff504031025bae6ae91fe3865e9ca271928be91c0d1dd1e92796c609a327ff8b40d4b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d513d2f8e14738f575fcf9ac86d3bf3d92d8a153300d9c7b291c73df7fa61367d0f1004c0ecd412e74e5220f0d882a5fd00530c71f05cecfd6220d7e85bfe6cc8addde51668f69f3f246b1697457970ee48bfbf109e34057eac00ef3a893e8a7314a2e49af04929c1a3333d8de71f7e8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacea899ae291abbc6691aa9d97535be761f7df66f3d914b5f29cb894e5fd2cc190a522a82747a66dedd309b408373cf0f13d91836112b1d482faf652e4c6e6497d3d0cbc46415474fc146f6afb384800ee21381909ee83a110e1845671c7597c23da58964ed5b094e026c247716de013f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81511980b869117de24e16c840df69560fbe68637104e45d22b1050f11b4dbc8ba07feca8072cd3cc8ddbda5cbbc4b430a9f501362c8c68fd44dcbdb029ee94cb93082b14fbd8483d0fbf19e43b647038f72790aeb04b9056f769bbdf6dc0cc56fe0c89e98be3e1d3fd14275a9bc7a9e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha037b228782ff9b48e9063f41037899d4b57b387cdf1a004d6da8694b79b2fe66aa176e42888c8134b9d025f582b3b8aa77e2f58d3ea641c0d1a879592e4a2991654c5d48107a3e65a9dece9cf1b1ba594d47f858005fc513ff7acb70d1051e66119c60cd633341591392c840b1cc3e49;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h262347020964efcd21183c50cf964ab5ca2e26d48aa0d22915f2216207fe7e512984c3140d966ed12e9d9a42c6f437fa70766a93b5767728c28eeb8e290c675840ef7580ac3a0917032abfdc0418ea35b93a3431e49c9aa68a4554169cbe40fc7612ec0efa3248626883ac63eba7872e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19a9ae522580670b443ddaed28d2ee9d865d72dfe446da99ded39e02de3f4e89e94caf7c2af2d393540945f164325d0d25922c4d7a6d7530a423b7202a460b8ed3f7547cb7841e83eab4ee6a6b86f9031008a38e842774314cd4fac11b6ea0ac9314971b06b57a16f12e6987e826ef225;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c76842562eb5661281a3791d6932196f7073172c6cc8aa4778f5b942d69baf7c599a78f26396f917165a80f3c536d3471d093c575471730f0f9825f99c35cba352fce06fb408cf4a870828c03b145b63b16fec5b50c530ae360137e38373c88a9d227c0a4e9fea9659aa86e667ed6ee6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb62a810d370a64eda4c718200b1e3d0c65bd92adcad94b499d4247815ec2cb65c7950a259faa412db62bfb77cf50583b72999208f8a0c2cbb8c400c6f06f91b12460386d89d40c27204ed266ae5594ba0a228e0107b41c8c0755f5de432077ca6c36c425aecb1b38fbf3f6d6def92658c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2297882ebdc8836592cd6437a0e6e36da790a3ef783408e9a76838bdea663899ee89ddd42126a8dd6656bf797d2c13a3c8b3cf94805575635bca9375975de9285db6d9b493e791e43ca619795543b7d08b79b82c93ed1ab094442ffcb57d1627c67a8f2c53e962fd1918fb246a6eacad4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b130299ecbd8679c360d5e46402d7b49799cdb36d2866faa8984c54681a583ebab1924a00b3c08d42b437c5acf6d1a6aa89f83981159e0039ad7522fd0110b86202e286dbdca74fc8cabdc11bb9a0fd636ecd4f82c01a7506162d71ad3dbeda93d3935406b15d6f720828ea6b233e59;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea761901f5609c7724dbc6195855f0ca8963403afc91b45af8af138b6e5acd12f3d6d14ba410ab2a0ee3add496bcdb246c6a59f7e501266a019cceeed4ad5fc8b6319e5bd6d28f639441a72fbca6467dc0566b8f3733a242834f33c40de2ed679a3625d514061134259a75471050d97e5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcee6995bed333cf0bb46fe1b3f0d6f4dcffb4ce87e9306226dd88df855d99876a4c24e93ad5e1f44620aa981c4df70f83467254c569b3bc4423f31e1eb3cc344033e9dc452dc73e98cba37d9f021e2e1e73e4db53b9148078acfee9c1cb3bd862a2211b9ad3bd030370bfccab907da3f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb595ffe917cca093b99c650431feb07d939c3d27f98dd8f7ee263885762227006e1a4d18d5c02ae181f35df5458f104ec87069eea28ac6cdcd0ef2882bcbff8d56844f8be240135c4a116044e281c0304a1f1b610e34f5e998523bf0dea31c6fa1f5907ad8a7b9ca7d686aa77dc70652f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6025b9dd517c25a6d526a5b1bbba6d771cf554de8b33eeb0652e74062993ae27ecbf5a0e7bb67333ea544e49ccf1da514f36259fd73d36c5425741a367baf4c04c6435914bc39a7ac624627eb489d0f07511a57779dda8b7edaa9c601589406ddfd03aef3568a5558b64ca4dd06ef06;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6eac521774723f64bcabd6ddfe93f74439d3c2f3438c308bdc745c3e384adde022bfafcccbbdf4102281be57f26d12f0484d0218aed66c75fbf5e29ad7ad3a8d0210a7030feda8c84cba7d0cf32ea85cf1ebdc863266f6338bc97c4a81f779098aed6a29c563a6efd6afe98f1d6c2fe9c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92f5fe82acf225226ecf4ea83d54c0644b0f642c1815f0a585da25796d5e0f769f1608981acc85fb9efd195aa9450ed3641e988554b9118162d6439f802fe16de74eb5f453b8b9061b695bb3542af3dc373a978d3ffec0c033c29a8e8be708043f0193675b9b96ba2a39f85a665bf3f3b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b094373954cc03069e384e88b422162ca1f3936c3057a330fa098d3a18b9006c96bbb530290c9ff57d6a1a91487f98cc6ef0a84026b12e2c17c86d7705a88135184b3a94b85040c50472dbf35d50c2757ee6edb9244b45c2559ad04f04743f5cc28ce090966d8005592c018460b87ea1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fc9843edfb008f3f7f2449c6d50619383c1e16608a4097031e16d8d7d70579682ec7ab4e840928480dc31641101e4c76c7e235a08a58833c3d96bb8ce916381267408a72b1c48bba0bdc8427360d718a23b9ed99706288cf21f3303e139236601cd6b54ee377c5786059ac75a580665a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdf2fb93e55a4aa3aa27507a1a445053c32f11f1f64f6591952d5122a24db73b57e54416e2f78da956855b35562a6eaff7aea449fc4b2f0843a1a43eea7721c15ed50c85023af7b2c4b13feeab14a85db5ab4a7eae848b1d9c9eab67c6ece07234491d0518f734f585c1f2d407a8899f0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19d34ebae059e3e4d5348086332bbe2fb0cb47ba0094320e680abf01fc851a3b40622aad7fe689b562d4411fed603c96f1248a794378a9763222c3aaa9f2a04b78dc7eb62d9c47eeaaad9eb7b6d3e327f01cbf5a7e3d1f70e25f12794860162a00c6d92cb02650603800dcae177abadea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed146d5c7e86e7f6a1ad2e01f046bbc710979827f98810b4b89bebec59dbead194ab891fcc9ea3880e94e43c80236b32a9a41e9767256142be821baa3cee05b8445cfbd5f0df9163ce5738987b9cea5d47ae9b6dcd8004738de9f5b8f3ba7eccfff7fcbdcf6d8900bdd14c0889ede0601;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h910a5441d321098b1a09534bdfb9e88ebd75f3daba763ddc26b14b190ab4f2ee508f002965f2827482e86e1d3fe289c0c68a061d388dc2713e1f839cba7994316392ac9d25b2398b9f80e5d272a2e2fc140931eef1fc9ef94881f774fa07fe5a6e522d1030ee0b2abb5be2cba23b365a8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17a87759da8bbb47135fc118e294ed036f45d08f01485101d4efce652c64368dbd50f26ed19fd3389ee8fe58d0188c6dad2000a0a13cc4120204dec3bad8d26100307e3acd7c1cd83deb10240a9fc754282ff9b783588ab81929431926ccdc76ceacac83dc068cc74927eb7915fbdb48a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72d48483b037f2e6f08f395a57fbb37deab7cac22e34dc600f9fff53f7d03727aaa200d37f1f66ec62a709176b3e49c1a426761c9c90e5b9d2300c21ec0194345d4e63778dce3a85e8c849fc0ad21b99ef91c6639afabffafa7f1e4e1cf223f7f5107b8c7c5d99f5bd1f83e1a83a9762b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf16018a5690d38e709d79fb8c373827e8bb6ff083443dd7ccd99123f47d7f6b50cb7de44062087b7482e96770868d150c1f16e4e1ee37ea3b23d6ffe5e8a683c34d53ca46c34a88279b9f4f9e1a8f514526b14dc8e13fd7a5de5d51979dcac6aecd7a57126aaf96a98c0415a26793aab7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9bdffbc7dd1b9bf38449388e464f7591e3083089dff700dad0cac8b5bdd2d6b5615352a572d6600198fcc55f93b8de909ccc0410b7ed8c10733b7394104c10e2e607eb247828ca7652490fd718ff49e58dce6dd3cdef3a93f0fb5085ebed34462b6445c1261faee08f324e57913890476;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b40a45dd5b368b90a448bf89f5317145bcd28f1440cd60f274fcc875aa3e5382799dba3a092a358267d7b530c796c2a7713ee3e422559d1114c13f414f09e4c68ec9560b71d7040e0a5734092185d4b48eda798a5546d6ec6abd7508bd2fb87786a4942ee454092e6adc030c15893d8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1dda566275b913a40b34570f8ac8dbb5867075f5da3c8694bc923b0b1bde7ffc1da49c13f85cb5da6e9f8553d5a946aaa6dfc2c62d50d207be9af90cf31ddee6acd0b1f9fc258449958f503a8504301f921f21ab14945d8a6f03fe621afa74ced9caa5a305c9b8df7e2f18068efe1c67b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h983dc86bdc0326f3070ade3071bbf9829b031ee7944d09e0f956a844e268a44f525215a342a31e5790b549ccdd4eaf8ba11c25ad87ec4a6d1ee275f0c13bea43b9fe3c8ad5c6761f633248a1ce895d3ab4a9ff5b77d4a47205562a01bd807e9fc5cb9486897be15609ce3c30ce387170;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3bc33b60f0e0c20e5d8639b4c947df811a776f87cd28cd1ad57d9f2485379cc719f6411ed09c24bc029e7c65073b26e6bae729f600ee87fe7953143afe85099a24d3acb65d903137595f3dae7174e2bfac07c3b40db5110abfa409b6a6a0b1fa3df59f3668adafc2ab5e8826c2ad4b409;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h730eb3fe53cf7615389ccb456ca324829e4e39f2091130ac1acbef1592a7604aa8beb8eccde2e98c7fabe5bdd2201a40e7d31a14e1c5480d1fc107c6e83db585cc6fdf79fcd3a90780db41bc74e6e89836f292fb2eaf34e9c6b69d446ea027fc4de15b5a97bf0b480cf0e9a5709a26206;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1b9e1419008968c47bdb3c0f4250f29bce972c2978d7f956eb574d3bbd342bf8e51a8f6b9218d309cd6041ac72424eb9c3f0a3ce090fd2e056de2060c891715a923ff86f10d0c4945ee9070dcb04dc1342b2d781763f9a6ca6dcd2fd4116c511aeaacdb4d6468444d42ab98bd5ac28d5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d9109154f5be93f76bf1ab08efedc39f828bc57059d1827279b1d0259876d647f06a9432e00876c3caad5baaaa12e5f28b66a6743829d3fb8fab19153aea92b475e3f1e5eee4094a93da7f4174fe826410f1fa449c8cb8ceb9fb9496ada84722bd5a9c58c8cbb0d12a3f927c76d8fcf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6043867441a9b42c63283ae310af15cebe5255168801df9cb456bf2ea2b8351e672253ec121cc64fbbf87dd6eb4c0fdacac2cc1658df361da4aab31c94beca291ff05a4d0588351ef356aec0f658dc2907bb0503e756a807ad2bd01d2c3125d66330464818fe1672d6c73411f5f12d17;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb48c65947ce5e27ebadbb5ff5f0d70c2312c595bdb2fb9183f3b4c635671e03dbfad28198099df50581e596c37e017fa9f32dbd66e9e8454ea9a4e526ac2108bf1852bdb18e8910f5a32f84a03343c0784fe117edba43dd659699b6d5c19fda037892adf2682e87c4bfc9e9cba77cd4bf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ed5b6a7444e21f5f2cf7f5d9dbafe662eaaf146be550cead234e8795ccd3f97fee17656d226ccdc7f8c08776e0264c45f326fcf9efd6b1f19c189c3fa52b8b3b3710289de9feb8a280ca83a59e45cd2255f8e185476fc8367f2cffbd3b54d609c419e33f11e96f9434f743b2c681f127;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c5419a5cf471176eec2e4bdd8ef1ff204a2977007c571d6ff8ceac73aec53873affb0cef1b5de4799fd852ddde6b857cbc0e04d5edd2adef785d92c827227182c9e3ff93805e7119ad06973edfd91ba1a2ead0e326eb721d318aa62fbdb337146ca2294732174c65d38f272c2758e22a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf085605f38f83fc020a208edc1357a32a4874f5a9ad1e1ae72076eccb5e9764e7bef22a89a97bede2a956b863d747fb3d49bb31310de143bbc8672ce8c60168483ef57d36d2374612de056a1a964e8fc2c665627b4ffe6c7bca1843f3b8c44fff906a443cfca988524993374f99ba6a25;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5f49e905bb9097861a5bbb5eacce9fc069cdc1af18cec55e53b1c1c09ad23558ab1a345d0363239a16174b7d4c1e72a80bb23e2fe60502094ff14f6aff7d50665d5f623e4cbcab807ea85c3788959d8b06575eaa4dee95b3c79fc7a3a6c3ecea4ec2465b0698909b05ae78381ecf209;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9b50641677bbcb09d6dca82345495ecc773528fb8f2e191b1f152f81cb36bf6ecf910fd5c8fa05f131065087f12c8b8ea9adffdca29fe9186d4ee26ef7693a5843d0e62271749852fb48f3b717a91916e3398f3aea51211b352ab8e09162c000456daed8378543af9bbbe6f34174b496;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7f1b2d1febb9ee862c993ae2bf513649eaaf0d809b2ad8b5cabc5eb9d6040c633bbcc4abf646560220a9299f227ef577d117e1809de3c3cec06df781e1e2d27516720907149a98f492d02cb54db35152195c390882291b6d9ca888f29bcf6dfe61f0111c4cc3b70f556927c3878fd900;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c91528f65d0ed27487e0c880cfb1735c7ca7fcc2a07ec36aa41565dfaf1131b7cc34079f6ff18d4fd68efc26228aa37a7ae3f4dfd9ab4be0c4126494493770d037969299ef1a2837b85d2ea44b71b6d17ada7bc484ca746fa9fa76fb5cc30b3a816b2a50405a3a1c271c3d54c9d94d9d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5673a3638205ae3edebb38d22f6930d9b4170426b6407e0f5e2dab52d3beb77137b95df61f4b977a6fd6357d48dc24958cd1cd5dbe3791107e142192993672295032c40828eff6aebde27d8793508d411c17174a6bd3a9ee1f43c8826224c9b0235585ecd4560dfda5bc1591b7c83254;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d4d2d28c4b50515f884df658061bbe56ba2c382901efde9e71b6b1d937c2fb40670c1601aed6ebedc41f7afe27747dc415f1a71a6ccb26f53e92ed94b86d5c4d31ec72cc0b3ed1e6f9d61bb748f2d4068665583077e9b69e959cb3dc5f3bfac80109d12d1b4ce97d41ceb0f4f4581998;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80fe845900160c9411a5021f6fffe47d924dfb5dd2b4db0e998801a441d370515b700f967fa6d793e05df4ce880925a65cc26daedd1df714a2411cd50bc7daaf79be3cf5eb3e4fccc057818634817cd35a8c39d2b54e408975610d99e5db0ccf2a44c31bb3a5e6c3b14e2cde16b03cbe6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1499dfe9b31f71144b429e7c5dee53d630537cbfbdff2f9cbf90d9a280b7e587184a171d11b3fdb88fd63ec56a8a33248f6f78d51321ebca5f8ee46f7464160b0b56901c91b1ef8fed5f71358856167bffc06780cf77bd3416ccc5b159312fea2a48a8b47276d6d13dde9dce6d41f972;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc0aab2d262c0070c2b0c1a537e63c17dee2254ca9a017b286ae5ef83df1fed42e9a998df8a8a88435760aec46bf02a79a80f5ba3e411fd68af34712ba0714827781141bc0bdff575a0f013a8a91f1098a43498360dd6783999d3c881a8282527e6186e262bdbf7225fbe0ae52dcaff117;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ca22a96d2efeec08edd2f57c9aa4a44eb4511b3ee5cc9565cdabb005386fa43c27a77ebf2f12b03b395b81e78fa5dde1ba5d80f6d48c9179ef9eea7fee050c6d2a91e794fc8650a646260fc2792ec4c5efd51b845c1db94aaf7712c92a9c7c40ef276a275112328d9a5b3007e98fc75f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35d5a02e31c2670dffbd124ff42ed0ca70a13d7e455e2094cbb82aa6f8df92d67705d06dd863092f62c7f2fb34625ced9c59cd47da26c182f91989463d32fb49ed6f8d8412bde05c8e6061645d2bf51f06d0ab36c19d7adb65ed58eef8973f66a1e3b8fe1653b393b2b2ed084c46a37ca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcca3a313dc5aaf2ff43a7075dfa231bd72729c56ef60dc15c8d760d2b7924af210be11cc5f5cf94a42f772504c33317847849b02a6ce4045acbb879cc117206c1e141346ca2bfba65ab0347148e8ed427f37749ce2d0f00b123fe0309ff5c80f77cfbb4b945a4ec82443f6cff2c6d89ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9252a5c47df7f969f125a7b5722d21c1021ed20f7f49549679cfb12f992b0027dfcb346d8fe9f0eb7ef516eaa6fbca380e7e107a2c9eae4192a51a08084c0863faab0eec6ac7a4e4f3db236417151ef8363e1709c925151956b608b675c8159e9d9b82e3ad7f86e7c4e6407b7aef843b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h861c16f1428a0ca0a2c2b01268e01a0824fa83588bc947880287680d4c36c05d121d526c5b2ae136ca5d884751d8045e9f22af0b71b95728765fc92ce1cd845e9c1ac2623db3a9397a5d9e57c9696ff79f6c410f518b287aa0491b7279ba2a5b24637e1360d238573a8a9d36b0e4e5fb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfe84ffb670aba903ae9f09a412ba8ecab17ecfce39bd917817c840d062129a3ebf7cc48f80d00b5d36cb605dd2982481736529f5fc96577bf32d7a267d0e051dbc1f2b0f1b5f246470678b437f3f4dac4a57e685691d6f91dd8941c518a75adfb086e5464ee77823f221ab21d7bf73b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heee7f21140a71509b370203add07cbde01ac674d3bb84fe7a219fccca0b3970cfee66f3109c2014090290e29bb8b8ff6b3d790d2acced82507a28f4f0b1edb42748fb9b0e28cd799512730f27756fa665eea1e3a042c01ace5cdf0c22bcc2e004168ffb81a1d08f6fb0e299648d3ed802;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e3919be54cd60dce2a28ac5bc2141809b1aca1069a4460b05e9efd5d735ea17b422ce947b91b1bd4befd5d84a4b85e45b646307458d17368e6d4d1c306a6276e63705a996f2cb65112dee4735673fb2f8879d6b910c4dca211785672836ac7079bad8563ecbf5a80f9cf694539f4a425;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc46895cb52e60b084f946429cbe1a1114ebce96685b1e502865945cbb7c158f339cb4b69da8efa9b18d5d37798e17ae819d9a02dac1122247ccb07a3692754a0e5c61dbb04a4113d3456c83f6d0b63ae6abe2d08dae373fec3637fb385eb1b5386ee2f202cb671969444213c93f34e5c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81c614386b9f11a1aa8d07006b7822755bfbf6450380048782ee9817e5321ab0750d46694f2ba78318ca5ca189ed2ccafaad471a1c819a1e3a192e7c6c0149a63a7b57a5c92520cf5f1124c3af630bb3967bb6d234117accd36835c21ea4b14228e0259c39f68f848663b8a7cbbccf7b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd0949ffb16e3e6f7cc2b879ff7be99f94298bbd7ad502e6fd9d26083fb9439609e55af509bc1e5a5d367c500801ad9ccf1a3dda3b261ec4e0b15b4a24e0190201eab3f99b089e9bd21b8de3b655c8349f43409c1a46a1022be9dc348e841e707f3e2bb051923ee95f6d11abd82ab497c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf95b19f1d874a6b9220bd20fe5116143f1e49d3987d8ad26d25d2dc683aae48ff9866d8f6741d8f25c588c3f2ae14cbe1704dd3a8c9baea1c2730c074e260ae7fe0460821f67c5bf86dab77cdc413ef7894380cb93d1804803327d9fa0fb50153f99a727e35f2d5143f8702c373fabf7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d39f64304e6f181a14b8cb395930b9e0d9043c9219de1612388505c70a33b4286bc313097e0c02ac96cb25d585e8c5ee6afea3c1c9d3fb7f2a1a52baffde4f4efa1983767b32873f7d42ecf7875e066296e577c3f394059c0a452ba2d2ba4c0870798c0d3bbfa2ae7861c74c98c2ce8c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc0f9d6929e51dbfdfddafd51a6f86c888603f91ff3d401d285876018d2877ee01d57eed653d68e8c2bb32213c7808f48e25786c8d4826b346948bed9b3dc6dc4b2cdf802ffc33449461f4133c5289720ee8ad6720a8081b02dad96b75852ad8071f1915528361ab08d7d7b288a753b98b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24c1725d5fe25462258b4c9ba643b5bceafff55ec23387da076fdb3f4c963f4ca393a68ffa8b76c2276c207a86fe80f4ea0d93dbed535318d56e8c78052bf63255eb7bee9152b631f9ffda9f46327819e6fbc95a059d96b6d3a41ac67131ee6d5af2823c695a23fcc2fd5f9c5b97cada5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c00586742f3c229878747456c46ee6d8f4d820f8a6f2d19e8e13e5a169f8441b1b847acbd8d8a9f430d669da4e179ea638b6a0ae7191c4daf259c743a6a145fa7800e4a544b4ae2294703db385ebe382bd71228ae4a452e053075e2058d1a6e55cd1d62ab03aba8286810143d4eb5859;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h840afc63b60019ad7c0109b29584c1b9324ce43402902e26c08034cedca7a116ae086cd14f4688bca96663d4aaf4ac1ff811326d92cedb40e6da1169dcc3d9efe62d7fcd0facbe94705234f6c7f86ac4c0c9de80e0ec40585b0ca986a02020028422e4a2831c2c13fb811d56a8e5f9446;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b7dcb9126aa6e41b887bb0a4c7cc0e200db78073835506bf34c91d28455363a06601f3c00b063595cdd8e98c6587e8097eb39b2e28b87ae25ede9b2ee266cdf4e76dd365debefda40ff05239aded306f9c00e119ad2b6eb7daf631262ff832f909067804d6e7d7587126831a282b4634;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa03c8d8acecf11354b4a179db7cba1d88686995574894e446ebfcb6b3f2f828c29a80dd646363be3af9bc0476f31b1f592412c320842bf3c7981ccd4b101501ac2cfc923800361b550d49e465c4c2510c61f97260e5eae0f526821f00136438fa368b077dba7481d114f945b8342c33a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce4d9d9fea2a04a37386ede0956fe747b016f3f892c3dad140a17592b1af35b05d86859c044bcd3f73f23bbae71ef8a7a2e6820a53cc62383c4d75850264dbd268604d44b1fa45e3695b6fd890796b9d69a1cbb1237fec66e3a2aa34740a188de1f9e9cf43a4a27a67044d9b712b5289d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7986d4ae1026b9f3b595d24a77f8a39780b07d5d4a3a690225cc1b8281b748d2dc37498519ad954e87adf1d5184d8882c01ceb1d318c493d90852b88e59dd081cfa5b0dd872e472157675b9977adb81df7836ddfd4a7dcedb519fad4385a2dfcb16492769ad0601ac7839d89e5b21fc29;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ba5e903f60622dfff9edad24a629f2fc6fd127075e5d829de3e6c997cb0ab69c2b224ca199e3b640085e4c8961146ce8829ff6113df7430ebb82c765b8443adcae654beaee224285bfacdbfc68f82c4616e04e0bce84341015c735cff95193d3f781c3069e649a4a78e53f9de824db64;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha0f994b7dff98e3b13af81b0e34688bbb5f3bcb42db4c9ef6eaded839198e402c7279ee953b6dbc1c64033c42afbf6769b39fa38c9e839db278026e53c771ceaefadad57a16ae6e9b23d62a0644864b8d1ff1dc075c9f882bcf2cb1127f7eefc96219b67d3c9c76b7032952b4817baba5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4ec9377bb7e6bc917148f070171f60bf3e90944bbfc549f47e358b690efb9a332bdc9fe2391302a5795c7a7abb799b33983e642910da21bd3c175adce876d90b20860e18610c9fd523baa18cea64952575935923bb69d29c2136e09805cb9a0f458aca0027e005aafcbf4d68a31231c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h673ca744d50067d74f05fc5525bdad76a4f7403cb6793e9bad9c4c93a549e1e66e7a8c34bed41f99fb1477a92408a89a20c172fc2c25c05ac829568ca8a6eb126cc75ac85adf965899583d7823c5313451418ce0d75ca62322b1f93e6a9d97803bd69888f27b61aad41a828839abbfc28;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9857d5475897912fdb42e2751c894ac7db4ddd7964c264d67d8a2a116d0e23605d9b1768a2347f7eac12b59b386895786b0e1e319dee5f5ad9b4078d2c8e409368c727f2cae780c2cc5bae478a64ad2fa13ae7914f889c567963af4b9bc02109c11bb327651d65e90ab5364d4ee71f9a2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1484bda48848e9c4c3626d2a52089e298a10dfbe1be00a6eaca3bc423af13f930466f6cac03db2ec4f34b14c71c1f1119bc872b16fe5463d6a655bba0056406f3dcf705ed6679f4c7785e49d5481b74e28f9905359aeadaa07ab16871562f9bf5935273bef9b017e87551122ab4c60b2d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7305324b5f63a02d54895205f78874215d71103e705c2f217cf82791a9fa38647597f679ada42461d6ecdf6bfd61b8a44b7d8064944512ecfa6d03063a76c063f4e42ef3997f3ec1428808d9dcd2684878f873ffcad92da0a9497d89d7928214dc2ccc714a38695fb58f709eabe07c562;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ab63b3b6727a133a2ed174659ba77a2bd1e24808ef60bbc9d823785a83d8caf8416804bf8f0b5744cd4497162caad5dd49eb6f5c4a249e541a41bb8c992e769d5917aff60b55c50df5745956a56149a95c3ddb3ac7cfe15702b6dcbfcf69817e11dfe829ce05969740e0fca267b7cd1e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12c5fd305637502cadf0428f149fb68418dd58f95da1b3ea043addb901698f00bd7ba9f9a083fba9d0d93adaf4f53c13bc01ec45a14bad101c66831c3172ce79d00e4e60d1ddfa08c51527af65c21c6de050bbca8d7316a31110007ac3f1796ce8a62c38ef1aefc98791a42b47420c255;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51e13373279f3ce60a250108cecd1c17bb18311e40bc4151ea8988c7a47137dcff39692e58988218742ca843f6b0409d76060b8dd1c1c7a4e7e8d3d2045a8a5937aa5fd5686fd713ce117438b88c418319c60b9b6466a8f5b1d3e6062921fcdc4455d8438347f22b57b0f96de932aeba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bb94fcad3a608e2b802bae6cebd91470e75182f5f13c2de84b8a6022715628cf6c1bbc28d08824ab295d13660104f1a51f786e3e8b2c82143ab4f295d3211f01f147278156fd08db1f24792c28df94a61fbffd3aafc46bde46746c763ce1e95dd744f1b7de0b934e9a2a43d062806a51;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8a5984092dfdf15ba4d8f0640b9d26bc72fc2077698096b3a0e18e5e8e2bf7b70099139f7647fa9f85d3ff5ba5b2a67ce9cd4e663031ae611973d8b76ddc085933bd693f9eb0fbe418e22067fd364e5a5baf8aeafe48beb1353201d1fcf3616c5097a8c0a2885b3e87a38c7af3051066;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4aba8de0faab18de99b35157bbf855774e593a277bb0d3d8d36f6a30a393b040075ea1740693cfa8881e06c25ae1aae9ac98acb069807d16c88a079a72f13e993c704afea99c76e03e44c1874cdb95b4e8ec5c8a8d32d16b1ccfcbd8e59497adecd38f54a30e6a0cf2aeb1c73fd174eaa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2a6484639c34b0671b281ea550e5118b1ae40be5beab9335a0ee9fb92855738bd88611b2c58f6ee79ba084dfe7c118a9135c8f4b2dd0222fa7eb4cd3e8285e297687f7d92cb7cfcbd2f2f983869fa29bb9db5c24b9ff539bf09a1962d3b1c6c375a4fdbd07450e57ae88104691425554;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha94c1eaaa42eeae18c5d09db8f0535c8680b4b55a4f0affaab332f7598929aeb3cdbdd355942082771ca9a9fe1301b8c56ae0cd914458689c222b711a15ebef865007eea05f94a491c96f230b2d59bafdfcdc2d94e3e4f94a735c3d6e1c2fe0b8082a144c8d50d6cd5a6cb77a1eacfd09;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1a5a5ab84a1caf7411d5251e3e9f7ec631b9f863a4732921806ec9b1924de56dafc7b0a8f6ba118c4fb7c4b960fe60d6a21de5cf10b77fbcc50cec7c5941a719cb3f172df5c78a791d7b6e7131f04f413410d42d013cb4e25e0d007f1ac0ffc34f4bae2af11ab742db15d7f5834d69e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e80aa61ad4832ca8ae5f1f727e6f701062d208a30043aa6cee7a0ce5e4a6396a02b4c5fb8b70b36a078f463c34adc54f11b2c2a55390324dc25c1f5bb4727365f6bda6ddbedf0b411a52a6c3ef7216541a1e25073e8b07153c07bd467c080840b77207eee6794f3e2f2e44f712555fbe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88748929a98fa5c05b8ab5403db829facfadf61d1c0eaad62e0c79a10417eab209477b961d69cffd9b2afcf256f7eb58a85bb0dece53ed8d96b675060dc3c7c4bfd352cc9841369f100fc0dfd5c4bacb57f49aee8a410151b01d72e6afae26b7c7df7b00fe84d54bcdbeb2d366b8e5500;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48e2d34bea081bcc424d7d6e34386ecb74d8f323bc74d4159e5e8d2bbff9bf4cd0f7d2c8d5e535b82fb57c0bd4500278e08403a4fee5cf1287d516f6dc678a45585d9b240659ef69404b667d52be0abcc9f8d4c1981211aebe9111e488abe3bf292e208fd1d953a341075d2f5f61ff554;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92837d1cb865edc0318af8699cf68e2f0b279b37b9fc90501c1ee4516859145f349de2071b1f76ef2dadd1c58cdb844931817f95a9c6b59edf3d72d41affa83da95dfafe206414c722fd1889b33028622096a41b0a96ef3c7d801826337f1895ecff551c5116c66a2db7fab31320c5350;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbaf22b2378693c84c9e5a6a0fd43155becd9baec54ea25128760fbf7347962040d16cc0740e8a342d6617d349a8629d5e2ddfefffcb363afa0ecbb5ec6c52cbc2d27690a40c541c0b259e3cb91b5ca30ba0b1c6bb32af5133d2d28daa7e93750842a2eadc9022a72047c6737d91e09f78;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4b819f87855c471a05a462f48320ac51e6e6e6d95adc2fa35a45b53ee4083c5ce569f26894c57042324298831bc707315a89fbedfae5ea462d10d36939128a411b838260288bdccb0ea11c1bd7f11f369413bfa10d36ebc7e10e3c98a82878ab3998fcfa9a8e09ce62ef4c75afe87af5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h575e22a896805c1a6ce48aad7b49f003baff8a2f355c3016a79e6e9b1650b05f60ccebaff5135bf724214a8822e8cb55f1ca9b5201bca897eff5ec5af847d1fe41746546562d3d587579850c5b65162c17b8d0189294f4d088e88399985be1b2fd21e110b8431371d219fd46b380625ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2897fcb40b5ef01ec01fda9a9112e22d4a8b7d743c4d206db33b9acb212d1d4e9198a491b65929a5447ea882a428b70a07a4da6389a54c0a981ed9a7f7641f8d5fc2bc4959723257a562c2d5edce0c09f2fb02b566074dc72c629b5e0937787edd1d609f997bbe8898427737cdbedf35;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c78d23459746a99615cd28084e7de175d0064e1f6657aa74413c165b20aacc29c79218dba29b648ebb89de92a42c1e33b73fbaf169dd0b0a7e00f01d19ac56b7e77a1c254f8f1e4b635a3c30cf2c105c397d9552b87e86683244ef6417113435e984559724bfcb4701ddde387f3fce44;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8497b333da551671f8dbb8faa5a2dcab9d3106f43f07d901a73d642eb550959782979f31cf8056d49687be12f118244b7d79caa1b3a88338f2fcfed2c64ae85e343d7f022b1bb7ac92dfb9780df7363b065f272d7d4ef6cc168510a7f1d3cce0c8aa67c43bffa2303b0148edfc68a8b68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f8e867d2d86d998aa62435eae853136786098f2aea10769cc33a2eac03c1229fc218207b1eb70851b09d6bc83148f5bdd578b15b128ca6d54d4ccad85970cd172e096070d720f1b0932677f149d20866538a864c0c500d70f4eed3ad57161d1d669b89c8dc3c8f7f4b53c714d710a7e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha45701fe02ff787fa608aa47c440e36aa18064a5ed6bdb78c5e367720f576dd5b5d8af1842bfb4d9fa29cc21352f163e5314740c73b87b72479fb53bef03677030e80d4e9e3e20e84be3e5fbbd3691b5116be0163df4ec71ab30abf510918d46888ef42d05cd8304e09c610e16cfd959f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h709541b9f6dc84b7fa8eb254a3127e358992489d0de6cbe624306fe47a26746f17bb94292684d88fdb042c866726f1e8ccb8ee5f5525641cfd2b37d950d96246f04472a9e37c053d74d44a2a6dc190c5584baf5d52dbefb1af8be2dc8f784ce9eefe5472715f31e31a3bfa9406127643a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb624c0cc15d2cfbc9db3c1c69e1832b7419e962c198d8752fee7052f2ff515fa7a6a9c8afbae8da7ed3bbc4d28dbb02af801f835f48275c3189fc15fed3aff100e97e36b21d4e2563e21df1ce70d7bf5270ae070d16848330dfa956eb93e8e2f2c8435a74ebb20fde5c279845a4e4ee7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49e540a044f7913f5bdb67189ef022e658f57967c801992c6e7f6c65c1538ddb5e7713b69b6ea2cabb8616498c22bec8420e2111cc926371f9ef121437411e045189d61dce7448285d3a096445d8b3597cc5f111309820787b9df6b2a20122095fda2bdedd83a9526f9f6591659af8557;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5bd43dbe7e833d21841d853b48273504cbcec6be42fa29ad330c56add05495de9d1da8e0368c1cd760865bc2a2deefff193f3d5e70f5636c82e79f9cbf54106062e0ad9160d72e9065e07a11d8941e704a5148b512d5876a1746f5adf82b4ef88a111e5829d8b4cff2ca7ba8d07605ccb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccf284bd7c685fbae4ec3ccfeaf6f64b57f9777d40323738592aaf1d8b92d4e9252e104a945aeb7e5c3ccda85fa23a650098d805bd06d7c9d3b5b296efa00e7a7e43f686d61741be9b42c2a2cffb0b6804bf8c1354f6ee132e8cd811a89ce916eff97b3e5aeafc85350201b6f99e2494d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha45fa76463b1f48611638fa7d124232ec811640b97cf2343c6decdb055af0beaef1ff70a05e1de1eb5d7207c2b2f6f2267a90e95552870302753859246d3d4fbb43f5caa682346d8ad9dc918b617c812e5cf120005ddb44a1649f7a9ff42f36bdaec1b1518d36b14c947bec5047649436;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc28720aa8d983d5f101b305d03003c9f8ac76ffefc94d5c3bdc9e7c6e1d009b31d0a33ae79544077b4ac0a95c674710a5416314d1396ee8a2c65dd2a238030906c74a36754e6a7825d8bc8c4c75ec11fba5bb342b76380483a95b3a96be36375462385c7eedfbcccb133a0c596dd34c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec4b38f97b7fdc7926cea696182c682c1456b9a60d01a85282c97c672b38aba7a5db6bbc10ddeee41831336c9f5fd4a3248c0109df9367d5a681832debe4ee045a7ab68db2d885381b323ac3527b6501221f537cdc70a9635dab75c7023263a4e0f9e70ac5b513fe14767f40df79b576c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c5679f0d3a41e27a90b4e67661a7b9446983b20e7c53b9f49b3665c8f0cd8494be84022b96441aeb0c7851a0eec2833cdd37c1dae2fc47713ddfdc1fa94c9b4c4cc8428c164731e0f55222ccdb234700d0b4b3edb92d387fcc2535092789eb1f5d551c7f17247af25da30fcf674a7394;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2879cfbf10fabb9142bc0a2c8760972549af2fdcc0cbe37a57cabb7c05b603fdc1a1d4dd054b3f6cf28f4e159b110fc5d48727727c877097fde27c591b8ec7b0d77cf4dfdb648f32a273b3db42456f1995c4be34535a6e8e9adadc81b5aa420ae7ef391fd4cec3d2a4d9c8932a726b889;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8941f4ec092c30f6f7ae68aaa0b9783041c35924fa3b88852bf21be53b187d31150db9d15414890357b07c581fa22a150f65b6a838a9d30d7433c2df515b24457864e697400fcd463e6e8829a2edb3b889820d761c5b1ccf3c262e449cc86d806c4395a83aca490b340f9f780d4ff7fbe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4ea93485ef698ccdadc9faac51ee00010dd1af5b7594aa57f77e622c75c17119dee91248315eb7016cb67bb4b830762a2ca30750f616d0395120cbecd68398fa579c4a06248b4fd5997890cb11e707629645f8eb643935d02c8111ae35b9298d5efa84d6420c234a5ca5fcb26d886901;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c333bd24ffbba0b1cf6b67223fcd4dc4cec881c686b958ff91302e8955146a730eeeaf9f3a7ec466124bdf8ebcc1f6c07192898bf6772a0e6b50525bb0b9ff2d6afa31ba8277e0fb9d9c659922c1248c74cd5b691c00944640fe8cb9c97b38f8a9cfa145a48b54d553da27f5f0a0596a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42272b43010672c2c16ac970c2c91d235115e3abd584e071beac522949793a6243e77078b31b114abaaca011bab772cf92a2d2864d41149f8a6c1b3f0f4e4294a088fe0b0044ffaced6d855400debe28dac5d42b9d66d5c837b9d649573a0b728992305344702bdcd7dd23518997e93ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h899271ca4ac034ff6deb446dfb783c34c7e4d8902dd45b5ffd9426b32830b24e20829d3d8ef0d7fb7ffbac1f471dca443149973417686167b225b511ca74b982ce419b800bfad29580081ccb83f118b638eb6e9202a08c822005f3f193c87cc990124a6e8e78929008a68e169198fed39;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d3e0df85badde356912225dd7b7553dc60d060d6bb9edcdf9d119b0f9188c583e6c8378c7b90e25c04508041a9f4eb4544041346026c133ccf6d1bad1f7a3cc9504a4f7f15bf134517ef9750fd14765595b525756fea976569e87762f6d0090b248bddd12fa497911857c1e663270aac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6b32c66c0b69ab84f01de65a4cf1ca148ea3f25e28574f02d988455140d3f0b1ca06102bf49ab39c87474bc91e7c55ef165f04d2110727f6a1c4319028a8f3e42df0f6cf2f16cf4ba3eab30193c48e983a032c9720b9a95c10ad66d01e59f05b864f62c5501674cf123fcd0c64e319f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebe4c24b2f3aace28441584bf7a5ecda3e72646568209595c81f4fb050648134cc6a42657330734d9b0e41c775fe45131d3f246998868aab69f5cf124c4c47dc9725c267844ca10492b5fc00d8eab78720b8ec50a20d01734db34556a189575586264718e1fadf3ce2a591845b0b0e74;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb1d53f5f43f559f43903890e7d078df035b774854253860a4ea760f8179d1702491263d5b6e070e9b7252b2f4802bf4b659ed55bcb71f5d921e613feb9bccb17f1ff7081e02c7d6b96c9af7a8c41e2c7d565aa3d4b06749fd51b36bb2ae54d0925263b90b327432fcb76d71ddc3d4b79;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h926bc3b590d67afbac19417cb9bdeef2374e7e06f6ecf2c08582ecc8682b21160948e3ee6400c9e776f376d0471ae121d685c9d62145bc62fa9fb46b5eaaf8ed1ddbf7e1b33cbd59a2069a8ee7a8b893005ebded792e69b9056026762c0419f6a06a516f70636bf37cd067604e6502554;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hceb5b0631f5b9db7dcbfd3c80fc7efb1dc0437ed61372ee1097dd1ff14a43744c4fe94abba9050a173ad33d498bd64d1e3c21b97d9967c36700744fbec758c894cb7e87d2bbc7b77fa7bbac53cbd20c9fdb79ac1ea5a59688197199818a09d8187354a37dd3250089c7be6076dd8ec97;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89431f09c2c6513198f780694142287d0cb090677f8354cbf4d2666a2d49537e16c0e2dd802dbd2382568e57de8ec41979754706f05493650ad6f97f1c2e1b56a12cd310f2fe07084895647100d687444e243d33a43138bf8d0c32d185912d106364a0d64ef6658c02836ae376b7aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e76857e5708f140860e9bef18c43d1d48f33ef5259f032d0401e27fcb00147f6d4ddfc789b7435a2f1548fea96e980b6d52ad4624aff3bd7241c4fdd80e5d2b1f9c1c23ed9f650907ab94774ab92a3a6a90ee8cb844d34a6436849f21f5889124f7b6e6441a2802e2403932bd453e943;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bb0a7326175039196acea5705a3e793597b6647fa21d66ea0a12e4db56d843dafd4b76da7f3918c4a353654af8894d181c66d1a87c0b3d73adfbee6d49ab804ee1dd1c3a870107e5742912617a00fc7ef506970c97d6a1a187b3a6cdb6e65d86389047b1fd74bfe31e25c01119ea822d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h772c27e46305e4aa46b4357dc82dd94f2aa08dc7913bd361ffffa3d06adc90c54f025ebd35c7f78d40759b8a16297f69d559a681ae349b69db48f27d34e607a5abf3da8b7c3c660649d1398b98bb39614792888bdb0f464d7cd59bbc6633ba71f37f4807e8fc9e2d5c5e5e0211c8b3aad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb45ec2426fc16c56fe021ca115d00af2639ac59f56ce3f855b6df250309043cd8c8a6463437c1f8059730db42400e4e8729dc7e756458a67b6eee9a1fe40649d33ebca2be889912d16f561b9d376450111fe8d7bf61938c795ea44ac02545441126407c4184f35833abaec587af10f2e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd042c5e29e158f6937ac2b3459fef11ec68d927e200d566c607e5a8d5b3b32b92eac2bc69bbc4b735e67075e5f368073b4e0c11d4fe42a3fa86c13c4e9aeec1a206471545925354e51eee08ea1eb15068967b98c97f8d1336ed34031f68b60c167f148f6aa86519a2c01d500a79149ee0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb5bcf2041162cf65e248a859f163064abc4933d375b0f18d2483a315abb65a05ae10a389a38f8e98ba89b9010eee45df894bc87469ff67089d0693b09f5261d8a5976c2c30a77faade54780e0b9d24f94279f58e3afedfeddd418b0647be2a6d2ddfd1fc72ce444c91f995e2d6a2f067;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2de05d8000b27ed2e7720fe6f982c0c1c579d7f242ce4e86f93ef3ab4b0c5110bf4e7a22035afaee6c4a66254fd1b7c886abe03e53888b12786c503c823081619cd9a94d15de86b87838f703d5ff73223c474bbae50873d4d9f89cdf383ea11e0c1ec932a39c31ecc875a5cd97eaf738;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bacbf5a6a483835b8e96f36169af565f53bc1e7bd7d4c100bad24fa1501444c5e3d5a8e318a9f25351261fe823d78e2f04311aeae97942eba35fff4598e2728f035f5f8aafb09b6d8fa7628f00206575ae0802017f6cad1703dca47e64e9b402ff84a5dae262981ef80af68657866054;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b2476c1fb1a218a9b80f250436a7707ba23dc7ca9dfbba1171f1f92c7b793cdc5efe54b72a1a9ddb41f1bddd816355b1e106465f4a9f7947b65a5aacb344a4028466965ebc7d6bfce1c612df89c74592fd921772aaa475ea31a88c7abbec8b0440fc7ba4b55de5b8e7aecb89925ab1d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82d05635ff1d38998f2c3d24b4abc0d33420c66d606a5ddbfb87ec5ff7403a26ada48e60c70f3cd18bb57683f13672216689adc361e9f9dfc1d126ff15b948cb94fe805c51b3278b62338087107ac992edce78500a90002f66679ac66c671fcaa296abb81b770cd504802140b76cd5f9f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc81a8ee8af6cbf927bba2e8043380d1c3a7bc71244be7cf91f8bbe4b3263ab8f038bf0e79237396130ac368dc44f5fd6fc7f97fa88060962a8f5b451aa6954180774b2b87f53b7c7a3c524e6f8748362ffdba7da035ea43835183609bbc8f719184611bc531922814e3d63f22c6061bea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8fca168000901938b889f793eded97cebbcbae17eb30db63a0c17bb84a2d276c6bd4db055c5871b69b9b3ff78c9952e5cb3ef63550e4cffc85abd7a6e482d10806133dbfe0ba1acbbee4755138ffffa0259a93bd17b88bb81383291ea1448612dfadc547d0e870adcb6edbd25a00fae82;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73e0f43ffc5e0e861ee8a0f14a0ec95e278556a1453d2030867438cee0285d4a29560436e4ffebf608359a25227b91d710693475e454bdd1c6f08f17de591a379594c41688ab4f3b0043d05bd99fe92546bb1311899d170f28ee4928d2635e0a76200d573ce504e10adeaf21973d9f0e5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bb8cb6eafa0807ae3b6a3a19a2e4ef2eb3149e536848d131b677403eb7e41cf924f7221b588d0fc640703692a3dcc5a9e582e09d3c15495e6ca0faf4e8759b47702f9332f03ca5979ec0a732e20a28059539ddacf027b632684751a88f07434b9402a5c635d65151f8c64f27116d32bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38afd95ea14db726618cc51da63aa13a2fbe2c9889f81c3b390e4aebd6c761e085837ec7dd0149dab3819779cade9860a5662596ae32ece3442b66a6782babcfae488f7bca0bc195cfb8a59ebf2fa0c2f21d14a7a4a36b5b58a073b3994b22e2d3961f6fb6292d012806b3c40e6d678fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2019fede691057740c863844ef62651c96ee3901e9ac516f59cd5ecdc5d7e049ca255aa8ab9537c13622c5c3e99a044fc12ab9d35fd797b93b69af7865cb4e3af2297865531977a95076c144fa343ebd65452d54ce3ce0ca6138dd1b3bdf2153b22b3f759582c8e0b5ca084edf9f6a8d3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67b84bc41320ee142580be6498b398695a22cbe3d14e9c6d7a09b7f21801b23fda739db6949e228a395e005431edb87ee0194decfeca270e3ab2031e38a585a25cda56c8e06ed5a6a211e95891da93b51803d73fb7ed01411cb2d22e10f998b2250580f0e8be5ff66f6311210ecc56aac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3236269a1be49d156e9fee5a76f701e704882545c4f6a0a75d85f63f9d4d34eef2336392cf6e438cda67f86b0b79a002a3a5d3778fd619ec7a3999263699dbdee4af3475828d613b1c310570360c71a0e225daae09699f30fa645a4f84b36f13c4cbe23b2b5a2e89c4e87949222573ad2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9840670479fb1024b9e90ab9dcd7bd1699990a17a68873b1aa29f202bef276ceb465447cd8b4be66a8b218ec16470ffdda55093a90f0aa053942dc1566264e3ef9efbf32b75c7b7faed151d64f8b44847fb24dd374cb5b113fb73ed19d8acc5b02fbb91b31b28b27a1e69c6358135b33e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h881e324f96635583833b161aa752ee9b84c66e93d914318496037644d5c76cb33512c799667a314abb4ed3a8595572f15ecaa2dc8a2ea6547b90c184423c8be458e5da9915e9db12cc61761e0ed3aa99297bd1f4e84cf24f986399939d4c29ebead50213598dbee5dc60f7f155dfc316f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha055d5ce991a8f799c6991784748b4202cd87ec203ee75639c00db9bea844c182de51a27dd8a47a9b4fd1e0fc0c6c57543108209860802ba69e6ce0706c8aeb2989a741dedd777d85b1f5a20cd08afdbb230719390ac13d010c52f9948656430fbbce75449b31106db4e12a2223551b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd660ab264fe571075267d95c76bb8366866b6d0df72ef7913557981511732ba047aa725fa24b4a6eb9d3f7253dd4e8ef6501f9e378d36f704df2d470d1166242a40d8d154ff144de76b1034c7fa063f82350ec70334b55b6495e301f47d05471a411ca79ad7196e6b500b77b9737cae87;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4054896b86a46164df09b634e0cd8434715fdc2757505a23774c234f0771a37e21c870876b2e013a6675061160185130828dd1610e7e341d60f55338d5bca68ae1fba644ba8f1c8b0691ebac3f26fb990d13493fad1f598ad8084aeb3e63305e899261ad1ee110e92f4d42c6f759cf03;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea8f71db6eddf6789968ba3500ed5484173097802356d1ef7baa63897b37f79c4edb0fe135e7d38bfadabddb5fec3e0d5975b9f35ad231d296344be9e693756f6c85a87ffcd94c3460095a41d5eed0b5f538ab71e2ced5796f66917a7edd5d2b135194f340e310c71714d68a634c69b46;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5b1e04563257d7f3afe07ad39bcf56e1fb1c707d5a593029450825f0395ed212f3cc7c3f61457ac809f1bf00042912fd9b7ff00acee21fcd9d17aa79264a70f1e815221a49ecf3ec494b9bd25c8a31c6b58a1332f2ab4e23ecdd0e5f56edb7fa9f4d0c76ad5b46e17e4ec43d7d87770d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9c965a6a34bd82302f14c969b40db3b5705af669f619bb34feb52a7f3a98b6da973bdb2268ea945b54b173816256205da494149ec0aba41dba47620345c1e314dd2e70440151aea0fac2b77f00a6b7a231d8721345a3847033ac4332dca61c5cf2a744c16302fa7c4e8cd5017dbd7e5f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2462e661b3a25d49acd780f6ea1329351788897b8d12737ba98a1f6112b69ac7d2786845de9c921716babec887ca56b51d823f6fbe6a0608033f12387978cd9bf3bfaf73074152b4c0ae3d238c81f15da87a9386df372b3666c295adf72265901b0d330206857beda64bf6ef87328f11;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71fbcc158a909eaafeda2ce81dff7f78c72828c435570431fc0856f2ce0c0807a4a507cb3d1c74d945116a27ce5e1e9a5792bc13ff482c8e40a99a3eab2399125dc29a312d1f17cb50576b0179515b5c2ff05532abd4a2c426cf52d62c43248e7584ad982347b1b54e82ad212fc55ae4b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb09b2ed20c2821daa15a83583cd720c646ab2b125488a3427318004ce43ba1ad2281ab3d8af8e9424dab310e4c4d3d230a544557ab30da305971a6ead2d96076d6a16fb646d00bece79942c054762fcf1cd5bfc1ca868b7bbddb553d777849d2a90dc09b7d0c097e9a212ac15709bb1f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d1df522a152f19008047bc09a2ba173e20207175d868da6f0b0b606f2f2a53fa09b8fa6ac67dca55e1ed8169187de1fef592d1fa2efb12541a8b0b49a1b217427b3f9e39cc0ece81094a4e106b2470b6a1d166543ed57901b75dd10665f207201225562ad5560ed111652ef9eae51b30;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3f9ccdedb7f60df6f75f7dc5059d7f307e039328c82b5d9ac662b12cc53536c17b3bda6dcaa74344e25d86edbe9d791687281b4b473dbda98ded6c896cccd42950581fd8765da8be9cd20e2b2534ae0e9431b1b35add27e953b2bf34d4d76e1a033c5e14f2afa604e5f58c04bc5a5977;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h622bcbab2dfae4758dd4fd23a0715254abb1d6254ac2670f234283b8e2fe86cf726dbe3f261f6c05fbfb1701339da601182f17242cc1fa0630b1d506f4b8e71165d97106c9baabb4f9f1c64fe632df4533426dea3419dcfc7c3286031f014dbfd9fd5a372b6a421461d388da77157234b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39aba3140b407ebb93787028708edfd00c1345b12c3e36ecf4f7b383f785e6a933262329abcc4b3e46b7c4bbc55e5fa0e8da2a3803ffb0e5da19d2b7ee92d20dd8dd5cf11bbd44a9671a29830fe22b2d2beb44782b8a802edf2e5d644903678a9754790c2a1555931cabec7a78283613b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h151b22e05b7d380a60b73ae3c9dbaebdc502ed209f28f6212e88c2a5cbade852ed4c14e719324c720b8f04215774671c2b44c7ed8e31cbb37b535b4a91f64409fde90f6bd0867926dd4f8e266d6e9ba9f00d453c782d41f9eb1207726e4928aea9698b31bf292dadf019c935e3388d078;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfca6ee8cb3cdc92e0ec6d183d5663cac4e7116180e549285be94322dd73e54f767e113a0ba41e30bbb0dd839e1d7546fccdcd8275f9103b260969f375c5cf69dc21e14e2e52e5ec673e07d2e361ddc39df17dc14cdd917bf4187b4b2ea132a06850505a39fd41faabd6d037028463cd72;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9e908988c0f09b0cdbbf1d0f20ff91c931c136c16636e879bb8c3494f8459461c19bb740b3acba4caa44d7a91d77c7c73953e3c5d95aef7e326e5ab234730faeeadbaf93a30d59bcc54b6eda94bcec7abf9c7340c9d93da92e65d748c4042dc3cab1583bdc7cc6f8d3ae23a73012c590;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54e1e8797d9ac3f81f89d424ffc679db7a049312187f51904673f50cf103a3ec61889dad5ad54b18f1e80e1c859b7af531f12ee273efc74e8a9f2715b7afe6a2e521006c87da3e7d1e9927213b3ad87e58037611bddb9ca1da0873df2e401213736407fcb76d989de1cab08127668e6e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ce88451a5babc3e548c5664e673cf3697bda8e6ff4ce52ad3d9782288ca44de52d16f1860013752a92c68055e65c13d7c8aac85fe9f7de08438e5c0ea9ab360f1301c541ae4efdfb4649036fb62bd232553df972cf361eed587e7d6edaf019ac1ab46a3528b6495c911f963d2691367d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h450059eba7cb47f87dd74817806c7e1648c05f26b92b1ddc5bbc2c7f73290192369b23677153b683ee47e1264e2449ed0afe6d78209433908f128c4ff0c66917f9fc23a5f572037561a014dd4a168574ab3acf5e741c0dba902485ff0f0cc98789e4edf213cbea5474bf6750a4e75e503;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d381797fd73f7ae57db1121f4b784abc00b4ac5b817190867153060fdfead8be87c336fc9f5d908cbb838422fdc891a6f0f9a0a549e8405f29260fec364a11832b32f50d95330f7cf8e215e1bd90447c4971018d836002a601a10516a0e62b1e9c1d02d7e43c1f3c8ebe90e1636b98d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he540bdd35de5735360b278a0c54d7e95a21854b64a5e898a65bbade36b96d88ce4f59114eb762ba13a8a3c7bf36b3b41a554b411a0fa31d261e67393a333a012dc07f2ec6c6ad412a72146b77a0e11315ead182a5abb3046616bb8100969fd378462a8aa35e0ddcc8a887dcbb426bef14;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c12669b96cafd6571e1fe744ca481d858d6444c3b1f4c858dacf223382003d5838775d2d1bd7166a0c3987660cef17a202e16937d5a2d9e9086342f528458654065cbdc32079ff1f1ecc7aff62fda06594c7e0c5ddd5e76af2a6057598fa72ebf30518fb2d5a822bb5c2b99b259efb38;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7ea5539e19ebf4813e9ddbdfe748b1834cc2313cb7591bd2ec39215dbf1680aa112cfd57bbbb7fb65f38e10a27698935418f0fb2dc416ad18a5e302b2dd9621715acad580bb19c4bce52e8167d6d2b54a6867fb63ecf96c8531fb5fa0a7317b215929597080cfe1aa6d203bdf914d7ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4d4673beb62f26bbda19776291f4df01d53e4e9f5e57af7b9a298cecbf43d629a6bd1abbe37292f40fd8ebb23bdc6c0b4a3905569e8c1a60ec93cd6253ab1d1e55b8588a4bb23f8ab6656a0d6a8a7596030171f803cbda2d3e6538ceb65cf05f251bcde1904beb04223206e4326fbdb5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd5f6f1b8b22fabf4a5b2d71b92bd50829e23b32746a49f09c174f634a4334622e6f6b8d8ed8650f3a385f24cd47c389b336d6d726444651db1aed4729ec303ee6568f26af0360d8f3bd4876f5080d7140a144aa3d5881a7f9298eddc73dae7f84b1d839e440d4898b3bf4c25541c2823;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1324ff090b2f9883cc3fc8ec9a25652727baf4e499582ba526110f3bcbbc25f731a722fa0d7196f4afd79046d8ed8f72170a0b7fc0fba7951c99824c523d762489c96355e9005cc8515cd6755be8c8f3c035246f454d251bed636970c9c9ee6bcecc7cc76d2bfeb99b1f9a1ef52dfd832;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h182bcbcc1e264657f2b3dbb8f18c5c89be0c5bb4db35f4cacd4b9bdd09447fd6929872955fe94bc4bf404e94e37d86a1434e412e90b8bee758accf342a55925eaa71917d6c3440ff1a9e968c462d09a4e09c2b9e02b6b8ebf8465960d5d9da7cd31bba2c9c37c8b09757a3a067f2cdd32;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f99044feacf5eb3d415171a82d646da6f5b42e65fed5cc86839ef089a997e058e5d25eb9c348188a5823bcaa8969008d7728218e7f44322002a0b96a289e8c32056c4d3de7bbd6ea0613293887b70baed9fef852f29df42acf590e89e178f60c1edd423e63ecf7cb1acf8aec9fed6dc9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdafe8d0d678e983bfc2ea7ae35477736d0c3b13856627b5b2e84aa72ee7b82f0e6b3eb0572335ec6869c82398de1cd2d18511e2a78351a23936087d34292d53509f74d33c089e8e72341d8849209e1655e8d0e538ecc6a01eae8c940fdf882795fed4e7ab2f13194b0c22fb266f8b98db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h869216795725ad8ed9efa96378d8857109b39fa23a35a7ad8b414ddb1e3dc61accdf7ca4c6675534170326a47a6070160bc3acad716bc485bc78d730cd2add840f0ae0bf3a4ebb2ea8eaa6b170b0c6428db2ffe783f888876f870293cb523bb1d695a760f4207bd4614e49d072caa08dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a0f36211b402d5c87e31753b6f4d2342a4efdbe9041f1ad46d585b6377fb68d02a9c9de7112531844099414a40491b3e30931a99ef7e67ea7016dabdaa4742c47433a2d0e6805a91b8a56e1616c6876a6f21cb51c309c36b078ddec85353a0e3b000f3b35dfe6525bec7afa48d4fd38a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92844840b5c620c71cb0b1b4f5a6c87025b8887e80ddcfdbe65463d79b334895376a6734736b452e3bd778cd2ba39ef6bbbc003b795b58428e24df8c530d1b0612e10377b7fb3d1e356ed3105828c2981d32d7fd6a9ca8efd81a440520d74833e0baa700999174ab47da2f977c6c40d9d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce8c072378b7e96a11444e5f646ae01863b532d80cac853be8e385e96272df6dc50310deef40df70923767a6d3b1aa39b36a86fa8d7a94d73309b403a847f7e70f2077eb5c3c5ffc5738f89284d280e64d01d499a85714ef83dc4e82bdeb50b11dcfbe057f63fb98ddf32fd97df36f60e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h801d572b79796f9027619402df8548b4a7c702c95e4d4c2ebbca5d5fe98e4e5fabd302fb45eb1d3e60a73f82eec4ff80290fae957e2d4169aa17bb6a677b2429d7d37c279007221e03a708f672e74822320be84c498f8033b168c6b102ebef39bad9f7f5193f20ac3a6018171651353da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf6a985f2ecb3d4dccad71f6d69e3750a1968bcdfa49d605b623db2ddbab670b85cb3c770b8fc97f8b69009e6e8bd9b2806e1201018169256d3b34d4938b4939354abfee2cd2f8b766f1bf32cd2833bc1d15c58f8fcaf660506d345ce7aadcc801bcd6ae3b7b14967660307ad6fe064df;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6271d6eb1cc95fd7055c96ec67732df81be11af533a4b1fa3aed75d2301c090aff3ed424ba6e72f89b9e7715c115e2687849cac86abbb0cc8d43cb9f90c2c7a33683e45938b391257167159b6b033358857cf9ccca289636a1e4365ec8631edd9228f99cb6d6842d7eedfeed1b68bea12;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a355c8a02fe7eaae040391511552cdc69aee86c83933ceb488da27175fe9e9a46f28922643f996d0d9adb32abfe0783b4c3bad63a1c56f83918b0a867009f64fa784c86276675eb4b8f3b00188595b2e272bea24cc1a3751309f4857283f1091a93437bc40a4ac11eb183804e3059c6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65b9d6eb0fc97a219a8e4bd7b97ea0caf1379a68be81307a558be183bbe97a60751258c397ae931e0d777e7ee555622994b0ca67d08827d435626007dbeb99cdc676075a41b98429a4794e1ad12aea5bc0cdeb3f155318557e6edbac97b6728fb85c529e17b63210de0725ecbadcc9ca7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha903a72fed729d63bdc22b046506d9b9254a74c8d76c3e453220b3f107d12f7132ff190d94944fb33660032b78ba768555f99fcfd06cce42146f8ddb79139a2efdc0619356f81b5ee47927e161cde41b62c68f77d249f57541279f44e0a69865cc2ff1fba19ba9f764ac413a3bfdd27e6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h107aa28114b585f918c6099867c2bc8406d01d834fedd241504a14ca59e1ad05996d645b149c67fa7de938ecfb734d13cb4ca1f9448d76449551504db0de0f42e71c12c70474f07c91a403eab842a938bc6818e68517fd9166ed3b006e2cc1a429fb06a7a073170d0d6c9ee583ed2efaf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce2520175117758df52308287c75318129a40852dec9cc87b35ad53dea1a4523b0bb9d9e19479ffd9691516b1614e67157e39bb016406e2a819bda61c1da7a6762bffe994359c9f7bf4a161d0867ef58495f75f8946aef13320ea4ff10c2e97ebf5fa0858784b73c02e3ce549424d152d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbccf88fd087c411b61288c94b2142b9af38b9bb902a466b4be5c2e9f68601716e6b5f652a0c43ef2b820a0539678143430769a5a937142cbd65be820e23ddca74af3d6d013af768f47aaff317c9368090487cc18f820f67b084e662ff33940088f9e95f67e5dceec72f25ced3fbf26d76;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9acae85411131df49fa232c41265042154525d7711f2fa0d830d11efbb0923e960f5f5eaef16f91b59ebdade26389d41f779fe0bd52837659a18a24a624706da6d8af979a9b99ca4fbfa95183ef9bdcae09f9bcfd5c994a22de44cb9e7bdba08ef00b38bfc6dbe462d0fc1ba398ea1330;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74de3b934a6502ac6494f40c698e91d4bc3dd00c5c953e99179b73e2542b30b84d1337c30ff5fbdfc36f1a0caf5d020b0b0e55b7d5568ad8b6c2ce800b26bb5b15342d3566d23251149a3744d544ef00298b2092ecacc64cc9c1b0d940d7b7a538cac69ff1542571ce9da75a42fb7e635;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32043012099edec9b7c7f68de9a5943798d985693c9370cb923157a0f6faea5eaa8598aa19252f798e2bc446bb1de7d3afd6aa5e0c332511e7d4eada94002a4d7abe54f9f107c81cacd4daf39826fa655d3fe6f82c02e9770cb1605fd525e5654894de562d47482b013650704e8c31e7c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe545541c6c3c494c5e16498b15fa143b2416dc2412e1adb8e6f4e5db6b31addc6047fc6c41065d797733562774a3983f4e885da34fd50bca1066f98b318aaeb43620e5cef878e6594e93d959ed7f7b9be88361a7fc9c2cf1a434636bfea1b96f2af6be998c00dbf7f31ce77c8c391863;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8e1290860d17a773620f5cb52df578acad10ef6098502233f8a1421ffc4b37ec0ee5b32043e742bfb619b3f33e3c9f15d52bf9f2e217a584ac51920bd97e9251a0eb5f33888027235df08a3990aa69b61a26dd287e263b690e9b1ff669a4df7c7c17a0a79d819a0930cfa570c29b63c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e4588d8010d388a258c4067cb4334eb510b39b458dae265aa0e396035299cf50706e217fd79b5f821ab6a782359bcccfe0b3c8fdc4202ba29b3f67c3aa60238ca0a69ff23f65dba0f79da8ea79de76cec11ec5922377e729c811d9febba42877ec85aed550e3df9c2ce632c3ac1dbd0f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c4424e56474c61d207446483065aa890170d608fa75278f8e14b7403ede623745161dcd0e48e5ff755a1e4066345a5d120083e9668093f6e7b22138f0fadf02c403bd1a39d885aefed2790319e7f33cef781ebdca81ff56876db01ed354ac07079c529514c607e3d3789cc4e0ee88773;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c67b1dbd4a4cffc4a16d8fccf6d2e2f5e22bfd46d1a81709cb7a720d4a72e937852276632861a7fd39935e5849b1b8cb3ce3d69c4a8aaf37bce565167a6e7aed1fe4196e5ec3ef794a24f55fe0cfe15c09c9821092211bf2ecab5f6524e63141d7fb88e74b16bfdd958a5d0e92970373;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb0fb29020d7858be7d8fb928f88c17a50c0e0003d8ab66934004e8f8452662c54af40d5845b3188276e3377d0ff5a57fb43dd6fd71d8ed13bccae959e43dc1f304bfd3e830d41ab314e829effb8d4062b1711ab03060073784cad290149adf85efb9064e7f579cb4acb436ec2aab924b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc27746c5f2b4c3847a4ca01d13e1214f6611b3b67dc2749fcc19a4dfb0ca540eaa157d72d38d8d02bb56cd2d94ee041b9dbb9e3cebc234512df5f82299fb129cc2bf426dce8680fbf5b7ad67b6fd7a707598c9636ea1f641bae0e4e86a88622510ed1c67aa655c4311d561f547d18644b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84e88381e119b0465858d9e22a240c870f9561ddcf64db5074b5c8be57fe27514fccb00759640d5e25c1a2db6080c746c2cc3772bc1a45a71836f0200d7f488d7a35f9f6a53ab8e08f0421349428a59930210a18271ea354c3deb596e3597461c1f2c42523bdfa818397d65e8dde27c99;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dccdd152bc72add7a674794744de251ddf5f32e78df2b606df78d2ae6e264506ff719bc1f20e8ae9b887125bc8fd7ebd80b044eb74355966b845fa132d0858bc4abb181d29aa1628f53ea2c22ec5e45cce607d71bdba1cf623ddc7f2dfcb565b17f9ee7c6013e4b1fa6970bb09b26440;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb080b82bd9558165281811c64d3968957cd0ad3025a7837b78ef36fc0a35760635d2f7c3c2f8b67cf74343f3463d656ab12f3d5be2b5cd2908e81ff187d14d01c8813675346026fc59630b8fdab4c8ef645ab371c3f67616bb55f388ebd77ae0710e3f2985a3f4854f1f2d8bf27951220;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ef35462867bb7c28d443b5c483aeef814a34f2abfde903f83a1693f559407d1e9e3a50ec6dcee02330983198fb1fbed467141a3af5d296c1c4d4c38b4b4a2f618368df635c49d015331fe15995a7554595028f517e9a1987c106440f832e91f569078a8247d3e9fa6e63cd5a7da4eb21;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haaa1956afa166eeb00c62e1da410117af3820ca8c5eabc0d151c835c9352138daa0eee5f8b88dd8ee59052f9554c270ad7df32d96b543bbb1383bff46b3317a4c4e14c2314ff823ca0c79a3a9a774eb64bab6eb9a0a5137c1c4374bf0bbaa1fd0485cd2a5f88d2d585ab913fa6971030b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4cb94ec971c3acf7399012fcf9441c058555864853a9e693502a90d618dd9862799d296f76f8f071c67bc44b5c8beacc51a04ca60b6da5bb47a60513f0c917d24ecc216d7b83cec98bd61756a1dd5ec79578f84674721d126a9b84c6c85fd8261d5ed80e96ea501d5e1967f70d9beb3fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee24bd701ba0b3d820b9d57c9e6825b4f528bf76ded8273e30009fdbc8e005aabb573e15fc540863f68fe26caf4addf2c7b90279760e29a0e3d3740a7d72cd48006c28da26d2a857963dcd83aba620f60403c6e034538e7e4c44913974810f1651d19fe3c12e35d820f370dcd5dc56c64;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a365771af55474f99e97418d366c7179c3ed03b5fc06f8a093ec3b057ae160c84efa82871081210be1fe4d5199705bf41541c4b683bb21f66f9208ab9c779cb7fa8313a5988ffa0639515aceed758b09bb617f968cebbd46386b3c89cc85012cf1811ce21874e9ec9a2c6607e582dd1e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55c94bb91b04cb9a6674cc74337fea3a0a253285343cf2ed8f4a5a83686775e70b1f2ac77f75c0f72ff38b41dd4e40ebd0942183601a687386f22d070d9ae197a6ad6560ee55bc16787bef3b85de8325dbf1886f57869961041fd48f0c39912067e25d0707af69cd018a97209b5405e5e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he393d22bbca2f695c9840a217d5db845f75068d87e9e1e25ba5679a7a3d35d02d3093e84034d9238857a3ce0c17b7b2c8a8a6aa0b73f48c38518eb47d7991384633a46e57f9383191e6dfcec2dcb839443ac54be6df490eb59b87355dea85acdee648e51dfeeec5954b9a178dbe118c78;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d6b05fa6d2189d695d9d65efac19519136ce33704ac32b36c96322475b5209cbf946976ac05f66c1c5a46c49257059bdc66b016dfd65f62011d4ee849720d97868ccaddaa9d86f9688089b6a7ce54e06845af3aefc68c83cef66c250509ba110f9d7f5a1acb53eb467d2117698ebd90e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c5e1ae656c668f619b1c1133874fa72cf92c4d46f5a62a729c357fa2d9ad09581093038560a8f29893a485c430550c159820a0639bb1ca65680e2854138e85dff3c60e54d0a9ff0e643a6401d7e22604f277b97041f909650ccb101a6e361e48084f9a786d20d2fcc5b4e35e34b51de7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd204a41a69fbac05f1a8ec6b4ba469a01d984353b8e52c3b894e88d23cba793b3aa4f37d4a913fbe0dee7d58b5a49e2504de24c36ebaa1b3c8bf54cca24bdb9fe4667715afb69e6b8286ef8041be5f1a1c081c10ff167367f69e1ca9f697d4d82a2b9e5d0cab9b4194b17a98a5cd3e78;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7428618cb82bf0b95c44f7624f674034eba97cf62cb8671254f50e243777df8d5579fd4623cce4db38a5462def1ea1721069e830a339670bd4aa7660c4fd6338eb30fb3262202ea885c90d7b302a9205188cd117e6b27c4a78f031dc30f12adfb3417966a783c81ea77af34160a70aecb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2eade3fcc2d172839c09ac87b8458a13fa6f0372d59fd8ae8634dcc92229ba22dd610e5e68b2839359ea2de86627613d87cbba5bd8a57219ecc8aa342c25639b676d9e6d1c264dd31e4a887998cade5b038094ed2a1db63d40fb9f9cc2512b160f14ac10eccb662c062b3751ce56de1d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h293583f67ebe2a105484e975989f326e0e20752bda1f09515bb2e42062952a8c2ee897a81e8d6396113a3b656ea46e05a0faaef30b1d4f95a8ecb7b85c330cc38c3b186f50bc820a2a0eadeb3e21f4ba0a486b2acd76e38362d2de62111888d0d9dd2c3aff4e5541336959db5d8612196;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41f88f7560f65fbd1a783d80d0a6495e46e0653a6b7f873d4b10385bdd0a4d5c6781836e9c74a2c402aa0028087d4cbb90c420b09871a85c7c9112c6b75fcd92a4ee204499ebcc38d5075c6cffd951653876798c62159f5f81d08cbbaddb023d754626c392eec1bc56a7a61953561246;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91491e3e5620e26c5e67e887641e2feeb2c1bc865ccab88f803e6080d43a44d9c817c67a4d3bc0bba071418571881b326514c999e0cc8342995ce78cb56595fb15bfbd43b8b2c7b4f3eef2407421e20c08ffadb155e9a7f9e7d26a6b44164bd629b74c23188d961dcfa7b70b6d52faf10;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4716756d6906a625f5980f70f1643c7c03bc811a8fde9fdca17620c0caf37da2716b42026241637f3f8cab9ce8f1766ef6f727be1e34587d2800d3a30bfc0cfaa05acaee053457f97ea92d154ca7386aac30264b6e632755905f073c76de5e77e5af6f52e6746ac51f20de5b38493b66;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3ab8b6692c4cbcdb4faf7b5db972b437ed2af86181e3118013089c7267c438fcba147d1898ac17c0bc5185bee339c81c5fc4354aa97f8bd824073a6db5723e3cd1111dfc0baf63ac4bf50ba34026773190467ee3f9c9b78f98795e17c5c537346baaf3eda9fc22454d03dd2ee56860ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9fa0e359b6fa436e67a6f9f4ad3a08f9617279b88ae01b5b5a7567348a4449a0dcbd165ecb36f547450e365e598ff1ecb209e3564beec4e0df91e8d0db5b1852dfe931b4d1dfd499d95a0aa0a0bf390995c7de8f4b04eb8d7130eb9b01fec89a89a75f709a86e73c2673f3aee95cac9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6b13a2e9b7a5f1b826cdc8af52c958d5035cb2579785c7a326b5c249ea4843e482c8f5aed599f204af1a09a8f003824959b5d1891f0026303edf216f324a34bfa0dab73d448b2bb66a5159ca3067f8317ae23ba27bb33dad202b529d11821483f79f5a52921213ccbfb1ab1513d64c06;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h429a0abc891ae89105150b7c1619a0cab9800da869dcc2599e1494ae8e49adcbc6fe04162f77babfef07078c97b6e5e32fe044013873779ce8a7dbe6735f647f42ed7afe941d6b98ef32099a96e866b4828b19fa6e9128483bc831f39eaf8b6cb4349cfed7f6b2e2a75b287297094c56a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ba5136b57e3a9ea29dbfc57a8ebb199ac73b53eee5c99808d55f3026a28a97e64ca360301f4809e9ac10e458bb4109b06a3cd3a6dd458f54f8c900d51a4902efe443bca8b85bdae4fe2a899070e91b08684fcbc3ac8e768183d8233eb80e450b10a236df346ea32c1a3a2e01e0c6d405;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'habc1c17c522a23fdee076a0a635b3e2a9faa49fdfe222ea01224a1acad6f9349b6031460ca1f02660e68e035a611b919222ee023a5e6c1ec0574f76b92725ab119e7f086b2b2dbe098eed9487356bc4243e5d074300c4ec5d23c2cbe0b48543617932352b69058a8630cf8573c524d294;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h429c657c4d83f056870d2cfea6c810b9be61e50fd90673dc55bdc0f820d77a34b6446b4fac7252d28f00ede3f7798cb309c63de33581e61393f3af9ac7fce2b9f4d6aee243363eb7498d5529870490f7a8b7b09905e3db76ab4273dfe10fd1673c03f43b09b871ee81167612f8fbb54d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he05f3ba041e59b430cd9ba72697dd15bc638f9bbeea1fcaf89421e498832305ffa6d20e365cfa55efcd458c6099dee1d25e541e9df42ad907bdbb9b1095fc0ee761ddc678758b5b3f597d405a720b9f3870d10eba6d8579edef7889ce4c5f32b4cdef591fda54865c868a6c588232b7a7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9773605a9bd87423a05e8d979726401037b0c50473313c0d472c477374d4c565f2cba462a468024b6a65c49c40d7946f827471c169afcd0942c4d3d324713c0be618ab0e8d4378e045679e11c2c549e91c483b25d8cac5715ccb8ada88cfe6377f8bd33bd1d412f04263586f0717a7419;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h120a84358462a58787e21c117e784a7d773e994a3d65c68bb052af3defe7bf476bdec3025e30c995586afd66cd6ff480a30e95d3f13fdb27eef606dbc557df0798a492f0e0b6a9e08a24ff6dc42cfda212a1638d8946f0d347dd85856abc8844d7daabfb0a882c9755fcf8c9ebe18435;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86075f18870e59d9cb689e2da4e2b719c31ff1322a036edebf6b84d922a4797f3d80f714ff69e5883b5b2e3cb9286502d64d35799b8c31514c17b1cab2d85ce200fcc50d8d849226536d22892cad079566e24dbb394e1b633f5ac220a8a7a2406a0b0f1bde1f0d3f34b1cbda4f9f39824;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33a33779a251ca6941528b15b5f86013073145aff2172e8e5139e239b162420e92d3d3fde35e04e5786042dc4c44fefe78c1d8f3f0c6d38c195b3390c1dbf449d4e90d718e9944992ca6e002c06401c9aa0336b269e1808991e8272f973b08e88115f0cb70ee234ef38e65a0828c19aca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bc02afe46d680dd7146ed010423292ede4ae8f3ef5220046468961b34696e8b1b1741a91a3fde3a5aa98e025be703eb53aa69426762fb98bdb157942f707d06a714e64c1771bb001e6086856911d0cdda5c12298ec81c2609fae7dea18d4223a2c7fd9ce09f72115078d636156203497;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb7e395c9873c7e0e4e36e40dd66b2f923384d4919361700131b311e4bfc4fdba6376f642db24b0e6eb7a312a80ea13dac06328cfd86690e981e23a04d28fff104374f1a6da1b07bc3b09c761a35745245246e7fe7759a3ddf8be7dea5d8d0e3a97a603e256905c7f118e363d11052eac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c99feb7f82f2a20a33bed1edffc9e256a30311fcc536b669753448425b74d205509cc2adfb8f6c48d3a3444cca33b59059972813044f4f06af9eb385341db8d219c2a641a1cf809458ad32bff3953da956c4f31c87df8693b5604ae42e9490ae013db20e9333d0332a5434e2a8ecf078;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7256db063c1c13b41eaa5c5786ec4ad41ea5f04dd04cd3963e4182b511c3d44e65f2663562fd0eb434c4f88152dc5840f382e3765ef936b8732873b609ee91aa963b2733ee225368b57ae3427e370db27a06c72cf03cc3ebadc6a5793468fa523c13e9aac1815943f05894e4e2dca8236;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfdf539d0e54a4fd3e52501c47f3b139e1248f728e1854cf40d624396089cb1d90193761ad34acf0e8a25bdc377f473d7309a326897f248fae6230559b831f9f79083a7f14893e6de1cc864d56fe7eaa7a9292b8915af7bb6e5238db12ed17e3ef69bdaf19b88409fc01de8d8575900ed1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed99fd8ca76ee0ef694927815ec7925a91e1af6a94e71d3b5c89af9d65271cfbbd244d28143d324a77e389344f855c0caf4e18cf8e9ba2a512244d64db8a0fcfb3260101a842597a37c29c318dc07ead9297783a7a627469f94fb0ad296906a0d20a7700556f4ca40ce8c94c2007eecc3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0c7e0816bc684cf08c3c2275f8aebef2f1d58a322fc6899ad8498cfeac9957c1d4052ec9aeeb60a547b9592e86200b2882f3c8e77902e0cdb0a55a32b8c918640c69d82aed73487a2f8ff9202522aabde974b2acf19c0c028ba31c664b3287063f280acd8e04923b2288a3de453146fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f72713bb672b005f8365d7ccb22e283c4e0629317a89951e146678eaa9738483fff17cc0bce2cf155beb2e702644e0d2077150fefa27a3326519291a41895bf6af7fd26c79a9daf4abf525d95adb77cad6d218f4a9b8b4f648c6b9ed8e38c49b8fd342877c697b7c90cbad6bd88ca07d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb91e9a52d5085ae66b502ed67231b5b49dd99ebaf01a1b88b732a96c28a98ac7e4f8840431e54d56a40c73a92668790de3c609cd6f0b0a57d4be111c94993baf94071e06f90eebeb55eef262e3f94017fe23edd310490b283a2c3f2c99ea140169d08316422eb9f78f52254627eac046;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9aa9a07ba4c3b47cdbcec453bf312b40776ac3f10f883dff9bb2c420a432b92b8f82c171b5404de0113469f59fa9e70ad4e7497ce2cfd878ee800696a228aee395d34bd8fb633458e674aa03f2865c25251101c09c8a45b26e6aafba0ff778fd6ce9aaa96cb3b77c831e988198558f6cd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b86528c5de7365791ccbbb76c58a562d0945acc0d2c8bfc4b1fef24b88d79e2dbce3ef42aa14270a3979d503bdf315063ee67d2e8f49f95056c2c98c120fce895f7f6b3eb341cb896bfee1625a225cef990707b352a163a6b7db60b0462ce81034ef7448340dfdbf457adf79bd1be55e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha89f8b8660332cc3413a7821ac90c6203ba3dd14fbbe37a7b97006453966100bf1ddd5940bcec50d30dc3da08030c7377392717d04e525f9f56b6ad62763e87fad2261ab8fd41ab79b92cfc20f0a308c3d3be02a24c3233742a7c55c997e390d2cc4f289530cc2de5a1c7ff5871611061;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h278a0c19a8824085a503501bfe08e42be52de8a646bb7ad8a962df00d22cd9fe9b4597fcfe52038d55970a10ea45e4d85052ed5182da1a72b33a0dee096c56cbb4c14ef71c9de7da4b38db1eb1d6ca1eea5990125f56f42078371da58ebff525ce68415fa002496d2cafc96daca241aef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7f35ea1aca0534288d5a37f401d4f70baad72ada389624725492085cd4bf329e163fcb586cf4cf913387b4d2436ddf1b1e770aa7a6efd2030af343698e083e65c04a670f450e2c12239c911e4126ab02154cc38a9528f8f0a7a2e4a192e7d63f392aaca73171997da2f7d38ba5c11243;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44915e1ea899a42b125caae3688ed23bd3b1b78aeb3834aa30b593f59282cc67e64d0f00a4ab5cf9dcbe5f6ae63199deb1c8afbc9ee0db799e9a0d6f8d4d0951b7154676dec86250d7c7cf57d3b788826060471584d87d1edd85e07097b9a03d66f9e852b27edf92d3b64ec5f46c2f39f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe8e4caab4ad5137db1852425e30c1a882a196ce483a9f41bd0b855db1bf241e3783a7ca00c99dcddcc30881a18014397c6f643ca2e1091d6970ca8ca1a59ee81a6d6fa63f06c5e98c30ba78d1fa6a8408e46355add2bb1a9fe034c9d29445a36cfba56fbe9ab2a7eff6562de30f30873;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59529a85d421a7bbff643b625e0b15ca38e06d9fe8aa6824f28539faccaf341ce3af59b218dfe911f2caf086d7b97918da756cf23d867b358bc44dd9451e9a83e78b54d4cba92ba27814ecb316cb04168c1f9dedf15d5dcd94819ca9802992625b56caafe52e51b414f2635c44d8b6761;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e42175fc3d5d9079b8f64354d43ed0bf908977d9117d12073a26e749763c0bad363ce2787fada210f1406f427be51b667109553a07ff71797c00ff4abe37a7c57efca590c3218a807162febfeb18962b87381e856e67ee7bb61da50ba5a74e828e217ec044f304861d48dfa2c73334c5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa63660f05588da0e822f27fe0151ecfaab5d092e361826ce73b2ff79a62babf354d28598e41af9d273a964c74f7512486ee0ce0b23be27e933d37b240c9750f02af2c5e2d9901aad0a4d4f926a0ec48ed7a26dd139eb2c619fd4fc6ac0e9df814d8e85bdd9d1048fde770910ef0642f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6642f920dc923aa0268fbad4a7f913ceeba9d34ffcfd0afca7a6b79b7c370b3fcdbc9934dc4885db3ad5f9823c5356935ed5a945074c966f9e22b760cb841be0df43cf14ceedad070d111c60c9af22b0f050742906fac4ac7fff26ad6f35a1f9fdf51c692a2acfc19853621a0186ff1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b135b04dad04b0d22df0c7edfb7c8499b62c00da1e57304938038a0da83215a5054a9ce2fd6c96758c51a42b7195093a7ff03201f220023e312483fb0158985805877d72705cb5fdf3f19ea03bd0934ad148ae4f2d4ed970bc9594f2230c9cdf45c52b2e6c74b69be44962fe2c8342c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72b536de446f9437de394da7fbee7cf10f2fa7e22a2e1b984b07dc77e0ce84823135ac6ac263792252c641beed022d1263ba65f7bb8aecb03fae0dcc1cc8089efe42a1bd2767b21e6c796ccde6688651fd41f6734c51cacce53c21eac4e47cd3aabbdf3117d6ac27da6235de9c79f9ecb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac186aa804cd6b7e144403449a6a66aba803d887cdaf9f552004baaeae40423dd611ad413e0c67859af4d05401462d7f615b5b172a0770b4b43b74d1e9520d344a7ff98400409dd6e64565a9eafe96ba32523ac8371528cc447045762a516436ec389ba2dfcf5a6d412c5cd3e70d4b3c5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57c57c79249e4f2470571b94f798b62cd00d9557839fb163281cf5e9c3b41f945529a7c499426f044c8b5dd77b0c60abb481309deffd2a5594541c313b2a39374e30056fa7bfb6dbd64a60f77755246da9214bea11a7aa3b32b80f9003ec1d56904f33ed7c32292226437c62da93fea0e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2702ac776626ae4c5afb3342b6a84a82a507efe4cf4863ee7f8275d87615e36d9ab56c3919debff77f365ea272133b76836a200ce0b2479e670013a2679e87631052f3510f66602d4378d2cbcdaacdade2be980b0a386c364e389498ba415404061a360e8fbc51cf1b78e8d1b504d81e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha453637af8553242dadd9ee07279b0761feb70c868702837a999c9de14fc58ce455ae7736077e3012d25b33bcaee0980be450539a6f0883057a98452aba39a1f99cdf9dc5fb457d0b1bdc524a82ca5aed78681ce259d913cd81deb7705343edf0031c11907b3981f73104c28e90379f3b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c4abfe296954d94ec8746c8dd2ac596b2a67e8dae94138f7b5d9b403ddd3cc8e66a080f4cdac5a747adfad5700affafb8f419d442adc10d5123b64b56420ddb67a6e302e12c8c9085272bf98d25efeddbf693c3be419fcf6f4cf2912e2e3c1a0ce00d83a666b32841f19b19f129a4b37;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdaa92d827e8e1b3979b13d4263ee877b7d61c06822467164c617666cfc026b85363645fb50b73f667686f88acae7fcec5338ad821bdca754de07b133be67421bc13264a420b2cbc94da773530749be7cd48133a48a40bc9fba0667daaedb735ab42b83b929e4480b8d8789c612d80387;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81ccd137eacbf8cdd68211c689c6c6fea0e33fbc47ff6f39424a19341305e43ba25460766fc369bd72f3b93d84d29ae26de68a8e4ba6ae58a2845f93d90878e8af1c19c7b527b8d5e109101b6bb5df5aa1aafe951ae9124bb1fedf72acb0d4242d442b41e814ad6de40df57551a30fe31;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e45b12e97a49aacd6b5a5e481675a9bfdf64b979cb27db017dfc3095d6a1397cfcefe43fd4a5e5cc60650db69738f488b3212bb6161322df519014a1e9f5d3f5df748c1bf000175ab8c54583f699e6b82d770c4903a8928df6081bdc154f8856bd212d6621850143b5b1274f028f98c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e5c68cdac88e5eb36ee22c600c257af9e3c05df7bd98c5f385b398c95d3fd7ddb62baa7fbce2aa04a2e971a546aeea4a20e5a7806185e8e8de477a25b67431fe36b3625f65b611eb06d5d5d14598280291a745f0fff8b3032969cb5d867082b0051f660f4f3dbf68f3d9136b5e01cb39;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e1f09e02d4ebb9b045721668b890f4e6629cf9e844599e5219df80c8c18c7f05471ca5d6b428efefa35e50cc956fe606c03bc18c50dda2f0e605463c7124d3b38b74806056292c42a0a8a4d432d78e4966a524fc03b10cbdb8577975f569f59421c0120af341faa619a0a37078a6ce72;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6133e19d0f8909608d8cd487df6811f4913386351d055786faea72384b63a713906005de8f9351ae365ed0cd05ea8dfc3fa66eaf7d332a06d9cffafcc566d9dbb364043ab01848922b2ae9df79f83b4eef55ed5b928546cf4c7f0b130c5bea4876b0051036810060ceb6e90deeca19d17;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcaf5f6abda1e48a24644c815555bd8aa96980b16a6e613a12723f74abf932df06da7de4d24cee4b783aa43d28136434e365cb36694495c45f87aae4a5d7644f7a82445995fde6af226c2c3c0d2e588bf6048f2c3c49078fd22f5a50a1ee82657f8e3082d54b4adbeb6e41873cd8c5cac6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha726dd6512b27ecbe802b07f2ab98ac9e43935ab37df14301c3374c7958aa172bfad84eb965cda710fd6e8faea639e033e123c553b4c6c0bbba1dc1a7d1e3ef3777a055dacbc03ded28d7a3899660b58792514bb83d4f27b019264deaac9dbb3f55adf54de6ecbae6b8e39a5ca2be3ab2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10900c1dbda8f5a3bcee17874619b015c30aa70fdfaaa446bd4ce7ff4e4355859f63c6c3b41d32a87e3d4d694e4de16001959f1d2146a7ddd2d761b5d93977bbaf15a2dd75460f805468a058a4189138e34eb84610b1bc52d23b9821453d4bce5cc27fada086e3a7782a5be3d1fed63c5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4374d25f1e8015ec528e73ccea177dc83c60c8e4f3722a1fc47ec264e12904c7df787879ab7f6dc02192b21339319f9f377398f9f6df6bfb09c6d100c00a2b403cb3b784eed342ec98a2ea7be99860abf1cbd44a311f3a14755c23b12f1fd09d70cfee6fbb3f90acbe8789af74068944;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc627ef052c288630d59d190c25d7834bd39a8dfb7b69f7b020f8de599acbf43ebcce2a63ae7224d79bcc5d4bc614d40c7856e82695ba9c6fcd1657334ed3ce4ab8b4f1ea0a097c2a07cb3d0c5020d8c34db020df4c022ca33276cc20320ecefdd8a2d50478a016fc2605daea7c089a034;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5cea39fa4657829eee735579ce5dd34e017410bdcbc73a061c5b65c677534d8facded8c62ef2dc99cd8a6be1a1a1b2074ab8205990340d4882ce9ff1888af8203f31506fc76ba38a29b3431ce6793555c767fa76afc138482737838c11584402f1fe17282a96d8a6ba80405c1aa0eb9cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9febc0634547505dfc3c75e56472aa8fe85f6c96ae21187428ab85ae669b8b2a5a6dea618d53aeb4c9102f8a5ec0f90d341fef9ee915011a438958d53b5a3786f7bca4bf5a7414564006240e7864208fdd551f136eb30de39fdf4bcf63e69e42093d994be5a0e831af533a858f0eaa4ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49beee198db7d916985b7232c2fcf591dc8915ef030309f07031e04631dc60ec0dd1675cfce89b52c6e691a2f58e91ea86dfccac950d580c8065b9b0a29fa8ed484086ffd65e44218e0d93f7d7071d028573c8a5324055e15c63b6f95cd44b8fe95eec10e332e89d46f384382446a64c2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6b36769233fea205206d80dbe6a98c7f8b7d862d849f088825febe93d3c81b6005e9a6f996ce91a81e1424988adabd3c3819b992d01e0bf8bc7010670bbefa307437f223f8a56af3b94ac3a48fc1762d1d046c6172ddeb9db3ead9751c3630d45f62ac659f17f8b63050e6e329a1ce34;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc3f76b67e5344064adb3e2d85542003fe64b8d55dc26258756c27271ed325204a10e5a8349255ed1acc2d9924a9327c013324f313ea2694ba93307ee58712acd4da459b557abd9347b950e0b4cc4071fc0704abb4a8a6e0af15bc7535923471b174e53b352ae33993b78041cda1066c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5fd266703e9b28fc595a4240546bb9395f9f4a838109114a8de33b5e2e37e6a27b81df94b9cc7b3269a3880d31f6e6542a95aa9855f78c8cee7663ba2167fbd5add09c13469ded730a74ff405f360a36a68fe719204f5499ac8e2d390ce4e82cdcc1078d5c6ee515d8440b61c1b7847c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c1f04bb9a8c2eacac8ddee3ed5fef136ce6be6a7e0954e00f920224501e672f8dac8da20158fe1acea7c4d71457e73a8787f9d1dde322f9a5c53040af429cf04f07212cade0446c9644a20cd133db98696195f606290c12223f171ab0bb80bc752c7322741d5faa1c51e3138b9244f01;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f6ac3a01bf55a3218640fbfd367d0a096c2a0fe2ea60941c3db1a84f58cf67683af62d99f97fa2e06b33fba45bea349d73a9a7114b3568dd5ba662b195453395caa95e420bb0360703c453aaecea03d1ff249d947cbe76dff790bd1fe8a9b4eab3799c039664caca32c99fd2b5eff14d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74caf9270b36a6229ab1fc0cda8760438461c18ff7a2dea65a0467ccf54dd7ced5734bdf6d4ae5a8e41ea12cc451c66a5436b28feb8d0e7d62edd302155a9614a5204a146639f2cd85e0a0b9f39af4cb66f5b3222664365aa067141aa1a4e822ff2adeac3b69fc4a12bd876f6afd50529;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f03fa77b03f63061bc919ac816b8d696397cd3d479317dbee02adc7f64124fc203dc26ba16541511389f37ebc2c041912ddd8d8809e124b53dcd6f859a13dbea927d11a41c8c26e71f1c55d30e20fa14527a0d99497d6e8b163099336f9085573e971620b77eaf81069106787e0ef8e5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52f2525d9a2f82537072385046301220f24a825831300d2841e4957c53d190e61ccecd07dc268f846b5cd722c560fd56970ab183583e65d09796f6535cfd09ea31283635c5bb5a439fcb5e153bc8b3b4a006e808cdca8de365c4f2cb4869abdcf9b3d5fa40f04b8e34ca682b8542edb28;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2562c73c0e3c1612be5d2da85f7b358abe1ee09caddf1cdf28dd3a13958bd6531db1c73958ebc4a86c64af926a31b299bdadbfdab3e9b7f9b2db7813f197a677ff6495219eb06108cbbf833c3f8a5e6a830b7b511ec89e1c1cb6e21031d579d8d5987bd7ab40c9243feb3c9d6a62702;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h264ca6ba1a3ef0b7fcfebe3185c823884051d17d6918bce9773e5daee8b962ac14f7b081e95a15e2fb8143ed16927f6f560616d16b3f9974b32ac949475a63939da721a757a76c7a7895fe558c99430655cbd3f20a4421a18f54f767a3729cbe582c3c1128ac410b6bac29432a74102e5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12c6ea4aacbe10c403de663fb74afb1e96a8fb7504cedb8877d65f973029e8cf176cdddd878ab58febf1bcbb65523d2ef9da226091cd9582384b6ecffa085ff6f173e40a460dff486193113ffb5d520d1346a4599c6f1218dfa44ecef7279485427ffc6d2c0ab5bf87e15902f11a29a65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b456aa2fa212198ee55bb8a973340101cab9e43f7c8b5288feb53ba21376a765fd21a5fb53bec0440799846d66b1a2c00c4bb57c34c5125ec3b557185ecb2d91e276f708c96e958d88b88b497b2790c61b20f3f862130f49a281af640d3f17139fbba0bfcdf28bfc5255924d8abed593;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2877f1e2a644b538fec224f0116fd30883514a7955d665258a01df44b6533e1583258b1aa27352e52c32669a0d2408807d92267e42ccb8a75aef32fbc54c3528b9fa7d2328ecb16a89f4f652c84767c959c30948f08ced90d6cd7b6a17d064ef9c9e8463c4e06587eb6dd6a636193d815;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h825ed0ebe3fc50df35839949e30604c8921c179d040a5043e3b905c5fc16d93360849364ce033973c87d688d9f3d467d9d81cf899089244a16880aa31f67285a040cd823b993845b8e2377edd386e4dea7818aaae2d9a14736049822d7a6d1de25ccbbd08d5e9a8e68cb63eb534518004;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h276c37400a555851f68990c9a64f3a47d31a8963e71715d2f0e08fddd3b90cd6c24f8631fbbf5f3309c44c5d2d73b91062daff17555b7a72f876fe2ea02e821674c44a96b9b033af43d085e04af8b1d884827ef421d44c8e828e2b60d7334b25cea67d7e7e34da7e64b2fc48682a4bde3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe2ca802262894a1bd25036be7764677744a4686b71b4f4cefc7bf4227dde9846a6a3779cc995615ee634b4020b6ad5a027aa760a9d251b6e5e25bde62a8114d96f1dc4d8082fb590ff1fe5835fc9f196319db42ddb269c05bd9468e1d35da6650902b7a5d46df0a9f24e7797378bd05b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf30af56410b9df37a93abed4a752bdf8e353afc6d34497847fd34b08e67872c2642c0fb1b0b59350c0c2ea187ef7602412e41c91c0301c7eec1ad42d313fccc5fdd2033e82841c0da55f194b9b994b7fac89336646314a3bd66297806de2bbe8d780298238afa3010bc1807e1566142e9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4935ad21da0d8f9253c39f997280e12ac4e8ed3915dd4670b87243589a09f60b803332b5babb9266a220e513b33c573487d7aff716e065b936c6b7a3eac70a8fb15709a2d9945fc8321805139f5f073b8432827a9848284b57e9416b59fe40e62d7f0a84d6e27ca196635400c92d40d92;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h999fc3879fb4edeed2d8dd45a39c314fdb7be7bb4160b51253523f35c8f0e09cb4b50a28034230cd2e5890f406fe55f9693dd611986af21d0760367e344e56e369879cb1b0811ac122226da7986b22a03e58d6cc6ec19ecf7c3cb3d34b94b2e539caa45c5d15fcace94ea1a4781cd191c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64c1cae46e94d373db0d77fd1010c3d1a750feccc1ee35480fd1eea867393ae2789bc8a3c6a4c065b0750912ff5fdba02745b6696446b0709e73dafe4aea391eaf22f95a4569d32811c74a374cb11c0e0dacc0b9e2c7f136f21678e307ea50a4803c3727218b43aab49b7ca7c16207d65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb244d3d10597a3e50e1048df4c24c2ea30f412ef1f59d113ee49931b45298d91b97fc493a8e1a2fd9c5e8f9a3b64bc0128fb9550aa86a3a67e64f0db56953d3bb8cf6d8937b6a5b57e65613140fb054409a4c6c63a9d8efcad5bbbf610e8f01bbf9bb82fc074250fbbb0575e624d971b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ff6db00304146ab22ffddd42fc25ec361475a4adabafd00cde463e35640860348ce17d120dec677ff944d625d0fbcbe6ed9ea43f03f856fbb05bffb475c512929af5e48ea0a665b5f7f9005512d4fa707e324d12098975ccbd4e24cd1d48ddb4c30f2e7fc5634dbfde4af82aa9a4e2ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbeffd66dcddc055718a584279737abe7ebaa4f860ffdae8afb08ba39e58f2cb45ffcce3fcecb2dc7840c53f1099aaa1123e9086475ee7ccad02f9524e64042eca3c5a5e1d34d19b6117ff2595ef40a10563beecb459dcc45e60e67a19dbc1d9857abb2f420e1e7ff626cb22d854635f0f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77d875c83d4598e0fdd433eecc427036d8387e9fe085924d5867c4f23a4fc10a61da36f23a02074006080476c89edd8ccc0983a607ba3d0dea04c36c78299d43e0d77e73c40d39ad7708ceb037e9704ae0fde3e382bdbcd9cd9a8b43f832de1a52b4dd773fd943e344c769f6770648540;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf117691162bed50199556c97d85ebd4aa238ecb071409ac7ac4ee2baeb2f475859e37c19407e81f63303cfef27859a97cbd7d1db311402b58e8bba39937a3e340a0f81f925fb069128766dca08144d9e1ca947007652e8492100e082c2d0cfcbba86d93f95bffe8c26ffebc5808fb3084;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9d87c9ff34ccab3bcca0d1bdced2648a1cc5fbb9d57112b98b3f9ded441b79f4123639a9c172e73c3517e8ba40e04dc009d4b8433068c865c6bfcfc3dc11632972f519dfb645d4131beb87129de980744b7cec257a70de0f6f7553c3c4f8c006e08809cfdc30e4bb1900ac1164084da3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h407a401f334c8c33f142f8d5686775d994bd06df0903b8322aad6bc4fdd34c0e275e3bbcb986e1d4461ed141799a80a4b792ce5b1d677a620a96beef45bb9361f4cd343d3a2a2d884ec59d038c8364d56317c18a90838c4aaad9e8463e64bcd0fe8270ad83b6678e65e7f5c16e08fce76;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e6c301f4ca149adc5127a7a6487721b3ddc436e3f55f7517e4008083a23cb13c18a9b80e42a00485c55d00159bdfd61a99f14e56aad0b401ce8b40c36d7cbe63b73a57fbc8d28b198e04dcb3ee57e4a3bc18d62164191e3f302625bba0fa30f2adaa8bbb818670f8a265cbcf946c1b8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4bc7f9a7a84187ea09c03061fd77afea7c3327bff793a48f9a089e28b10787ea03c09d34c6b9c10789a7adcd71095bdf6bf8acb8df0166f6a1efae5ff27016e823bc2094d8ee2a5e7e0b2bfdd66875e5b6e75881ebdfb16ac0eb230cdf617e9c18b20b3a72a991ada0a4c9b9aa47eda2a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f3672b294b53d524b4fcabeb066d62abceaeb1153ea9e2407247d10ee305fbf01eefb0d5de91997c733ca08ee0de1c55f6ad0500fa9d710e4ca3c28bb323e7d74d0d918c2c1e61c397f88b6dd0e973510a63666061e227badd4407721f4be6d31b624afb7907614f7ebb61c31265440e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd34fa389741ec0bc75d88bc719631e57773158f3a948f21cafd7d085cf02745d4f6bb39bffd19cddd210ec14b3255f212350cee1732a7cba11f93b93c1c3106d362dca402b1ff02ca85427df61bf71f892dd59bc29a4019a329266323bba33d7a1c3f73c16fde52b2d2ffa14fb43be3c1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43561c8a8d5e542f928ce34b836aa1217584cf29221ec9ab8343dc44fc2974edaba93597435e2654310deadbd1dbf5101ece62bc71d4748a4d5a6ded22a7628c7b93fcfe2333b981a9bfdc11ad9c93e37bd3d959f19e8d691749a63beca1e573b6ab3e3309cf7f4834768095f6ebbfb64;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46bae64a7da462de80b5f51ae0bd52c713df9d90ec089fb684d3c26cdb5a3c76923f1fd73711412fddf3a066aa8340f0ddab8b614c31d0781f740ae32495863c0803589443088cd9f0e33ed29ba0251fbf6b20b97a87ab58b1f01e4569591dbf418a75c300b91facfef7aa8b04dbfa3b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a7aa27a19ac201cf903fc5b7a4089b277c65a9aaf55a3d378958894edf48c6bcbb7e1eb514513320e91fd9bcaef2e5eb623ea9aa3312cec9075c25c7dd68fa501990c26238890c5d27e61e8bdef0cc6d2fbc90474100f4f4237d97cfae6cb6a99d087642bc4e242ae319475816f33925;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d469bad21b2768ba99f7e04c40ddabb400c35352e4ac0029142188c51eace5123f3880c5c82605ac03ec8a07c17921c7ba1da5ee97c5f26ee1eb4a4aa979219fdd3752f5dba1c846b3649577f199623fdfed1b98e4ed98788aec839a2513e5e4bbd05a836ab148a9d9a1ff81c38e7303;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0bf21f269fe29b5da2ef9a3c0ec317b75a82314ebd39e272e712e886aec25021cbe555601350d262fd6b7ec244b196fb9d9fbd7d07b01bf70ef2c64fe2cd82bdbec2d812c8950e0c16ffc9c86dca759539fabb6a5b4430e60eb75043d96f361b307b01b271e0f22be4ac022df4f84e17;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c4585a102f9ea9500e4de86ccd9b9eaa3523b92a889fbf3e1102cd9e5ce5ab11053866530f764eb50782e6641359783153b74919bb8777e8499b6b076220a8e7d271a3394c273aee0d68510ab48122fa4db50e4c11d692457013f35f57ed7e3d3fc90673ae81555416dc9ad360afbcb9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had4d52555db9edeff25caed3b4e7f59e9b0d00e0b757aa8900bde1109faeac15e72c078550745c5667f55a6a76caa0d1ee005d660b41d7d8762b8d28bd7f17ae4dbfe90b29d977f3d063776fd77ba56649560a036c3665b17bf832e2163a34675f9a14090d91bfb4b9be4f383421b7d61;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d7043315026f2089a38fd0c8683e1f5ac01cc4426f62b0c1e38e0472c1542a03d6b71b69eb7f690e6a1aa613d4283e74d3ad09f4070111f0f8b89b7b4491512d8f95abe1f975af7ec89e3c9f130369892108e3d3b759d18d524dd37adb0e0b5f44ce3f249cbc24aac39b8932d7c6345f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9be36be9a441256d08875808895b0d9d81785d51ccd3838632716421ae77677deb97098dc80161ef0154901856db456ec7e72aeb6cb32407df9003a8b8cc043696c07d271540d79be7dcbbac64a5cffc930cf266815976981af143ec50c3e225ec151c203541ff9eb92a74c1a9ba8ed1b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6717f2edda3f36c0100ee86c4bacdff61bb45ff7a36f0b8929d83bf2dc4b54cf846eff52deb89dc57dd27045598166584fa7e00d6368d10c339d1da88e1867a7c848093a1892e19d6c353035f0ee7ebed335023a0fa8f37e61eec8aa316091cbcda065657bedb0e433e7436d3bb1c9692;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7356a18ea3427a027f9ff1f6523760d1bef865f31dd0230d308f151146166ac40c20963d4a4f4874d637e91000d8d533171e4659578fe1e8ea4e9bb538dced90be20fd28a60de03ee46b0cc67fed5e920374b0f5488358c0984dd9e3b67affac965f0cf2bd372ddada792921b3e9bae31;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fdad8d3d79e0c9bb5375c7593728894bf5ef0a9fd7e9fd40555a671e915789607dfd4241165f01130a7ef4062b38c48aff3ae55652344da9aeb525f409f23f71cdbca11bebe74f918d7d6f3f8655492eb571279227077b73d99120778237f5ca43d6e3462c6ecd65e7bf22165eb76c03;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5cfe5c6e8991966bbed4608623af9684bb19ee2ce29c157690d86d47343fafbe39755e38eb4e3400b1df112038bf5538b04ecc2060169034fccab3d6769e955db6f8da937f6730f679abca328a1cf67696fda7a4da69fd4bcc2ae4c1389d39b40e986850a04ba2196c238a5ff20746289;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h776bd89d3afd5482cee6439e8a2818afde9fd344f35c51e46c4bfc747fcbdbc41605a68baf40734566572c790903561556b5f78338694622fcfd8f10e3bce5ba69350438576a9a20e7e08b4b93529741de6636ebe833e0bafd57801087ba8d18772b66d366091e9ba7149f2b668df2b2c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hadcf037bbc145c404c6dc036c1a8768232d127fe4cc9be7c3c6e9da44bbcaff0d010c78ea670ca5f1bd61938712c372b2456949db8d8e25911bd36ee1e3c538ee7d2dbc26ca6b3ab055d914d3b6f974904d06e4cc498a3ac6c0768fe0f6ac9e7a6f71aca107b0a616d82ca0ff0db80d89;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbfb932afefd3a8c2770c13fe36a8a58f66f2a80b3c351095a4ceacc2b86577a86db9c2fc6376d57c6f0e649f63d51ffbab349557a349ce292107d841e79e68560543c928b729dcdb3aa18ec96bf7ea790105cb144c0ce36d0c6c459afebd2b61d3558e138326a28a07801160aed01b58;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h802e4187a006b1ae3401e18aff3eff1018462b344d27c0f9c2ce06cd54d080c83365b0d6ea22e0932db130bc809f0c7f401e43d2ad77d375ddb932db638d0afd65cb4ce93f1660dc49caa0dee29eebe207dd81128723ab009179d8ac731cc3a6298afc733f23bcf54c114aada3ea3d744;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3e4a2e7a0e0198c94bf3c98751b044bfa0a540937076b5eec05e3bfa6b4535928f39010fc021000f3a5d1deffb083b017282cfb5609330f4807edb2f908e455f47ff3c1234956627953f81bcd2d2f8484e10f6e90dcba0c9452bf5a55bb210ec09e633d7fe0d99b37c4045b885d28e36;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8d44ad93c4e50925bb72931cf7d0102f8f018c5e2f82dad92493a48384a3b27781e85287620469f68b33b2871e99760865a47973de337d5a448850a9f5512bf44fbe2270feef3d24c9ac640512d60d4b769eba295c357836bdfbc2fa71193d70e298932b0bba494366df7ba316fd9a6a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c98f77bd8e67d16e255a8fe90472afaa9bf61c6630ae9f5f837f85b65a47f373f5c2d4bf4b262503247f562219a124eac83db3633b3a10a52651833f7a513840fede6db829d0dc5c934fb0e4f9d136143e45d61571d0efd1ed2509ba118af586ec3cdf9c519ddee88fd9b8d061481c20;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hafcd2677d9f93bf8d7c896112046d52fcd7d6bbd449f21a0483cdee1b587c9b81060a3756eb77c6e3b7fae28393a09a6c437085dfc0aee15e6e934221231b9ce930c9e5987194556ae3fdc6d8e960b569419e338165e4558f3901b054f34ff8d2e8dcc3e274618380efa04d4e9abf96c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4dca953e338c3e81c7a3e5e0ec15169251877bac54200c051fae5cf46736f23e6c9d1b013912b0bc4c69c912474aecb7929e17182d7053af0a20345a9a02c7c8be3bb07c9e3c765afb04035a93b081161a8b6f7d35a630f511a710a612ae643c3da5eadf1fd1905af4a3bd3c59f015b30;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee80e1908ff699d86486225411e7cc68a37eac7d0be907710f96adef879fe53a7fa9106cae4a478a7b956a38550a4ea4c09972e60219ae37ba983ad461ff963f22981fb7f1020917982bb341d76f9d4f7e388ca26184321f4bff5f724297052c63271cb8cdb36585e631e976fe806a815;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47073e7eeca2f16d1ecc6d8f8310623dc84cca53c0bcd05c56d1714af3fa409b90bd46f516c76d48abab2d877aa395bf5f88c598bb0570ddf43d68f813a24e5f3893ba42e072ad39c254472dbc1a13e661201092a011488ce3d73b6d60797de56fee92435b2468b1e25b4191fbd650eea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h476b3c1968f45074fe4d5825887dd6e44d2a79ccfa89340acd5af17f248df036eef7cb66d024352e2bbd0dc9006515a343e7860d01eb3dba0d46927909130c2b0eb7a722bbc10259e9910a4467134e3ba62d7f83ffaac91c2d522dd83a9f569810600f7fa3c530a1e9c6bb53fff17f71b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb82288df0685a4ec1144acadfeb370d86d96512d0a990ada08a4d6deb9697ff6929a041456739348c1731f268d9932e8e84d8fdbabd536830c7b0568c3f2f63e30c993b1c3752feecda997b973b45810ae30971d6f619fecca944199cabe9d05c779ea1068d8a54d92e53b13663625d69;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ca99a8caad541a2c08baca6e6c493fd46e5686df43894da76690eb65c24b1cb38f69de8510ef3c78412bddfd9b946ab6a37f732af0e0530b1e9842d81414aa21bdf4c4106c6730fb8869b501397c6f8edd70fece866c0a2805cdae1ba3857f4e97af0953e4dacbb612e708b27ffb85e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1469dc43a0826e1e60053f1e4960c60653d265e3bc918606beb9d060ac564a9bb8b2ca38619cbf81d41e7db27c6d76711fa34c63ccead3c2952b9c1e4e2d49654be5dc79a3b139918d70f9664b7b1ee0f24ebcc45d660572c21f3dc1ad3f2eaa262d31a9b52554a2ae45fad95bfb4655;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha85333f366a287b18127c6e86a038a951f3a6e3cd01a3eac737e9869823e6ab68cb764d21cc031ff299e6703bdeb6e1a307c9b4d99fd929d7a05d3ee32b7ddf8e06437baef34f3a4f1ff88ba8355ddce660f99cc3f4a69d5b1e08daa19e3d9078ed2854a0e0eff1a6fc0c959055fefe5e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h295aced02a3d6324db563dc58e0ce9e5febed03c9e3935ea8d59bd86d1d4426799405961b9338cb80b2a311022521086e5916307ac71c3d4329210c8105e0149a96a099060f1c4189a69bfa3de3cbe72a8d00f5f7f89975d795e2c56e4c28bac2bd307e2ea409ae9dc408b9eeb39acc74;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b2e03ebde08a8bc54b3d691e37c828a408cffce0951211902e48ad103f487644873cee0343c2a86c19ac6f5ba67bef9460a1b535eab5ba628c7b4c2d22f3a229343a2f0a0486802c3242213da96d55b3cbd7a1321ca994827310f5e48cba5f5924e09af8fcf3533ebff0d2c781de480;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9271951e10fb5d9567377909a5ef616d00a42fcb1d49a037c565dc3e09fe634e437a86ba7f8977e74b251b01e3969454482266deb6a187d73b8e2e9177fbebaac76a6ec1e52ff0b7ed444668b07acdc488ce98427f4708ac7d3002d0a19d5104e29aa0731c2cdf9d4c58048f276b66b46;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha93a4370098fff56911d2af1d0653d5651f2988e4738b598b773c037a1e6bc55e6c964ac2c309956e07dbde5defbbf5ee9cd9c2aba8c505d5d13c30a1e479d303c710c1a05b1fa6e59164868c6cfc1024d4d7be4e18f082e6328a74f9a22603c4b7abb1e642b0bd5787dc37c2aa91136f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2c327e92ddf7f95769348ef68e739b97ffb010bfa623b1013fd6bc04a9def0a5c7be60a8967e658ec284122a4a53c12f69cfe2816029bbf06022da0bb9fd8d91cb7df6f39fc719449f8d2e2f25850658f02dc5ebaaa3b9f3b18678529b2778740cadd038a964872b64641fb8f64a16f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd878dfb274bb74dd1f29f6f1306f9ada14907fb6fe2adf618189fccac27e94340b008cdc09a11f0c87d2e2f13358b9b166c87db9ba4f65d1ac6ac2dd6818f97fefa6940e02f91005d285c43ab7ea168e8671c89c70110e728c454ebcde2c287c576044b4ffa47e8863d8f26913315571;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h812bb8b18cfa06b7ede06493eabae315687c43ed35d2de4018eab4328b64198adffbda2a8b3bcab2932258ee96633aa335f3d70c212bad6cc81d137a54e26dd779ef409fa815c0e2e6161e60d805eaa65716908e29bb926217117af53a3fb72838d0e0204b1d9eef1fecdc2f585dce134;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8100fabee795fb8e0593700a9448548fe13c9e6a7ac0fa44fb1b2e08db01b0f5d152c999299f341a436b3e18612ad922e0198e90665d81db2f7197d75fcf887d4c663d6027b90fd1722d15be9a131f68e8fc53f56318d41ef5a358b1580a3d6a55ad3cf4310e8a759d3213140de3f75a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2466ae36f5bd4de0fccd40e664a6001f0bdc395ee6e01e3119948d6bcd817a1bd1f336c855aa51fc3eaea15ab3190f0d4f1f9c413af137cb7602d25b8f948f96843dcc0da79c8f27ff2f8dd0c98032b488cb37af020a168319e532a1c243dc5134e6022928d86a6d7373c810308ce459;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf63e1622e5a6620dcce6e0c00be3c252818e27d5877fef964f15c3fc44db697f0128f61beb7f67e2d63ff3a2ba24a216b06ef232d9cd2a73ce10041a2eb8df0b776bc6b22e56c3455fc319972c67c815f0417a4ecafdccb40010149ba96fbe5001a1775337055862a22a456900c5d0870;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52880e427b8ab713fa46a1ab1c64b8a32126f4fa1714dcce4326290313655efd5c6e59950cac74825030b7724d14134959aa0cfec83c9317b21b91aeb7eaf05f7a7cf8a46ef8123d30a2e6de83c615a157a53f0fe49cf5195ccd522329ebf1204cdf09d40e3de8f5a8682ac4f04fab099;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2006d42344d94fe0e69a76be5c369242d59f69eb56057048e35ac613e1a72c906a7baafbc37e413410eff638ce19a2ff9162d902e842f079d881a9150a3796b721d3f300ad1e9658f3754ce38e244b98846734f4137cc8e9719c14a1066165fea64f086c28b7a4a72b4205ac8afa0a48b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6470cd40f0ecf0764ef5ad570754fb07a3cfebfd24dcb5dfbe13d75e498ca8655303bd87e9a66e3306a3ef540b1155ae96a4691b255009764f59e9a1e0caab7b1534741817b1eab8ca9dc8f30ce5469698bb8fc66069b767bac532c5f8320beab187fabe4b13eb2ba9383f00446dee666;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecae8a8cfe75b520febb6559fb3162d1036c2b92463c03f4af9f197e8fdc00069b7d3879bf47573988d0683e06de49b558201d1ce19b16b329d3add53d53f516f85ada9927c40f9839f2447e752f79e841b10e54ed02adfb66184d5ae50b225e5b18b365bfda374699276aead7d9de4c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd40402d084956d7895581ef581d2d864bc54aef05ca75580ae4381d63dc69dee1cf673423a306ca9d6c9271e97531add3e9db9226fe6c7b7004b2f1758d143897d618b85fc175ece84dafc8b0aeee10ef5f34fd7ba1d2982814363510a8eb4e54015a090bb140989ac327a03083fd9bfb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h262f7f180b7d059f8f2b55ad9b7fc236851d4f842777c86c62fd711007639bd56781a787127c5de5316ff42babbfbf9cb72f6c947a97085c402f08c9c727ec6be99641394daa53288e42ec6d1aa0111df5642616dabae9febf28829fe327e088cd26222246039d2c557fc9d713541992f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he542a6621d3aea80cc50000b33138178cb3ac03775fec948c8d273e0715ded26089288e6d307d21982e1612f7b3667388e76d49e5d82feb9758fcad67cb2bffbb240a97daf6f3649b1b917b0d37acd88a2f371a9def354d7389ce70864ba0b2bf954aad90a7902e48dc5ae7aa274d17eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h746b8d34c5cebe19d1fe3540ee8551d7d8469be21d820a91ff160560651f8a7d220b091a690ef8649b2fd1a40feeee5abd45d4d4dc848302249f0ac2981e4c3fba6f0a71a15d30348c08b3ebcd30ce4cec2d7909671ec8db7d50977633cee4280a79bb939b2be64b2898e464ee0ea5e9b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7021139f74d9125e68c9bc99d0792642ffc678018ecfadc59096dec3684ab6fbf75a5a60f56514dd0193f4fb84340ebc88c9dc6889f1e8cdc05b46d551e0c6ae7989c9cf9c447a38aac96161298644dc0b61980d41d2bb3a02b1e6a8309da0c0f03ddc926df508b06cf860ec8f4836b9d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd4650a03401483b12df95a34431ababd978463cbed7ebe29a0c5986659176c584c5641aa551022dbb5fdc709db70f6cef179ecb65a9e2749464e5ba86f557e1c981cbf3e8898ef98b654863da918ee56f3ae913d91bfa1ce0ba03b03cd551a38c4ef6f8f769ad2abeaf13d35b6e53f42;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc24cad7c6b5379e5742c69cbfc02be073003f733fdfae790f0d568c56803b254444076bcf75a7b7ce35356053f526522937cc3087ff13fde13c8c3a65610d512578eacb773b85368e08be91e7312ab8c93fa96092532c11d216063339a024238f2f6e0c3890611c76d063f023f36385f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha700b9dcb7c13e16ebb1b5f39e8882e8de69c5b68affd27b8db9a19d39d27e74c9fae07e6a191ec41545a1cbe4155c6ae47580aaaa9bee0f04636a0a2be3d52dd495c7ce53eaf30fb43732b16a834f3b9d2b968428a5ac615842bfd56cc6a609afaaed776210ce2cf05427575a3dc9be8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h845a9f60e5368941a189e9d5a350076e634777303c240a9cf65ddfed8aa8279fb70994e996883397cb8d96fdc298c8a3c364c10338da53125940f662bb9c360b24e36e7dc42784c38f746f56d888fa317155dd6d1f37fe27206014ddfaae29ff45737147ba5ee1f0e6239546a6ecc9d9f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd523f992f483e8bbe38e90915f17e2de501efcbb3e09692a76c60670bedcfc05784b3de3958d144d08059be13a0aa77e217acb51b2052b8a45e3bc096a9085711712a10b4ee3755718b46e1b180158e50f0dca368c56dc9a5ab66269dc2d91636e79b9642a612e03995d3905f87b4df75;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd163d60e2ca86578a7a22363b74d2ba29c5cabeddc9162f43bb7dfec1258c834885b7c483719fed08d33f340c922e686b10f3ae81354bff777898489bc33f249a3deade004044aeb36efc697eac5f229f07b0cf4c3fc1256e3019d99327c33640fe3309bd425319ac22a8e4fce194ecea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4177454cfb8ba9d2af7bb514a05c29a324184828c333129f52bedb2b786e6bc81ef18f7f3c9d06c8edb9280c5f527708155d50371efdafe1bdaae5ccdc3ba930580b26530f2081700bd49942a037cd25086319e11e433658748b21ff4ed4f4d7cfffdcab58833a878e25acb3a1000dc5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a2336297e0adc014fcf4300a942e85a65946b22ff7cd1034ed5b06a685f191a888c36d2aaef9daef0bb3bb4d2085b2da1e9359b3bc625674ad96b6c655ebb08ad53598016f610f15976582566b64332edfa35ce05092a1dd3c251f2e5d795c21825e8f1d9ab3b01c258dbfa202607c2a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdda5c66746a1f2528b9ab3f8d714ac6f0add4bb2a4cd802f1ec8655b306c6e6555d2e8ea6d9500833893fe82b7efb9729ce6c37d1cdaedc124c12960f4f879605df1a57a0106b902cf3c32a95636b9883bd38eb2a9bfd842961a542b9cd9437232767bdd9f23d4d1e78cd65cd7bd7e539;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7871b2e8b1a43b8a77616053449a28588aea627fee541016a2b9803c1c0e8315287216907a889f4cbfa933f8a60cb6cc5acfb351828f506c3ed8f8267c31b35b9a67dc2fcbdbaf9faf159110395bca765ed33bd05fdac627e20584ac5c6e64231c9b3a30fbb32aa98afba61e873318c13;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7fcf10d6603851f6d797980fec33455444befd5499b0f7f1b9d78d60d35245b98371b6c77da0a04f4d58a8d6a62df910a269733a41a0d2d691c369070d7eec42aae6fc5297b5fce8b31e415f9ff20bee9e0b04a3c315ff4dead9ffb4a3297ab54d842ce33b6da4a948f34fab880a91c20;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5eeac3baa5d09811e153ce29af978031f237c052295d45cecfc2043e38bd1a4305966e0c4dfadc033936e42d435aa9083477f49444311f1812d113896aa1da956221291bb5aa32ab4459208282be62be4e128eae030d0349ce2f301f68e4ba172c0805fb5c80d26ff7934170c5e817a14;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1821c6112bcf54669f56156b283dedc5e8bdede3faccee83fa03ce2a701796138a0c502824b37dde9151c35ed079399a063de50b7dcf258ed3db53afc76f2361817bd983476f1b24a9ee55c2cfd21e06302e11fc5a47977de94d622bc8d58f2aa8ec6fb481bc8a0a537b4cf12a146931;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbd7d514b04095caada4bdfa2087b274c347c2759e1ae09e759d3cf78be34adde8361b21321b423019ac63d39ed878f16b56d1d7d6ff586e7b35f0edc0aebca651ba44ed16e5aa95adb52b3cc6cfb68410684f7b163fb4e4146f79933fe64bc1fdfa786860aa8eb0b48277545c2aeb8d0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1749d8e3b4c065713bd8f1f3545faf37a59ded3051095bde7d7fb13ddf34219dc2f5e9026e0e1e6d01b8544ae7d51eb6d7d450eab3ac57262f82827168af449423a4448cf0cc9adfcf0acc2d2a629e8993330659df821089a70e50858a241bcd5b705d9d03cd00bd826bc3cb136a3204d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67ef2dce1f5c428beda36ae2172b0c1fb99d33fcbb229a15c09d8b7e13a7e791da1cd6cf4003cbdbadfbfa3be42e1e7e26f271239c36ae077349c78182c7cdd44735af0cdcfc081780697974ffeaf308ce412768a083239298ae14692663933facdecf1ce9acabd59f49251a7412f16db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ba71ece697a3be8a64a1343915cdd3955af74bc13be73e0cf97363ef3ebbd41bb4c32f36ba151120718a4ac4729ce0ebcf81eb800a4df3362ffc253f7fb89c6af3fcb6e43079afb598655df87e90085b3192a5980267c36e0eb73d1bda3976a5c0216bf6bffeef17ddc40447f40bb61f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84c472e20ad34b5d37ad94949677c1d912e4994605c9c70570eab3c8ab12cf8f67d0e642f3655db442211be0f41d1cadf84dc110d5fa9d5b4e4a7e0911c52c496d06811fcc9ff9c976c5b3ed3baf9ad545379b80297c0541fce2c702f961b387217714827b1fc04f741ba32086a638432;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15df10068b3f88a2fb01f49b7f697666d746ed02d77f1f5b9f228718d4d71fdecde94ba8c90c939bcdf578097ca588264dacee64330b5d295436d1966b6a14f1faaa0fa60fc1de3a665bc2f7b69185c92449a57e007cd80bb282b357ff7ebcbfede661ac37a92983d523d5d584f57f16c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff2e5c4c1c6dbdfda7898afabd6f504d981f05f5cdd4608b2fbef9891e594e870eb34f834b238fe4a20b3b941f051cfff030eca8cc642785a62e5133721ad2d6eda6e27755c3166abd9cd5a135da59269c0abd3c93fde76d8f47a491363ba4b4c87ae7db0d7b6d06a052a4e0a4b4cbe9f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4142d5aa83fd1f270676f1dbb888226a73a1f97fa5ee42c504cc1c0827cd285a77a2639a1c1e11bbe1759349838c838b916a603590c92cf2c1ca6877db343c05fd7e6b111f974b8698a3a962b35ab085a42fdb3a570517c149cdf0537d831c8c00eb17d5b43d17aa1dfdf1bf7af23a60b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ce4f65d463a14963d2fa22166478620c3d5bff5244c6b4f340a883b6882d1a7b97e28d2d52875f4b87b5730211f7ab4e9a64190b119952bd9e23f23cb26851f681a845991730e83851ed76a70f01d20a59a2e238d2bee24434918a56cc5f675ecd7fb6bbff04df55452f08d2f2d08894;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcda48609eb48202bf3d6365ee787a8c6f39626460505a20badb3426d5d3e528c9e9d03ae1219f73b40c079896f34a4f93736f868542da8246d540350379e7504ab6a41fb50b2578f837d68f3130e05c8d0815d60b0f32b274629fc8227678b2ddc53492c28680fc536a75d1a3843e649f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb1e37e3e7b7d673902d99913d2cd51a2b69a1840bc6e59ca896feae8b01dd03e71646d7dcad287df2b98495057a9c86cce3654cb7d2f0937ddef20e5967960249cc669d33267df240752dc8dc940dbf705aeaff6c1cda57ae342991e8bd49f38529e0d71d9c72991a1dcf82cf6238092;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab1c77a37f76857866b629eb8a3b13637bb245b6110f78a0d35fe7f3ee2662cfe1fba9ca8c90e67d2dddb569de6321dcad749051c70e0045f9d281102255913755262616679fb07bd36be55dfeacc1121d43c07cd483164e7f13a2287626ca2861d47d0006a1b378ae0770a6784834da9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26688080bdfdaaa11aa60cd111fe6261098caa212c35ff2ba71101030569cfa35981ad29785e603caef88063be958e35e38373adb221f854663567f407e79b08eb4b95f09d44054936ecc480487d58956e0568d60b62099a03e0e2597322772d7b3fc8d209015c4a487cd764b6294f704;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e1b80726b28d996f479d393f3a9e7899494f93ac97a022af8937332e88015e28c11af924b64a26f4b8ff80fc11f1ac96713e7b300187b24fa89769409314cc20b5d14493dcf7b0379bff63441656d4824491c0c7cff2fb897dc9522621826650064749a4c9e47ea4d91fd21e0ff9c056;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f5706858f0b98104c8ea959eb024621338e1a4f8863f2fc66707c9cf0f28107112167733701fc44560177c20d462847ac912f7c014cab18a677b5724228e3ba91c4cb40cfcdbd7a783f239fb55353603bc204a1e1faa72938ac77e3a06caad6c24f9ed13a052ff9465e3c48e1e15dec7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff7d0efa01de8979bb6f3212ba9b334a9557f065e51949258e5b9ba85c793ad42c236db283ff57df8e06ec5616464e977e81d4e9c8e6ed865947c5f09f435a5631a19ab2ffe4b3755e9228c6a8cfbcfba7286535a5daf6c3715bf94a3db1f7ed157568b7a2f73d3ff2d9553de5669d5fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h237d90c2f03beb58a319e2d3ae6715f684837382827b3ff874bceb3e0bd805dca3801636fd8fa77f607b642bce50dfea145e65bcaa2872026457256d37ac7c5d291208fcd062d45a2b50b903edbd8ddd54d3e6beed0d5632432e67c5263829ea4d06df5594dbf2ab871337014552f2861;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4d57f5bf0c773a3a5f9175a4eeec51d4febc283748344aee13a6834ead513966eb511c70692db845ded3866a997cc2075ffdc870dbb7e5153428c5b1134484eb8740d6b05460b35bef3b8952c281473d7388ff3c5bb4cd13ac9733679bf6e37c59b0848ff8cdac224c9f6ad5ee64ddf8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41bec1fbc15dfc6a4d91d8bb4773ed36c0a30727a7deeb88359c467c7bcd329d4b8dc15a4aec3c37be9df24e315296651c33062f279ec8e977133f3c1d27389f1297f08f91611737e7f3713c35789fb617f0858b137e21953739f10e6f5681e992161e4d710e6ac80e988da3ba653f510;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb670176a856762efb533efaf51148c425efb9cfe8e72721e188dcf1356b6dceca0200d1a3164e35370d11b6ffed1f6b4a608e165d89c1d69f6ba1bc5d36ec5bc68e16d86c99b2ac91c06a8721d7c3caf4acde5d894c68255c4374b1c55461578b2a2918ee7852676c7039a7bba6bf9f15;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37783fdeff640954047ff5035e4b2d4d13798e27f9d1911655f9b881f596730004a5d308af18ff2ea311466b7671984b3e10c8fbd1c8b1cd01d06552d628eb6ce978af21ae21af168b52faa9a0526fb35c717cba7b77e8c59ad96fbd17cf865a7bb8c50d6a5ded0e7579ed88b0b96abd8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5aab1b7c69b92701d5e8b08271f25f94cfbd4454629cce0835d8539aa86118b85030181d6b62e13d0ab87dce2761c00f7f8a1097ff007a1bf1021e2296dbb456e15077169118fb090ae2026999761550c3f7d6ac4a66fe54e111961f579a66c6f26012fd38475f98b677421f244e6679a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53c4207b914ff5ca2846801e6b01aaa6bf92ce5cae1eab240120c7feb027dbaa770d03f178dd14bf085286d705d2215b4382fce42f3a5e3507d5aaaa7f9555ec3ab73a7ebec79e02f98d0b4b8fb82cf44a40f3dc5fd048d76b4b3f7b7883a555e5fc84abd982925b2bcb2e1ab919e6bae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6ed1683a50d055dfba0d0edcab9ad5975f84996889c740521c668c4e43ff72f606bb32735c710d4b9e1463beb311cce8add1ec40b0fc74c83898c0a09a9a74040007e11887316cd48588aa2e6ccffbd30a39ec1d14cfcbd5b927f2ef98b3fe1a5c9af93d24098d97c336237e24c06c3b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc04f7dba8987e411b61c6659c2f2e0f8afc59f9b95140d522ed8938665a7184c7ab4b0af93d58a9bf4a057064094fa45fb0a8720744191718249946e1f55f7ca74d9feec57f4026f19112b29a9f330663f9806a18056d2d5809f8a94d2cf5a1aa3c08ebf99a21bab074b99e8995b6dd4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf35cd6594bdfaaeed972721a9a71daf6caccff3131f3388a772b9509497c413879c0df04a20af6710dbaad7c7ed402e4d7e0069e6c814f441c32819573758368f3c058ebf0ed74bbdbd9e9ac082290011767ea69bb1aa26bd395bb41370b8d9325a5b42ccca85354872d0af17ddd22734;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e4b203eb540069234d42a13c0f2a017e77d746e9a1e4452bd27ef5f996ad2e9885a290e80a04e5d883f3c63f4d9fd3d9e03a659bed6c14d3b6ce642229286442d66c2df91b6eda17c78136e7ddb5a44f0c4c205d2f39f4809f17c971eec007e5152e4cde117217a035c15c98dc0e363f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb24de8e11f91b03385a27ffd981471e1e63962be27597cb0037789a921bc5dd7bc61476eb6e14b36504261e50a80e0685a84859b7e911cf995d81e61b384f83348d12d2d3188b964c27059f849071216bddada9eb7e63d10dd7d3f7b75226ca905c9d631574d151300ca7850e597658e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h421ea2ef7f085b20ed7403c7486316bd09986f510a58b7bb5e38691c1ce89f346c69ea2764ba2484323112ce4be30025d661a3b6cbcf10db2efa1bb900e63936009c3bc893e467e4887e9e730a7fb6298d5ae90762ec2f3138a557bc6cf58897597077bfd0f5d38b4417d2f9459ffa5ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96c45ba88e9c891936cdc9b12297903830b0779d3c7317e9a4bce094d361cef6d5d1feedbc6af367e4334956575794d180dba9dfd39341b66f1182b57dca52464d5cef07b2d41558bc6326b6ebb9a2754da54f22fc991730e80936156253de65bb1256935b7f84caab3d00b56eff3fc92;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf5a84bb8012e14d1992781abe93daab1cdd1478e08d27952ef2d0fdf7ad0b0a12c59ccbe604759d8ebcea3bee65bdd7fe7c10ae9c81a6e763534fb421ecfd16489010c5ed90fbf216d0d313e5ac73c90ed9ae5ce1d33c7b7e03c1816dd448394a4c5743620e6ca38878d7a918e9d9bb9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f410199890385fa876a14e74afecd5cfa8dfa65f5cd7cb0c8da42a9042ad4460d23a9020d1319909aad069e86f7dcec5619d4aa13eef59df9d4fe526028a223cc6350fdf94fcfb7e159837132e8e2c8e0a7b35ccdd3899c1a01d7f6f0b0a4ea39970d296ada334b15a921bd29c95681a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc241982e6c5b5390eb78790d7c6adfa3762ddb5be50b9324a03aba703572638a2bc931172040140f0b85f2617bec141fdf71a70be0edbb9a9ef178b2f38c10d59ffd92d0a8b11fdd11b6f731a3a47a1e03b816af481e072c19d5680fde19f96981a13735c81394d19731e5f6def4fa985;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb2a1b8ea99b2dbf8afe6323e3636c89daab6cee0b92c7daf9d341fdbc55a3b10af0c4246228f4f8c31d3163334acac7371ec60640710bd5bafc400d3ea6d16ef25aecce8829a077ed5191a6eae3a8466c4ff1e911ec60b73b19e6e3be05c466d045c7f82121ff0e79ed4bfe83ca577c5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e9dd49f0a3951d7dbb9ffdd3a099add68f72643a8923bdd79530aba0a85d8d8f9aa25836d1676b8b7efe337354ba6eedcf1175c70206da56e5059c6348b74e0ded15d2dd4e7c37e7fb56ac4a2d2086399d47922ba230ebc7c2ff192ede2bd1703ebf8d4a0ff657013d0523796dc132ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf467d3a833ce4c34a159a27f95e437623d178e36da37415efd40d5b4b934e7ea915ee2ebce33cb14b6327cbf4cc884e392fac6f07bb09df3c99f435aa2e45d812d187d389be581ea3c07b94d3285d6c7219b1a28375156f730604ef3a1d6f693881586b55589689efae48797b701f56e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedbafce7db98692eabb19a21c8ade98cf27ed7e47ce4ddd0c593884b28d48279057ee75190077d59089205c3e60292ba1bac02cabf833452404b946285cb5fe28157616a33f4837c3da6dc682c0337c321d35dcc9ac0ba0a5b234f6d5303d8a875a9d7c32cdae062e5c029cf091a9e621;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14725e04333efa97af8d293fa49a9ec52ccc2756bb24b37fbfd0ce289199acf87cb9ff3cdf3575010f69223075423155c039f76e6b0d83176cb46fbe2a98648f3d076d436b052290674a12f5d8f3283dfa79ecaa378e05c13f204da1c716f11fea500fac3d151a3ff4d64afb9bc3ce4ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a982d427cda0a4804fb9c5cb6b9fec11f0f2df9560bb03b0d7d2473838d221bd260c6d761c4ede9e039d857204e3ce94ed52b8bc2c1c795ff66ba4ad9c474a18055477262c4e2442fa9535dc22c781d36ae761fbd79a69682ba5b22dfa5e35c637d2562f345a47f1ee4a94336973ad0d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d2f6abba958392a6c825d6b95dc47eaa556a30442b4d9cd208de891ebd54511d46ae008fc6213c1ed52586cc635b4b999f9d120c511eb22048fef673e68871802d2c3573ffb03e06b2efa381adb094b863d0ff429a5bca026aee5d4102798772aa798a30441677826af8cb66217a4621;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d7aa47e337b1020b6187f2e922c42bf8a032d77abaf2f8757e54699c2d4877a18eeb0a21f4eda888bb46227dda1c289c4d53ccf4336581190efb566251ff1438d43a0fc3426d2356a8ce45fd6d4fe47cc27db497431c9f5ebfe91cddd6827d6a8405f864086ab7d5250719510df5d289;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce41228ea775dfa75a68fb9136ef3f2da82098c1e94bb10d38494e32506aa6325fb9fe610bc71725818a83834e9f66c288c9275a888ce8549fe0f39cdc3a50b8c3fff6683e8403c686218425b318c9f38900a1c237841e4ffabc01198d7e54a66a80ca4e596d030a97415414704bddb39;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20f364090a9fb730e7ec844aa658686d496075460e3203beb80049503c97a4e338e9d57ea66bfe0c6f857bd8ddd3446559bca48b119be9fac94e5a536288b3247286b794762e1dd022a45f80702a8fa10f41ada3df109c185e40f78279b84727af274bc4ea042d752b26e233a54210239;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h449a942d7f6ca696c35e5d339b07bcecd8844725dfbdefd7b631489d8b1d0d21dc23811c1097a7efb181e773e00e46ddf54fe4a3cdd9a3af6fcbd5ad7736d722b70a4dbc29e9d3c3d54bfc2049454e3f5293904ed15600d0db7d0af27ff0c788fd38d0071c8aae5ab77dc6604d7146e59;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0387c7df6859729575716add5f0cc2824725e3673171bcafe490a5fcf1233b5059964b90e01a3ea5335ca0dcd6695c83559ec708d9dfa225cf8072e21c95ce6f00d1fe084bdd22ae295642b6950dfbad3a498617f01eae4cef60a3c10f4a4c2b925a40962571d2a28650ba96ae7843c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3caf662c06703090f766f88bbfc96fe0b582acd1553ffcb5560cf513f7a86439d6ccc03a889b0842f59620edc84766bab86240498f29d9c37c9e595c346856f7a68869df28a49f501c44cbd263030828436d6824244a3e4fd162b63a6fa58e95a3934cbd3212a2bee7c0ade4a32a961c1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h714a1856c21bb54f9b5b7047322afa8d341f9fc8f51b05bf10a2e293f9cee2cfc640bc865ec59d6a36a3b774abc1422a2668727169ce74b0a6085600af832843e3e812f7cbb78408e2c8cdbb7536c23a7c70ee4aebf993df176a145cb0e3c036343db6643399386affcd1e2e4caf8ab05;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4b410cb4195049acf9cda1832746e7956c19dce2e14011cee5fb837d0a80d64919c2712f2b18aea1fbdecea002b26230f4a10d886345dd2c440e614cbf068733b97ac8745124b9a7c9537ef81366b7ffc91cae383bb2683012492de92ea8d4709c619f37c461c8495a1ccfc739e4a967;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c2ee28354092f300dad9af2ba2dbd69d1e11c5e1b0754aa3882f6a2a0e417dc4e81b9949df390af205a9989893e7ee7da9149e646b8a5ae785a1035f039d47468c54e7b16a2dfa201f9e2deff2885da041b3ce7bf2ab1aad55c0bee839263a2c4fb87eb30ccc270ae395ea152a5dcc58;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha18561da4442b3cd25986744f8b01226705100e05708fdca2dba065e953ade4ac68b9d6f184eab814865d275aea118d37f1eb1295eba38cfab9658ff17e56e43dc9bbd89a1d8ebdd15934c42b84a2d6e692409d00d5cfd2b3a498f15f3d37e2ac791abd21bfe7469bdffa6f3395898aca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ef1bd2afcf6ffa588897675bfab1e5ed34f226bd5a679e5f0f2788ac42bfd3e688d9ce37978b583c0b1b331af6b75d8dedc70a456f1047ede7a68d58eeece53bac51020a7fae9cf7240b340fd1a3a22aded5bb757f1c33f25db0999694097a9e21103eb9e87fa807a9d68540aca7510c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hefdac02d70415ec7254c0afffaaa8e07a776c2009149c1ef6ffd80c7b8eab37d424733737f73ae5a4b78bf4be07553cb2d2067c03e32d41e96b6e1dce99d1bb1eff524b57096c4cdf7e220f4484d089789a6cb55baeff46d0fc73466683c6d56d0d62092c75f752b3a3331acd1b11f911;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ce8418457ea18f54e691f38dafee3b5176122e5b687abbb5c49a2266d6a1be21cffee32b13253d7813b0ecb4ce59b9d005032f6d7859967fe38a0bf5f3273b4255ddc405c00ab50b67c34cdfeb5575132f5ef8bd8d14ee27c837044b98be26140af33a207aa532837f3d42514681070;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h361f0ee3855c4f9bda0169195cf73061606251bcbe13d63dfcd1bc72f70ce536bc77e3fa779bac8ee4a5ce1db974cb39c9d46d50d51e422cc4f900c9bb650c58ebb1854313817be2197ef1e85c524a50ab43cc2d175d36de1a3899dfa0e213e8c0565d59bcff29534f098eb684bdd328c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h822e098c46a715c4756a995d1c97f34422fdbba032201b03430110f932fdf34e3bd271d9a7d4c1a5f568e1c857cfcbb7bfb22b211ba4af002855c0f6b4cd32c1b694d927341f62c2fea903c801f8d70dc6080f08aa21b07bd3453f3d873820c1f6f6711ae736273f009faff4c08a62bca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haba28e2256930d809d21e59ca9cb2a78b0fbafe338ea8b71ad54fac8250d8d83719a89d24004ade55518d23d82ed9909b8a130e306da327658e0f00f74ab0c9534d80f9ed9177bf9f7ec2fbaa268b9f3f9d1e5daca89a1f567c4afdc1e1a0c60c9cbce269b3b5723ad0513d2e649b6e1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1defa5dcbbc5801b4e96cfa44ece3688169df25b434a34f4625fe438ea89977f9b732c93f68344f310a4c4f74ba7e2965afc809eebf5ff17902eb0abae8342959c554378dc65ed99c7698339746837c58129a4705046c6fdd5a8923facaea910102ddf5ef056b7d431b007db2ba8b9a4d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ac572c40da25654aa8a0d7bdfe2a826dfe1b0634ea61ab19aa3830ba0c05bf59ff552612644a354607e0ed1ddebc79943f686f61764994becc3a6bfe2ecd3048a4853822765878ad9f3fa25ee4c2ae4e3b90388072a12c39a8432097c7742002c482ef74e76822e77492b860ae12e761;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h940e1b723351d27bbb3581f94dd7199e8efe22f81d26b534d55dc8236def31883e69a69a170cc0cb87d831e85a589c651dadd1a35c833baf1377d1ae95b2fcb4ab95bff65440567f9de89835fa92fcd0ec271d39d0311405c6d983b21defec3273855996d2fba3effc26fbe926f071e14;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9027ee4602d1db68c67112248f8427b0b08812131de61d0d0d66e730607fbf8a5682a29c0a4acb6aa370295cbd845bccecc866dcc6daf2ab217db42ef2efe76ef467b45681af64c6e84f829fe6717c27cc7c844dd4cc1b63ce0ea9bcdbb456b329e1d93ae890346c7407b2c0867e71de;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h463efcf5aaa442e21fb02e0fb71e883894fa079816e50eaab921f6b5b1a9d3c45899a1fb03472fb920344267cfc905a7684e699e36359000bebe6d532cac703e8379bab62007dad4b287df8ddba9ba29582e2c924b8962b932a2ec6eaa27feb3ac726359502383c6d32eb135e31542244;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbd019778d5fffc90d2d92e2d379c8814bc8f56fcb750f5afc48c8f61b1cf5206b040c18b7c855d6a0c826f9bd311c2c1bb4bafac4d83b573c9c35e9f1575f38207bc7c6fb2534f103b79ca6e74322732f91ed57cf5b077c049298fda76daabe4d4be1c261e2ab8d95f36af29512f95c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h960140096955ef3b9ce6c93380147e5297812d8805ea97ce8bd7e1ceeefdedfee532bd97e2b6b331bcb79745de19f16b257d74c891b9d82c022deb66a3ea482b8f0ec7709664bca2f0a41178dc0a6729f0058fd3d107b69dfe5650b0cab509d20c40d1d298edef81127d2f17c9a61060c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heda647f37d7c942487e7bd19fca33a160429d01425fedadb5fca19e5fa46384a93aac5f9a5196187a3c27d4b2a2422df3615b243d02dd9d175e7a5d5d13b68ba2d64baf0e19dc0ffdef53b2a99e1701cf8eece1e3f45c902579217ab44bb11f293181bed5de012da156be6dd698c8b477;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h985dc5e9fe8fc2898ea902d88b2942fbee9f808052b35ca619bdf88c94967626dbbdbd217d3335a1cca3b2397b36e86c12a6b0a5b5a9289aad6e2e2593b5454963c5b846d7a6a22ad170879c62833afcedc04469bf774227455f7ef2ce100342e4715df02b0beba2b88cf66db7266c2f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h533cbfc68169d25d301c420fb93cfebd31cba964bb0f98cb6c0ae4d99f34ab5ded60795e25444ab3e2e12d3f5f163414a119202a2d2b40e42a132bc1ea19def971ea348a3d7505c9b59fa1f1e4fa10507caaae6f8872ea6c8f9fde3b29042a48f20a933737a00779d749fc3c9431e1e65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70eb9758d976669b79087ce3764fee63ca5228b43835a45313d88d6d11eba4c55f164a684a2041c7bc414f190ef0fbcce654a84e0a530328d4f89da81f26923c51a35c02e74113b72b5c21121d7d0775b2b48168a58f9dda274a675d87704e5c22881e1dfe9ddce6e8e3235c7ce56885b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe96f24cf21c1ac1b2a6eb67e22456cfda76c71f690d588119473851e9b170a6a7ec41b01fbb9cfe3a1c7490df4a5c9c00d73890acd6d717db7f76dbecb1aab0039eef9062c738b0ea718db7edc21902b987fde8eb8299fb3118cda9bd04cdded7c590d2c79620a2b6f4964839aa753af;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3bca329b28348d1fe787a112362f6471f66c1bb596d38d7fa3742ff0083575251cb2ea8503c8722ebd04bf45e82c7fabedd1d1543ce5e9d09ebdbb6e0bd406ae5e94c36836e57df7492bd3f732f72f9a0556c5eb3efbcfad0b1f48aef019faf09c17a332fc9da765d04b363f92025906;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h255e25ebf6da1d1c624597a92e03c67ee466073f61d8b8430fa742036d4b92885c47b6c5ef6b3e41d8228e1214e05fdf3e02a21cb34289f8c875af5b81fff669ab06cac533bdf757a5a45c2a2c5af854ffa6902c4166a07ae080d9880f5737d4fa94687b11a4613d46f9cc74a2197d7c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7833adb491bd533d101b72b2eda36d31ed636249804d032d8cf5c1191a0b894ac860d6a20edfa227df598328d399ac6432da281c6700a161aad19a368770d3ed8893715850f3d8b385b32067ffb19a3bf30e0dab4d646d03c8dd4ec817e1aca4c709701191e9fe2de64745495f61113ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec873a579cb07d14a28028c74ccb31c9fa6db0578b4ce640cecd90e9d1655e87568478ad7129f02c68c4ccdc2d7a53e6a97053b6376eacea0f1f97f7b99333d3934aa2a236e0a3851f05842bf84d87670fda0d08c74a63d37e524ca6e1f8a043a4a759b87c7a12ccfdc629dfbecf76535;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h271e37dbf3e067ab07372143eae4b89f33dd7f1563fbf3fe7a62384b85daa51ac949ac92d1f60004e939582e890440dfa53e43d1115244b6736d7141966083ecb6195f5bbfaa248e0e1d5f18f76d8b70ba8831d198942cd7ddbd469ad10381939f466c3f245360c41d3516f9e929c0d46;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h371fa348f7f8f9790a6cbcb92ae698a6cc61a6d6c974e70e54e341741b86cde7e87f0d6f0bb06a7d96c45633c8c5142345a99100dcb97319e0f6fb0578d43b9da02101205c9852970957816bb2c59b4c89128f88aa39a937becb8df968018602d59f92c0ef0dea238b9686f2fe62f1f6c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfef2977b0e1eb65ba98e17e1d6735383e09f0e2c89a09875d51f346d9792eaf177008f15ade358f5f6edaf37c95b728d68126c2469da23e6b436a2d817ed7fdf26edeb87f84c2792b21f2d40cd6ae69813632e7d2f13de6fe7271a2c886f69446ed8d1bd34a9852b5c20d5d9cc7d778f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91423f065e2b98eadb9e82e8065e7897990d813c9ed394bdd066411579e31572006c43e8f39e749b89994c95ffca1e3ee64af5669cec47691e0e1d42ff51995966a3d13c46b8a0074588c7820c49bb5f6abae9234f9580a4355cfa94b5a2c58b108683c2fcda189e8912a8d0fd60045f7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0b616340b600b4ddfbf5d6c86008c438d6c52c394ac742fb1e89fc84864cb96b7742ba30857d9a88433484f6a1eb915cbb3cd8575a97cf4e6f1c102bedebf52efbd515066b74df9f9ebbb9143f32f4a8c2aff1a9abc2c59f99d38aa212cb10e43dbc583cf5cb1e3e6e1b8ed4c56837a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68268cea85fdb5f7a4f1d8d46eb796b3937b3b6214d732d0d98b40a54bd4c08460db44c368120abbd8515666d27bf00c05bb8cf1e1c5accb0f6fb35a589605b6a2d84ed1c86c5e8c2e5b8204f58cb93682f483d96ed97de43d4091804a80851da3ae9c90401fc19ac5e5a9412b4e65f69;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h887b604a9938acdf6aa62861e6df909441afa6f4931ab88e997aa14d07c68ae4fcfc56022759be22a0dbcc74eeb70f98c8515e49f12a56478a439f1c86d9c17ea050ebdfe03e133be3b5478a4dc96620f02f3b37771def8b3846d0559b50fd6f5d5ef48ed2beea7b9f98f2298517d653a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce28e8c66785221d0cd71010faabb7298822505c613524a239bd60662178d65372b14891c156e0f6fa5152ba6a3e2cc49a5a94d872b422f5c9e2c698c7ef5c9dcb0abb425cfc1961850883355c63dcee1cf56227000c20d0d8b62b4ea8f02d411eb21ae6c48810579ddfffd60d8c4052a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36d36149c94fe8d57ee4d47e177248a22243d58bbbe20cdea0bdbd7a2b7323f376961e20e1bb3fa24bd7acb4c0c310b6c237b4e6440cf845a3cf524c109667994442a6a16470db5f3cfac063070c09297449106056819770941e9307eebcf78d306cf67ae21d8498797b59da35ba0b80e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h703a62c1b19de46de4664bf7c1200a68272af9062afa47430c77630aabc5b8aa2fea3827f024696858200565c93c26a3ea0ab423b49ff664ccb5b0f9c8883c2139ed191c918911286e9805ca45100767eb7d67bd866aa7319b232ad0587b58399c745adc092728c084863d3f434589a12;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9472cc41e0a0459d9966f7f7be242a02edf4a841b2f8696557b5193e420202cd12ff9bd56c3bc690c6871a5653fc9a9c613aedd9fdb78ff81a9eb602910226bf27598bcf4ea6a17a2944dc9b11a5c4dd6ea26eb2a689984a7e301872e22fa0efb3583b39179a7bdeeb416e93c5123924;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8194afabf62aa52062ebcc0c0ab2f4ba70de39ac9670200d92eaea27274545760bb14485879945b0e2036b47587126cde8758a4cb50dcd094c58ca5d7b560c9f7b2dae4ef08667978fa64ce806fe56a3578e44d387a929ab2e533380a7e7acd760722b06c9e44f5796be20cb8a4865ae6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf78541702c2a7cee0988f87bccebe8b2b536e25cdb870d62984790b5cd69ea552ffc0997aa968460e1c1dd30b5b42001e1354b77b32215d336977776dd17c42408bfdfdb6a81d482fc817dc5a5326e7f8ecdb3110e60b76cc2cc731a82f652d0bb25e9eb98bf1fc8fecce11d06d342ec8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce105a5f71db501209f2fa4e1376f6ab34c185cf0d4f2db2b512947e4c41bf52b23d5aa818e20b0f4f2b621eb63ab012977682b0b087794bbbe02ecee0928e15595c82c31c54d66c8e763dd5e1eac8d94abdb69283bcc4698bb3e7974e0c5fb96299ae9b0919c74e64e5eac471ca380e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb76d00cd93c0891523105ac6727282961056b0965b5c834bc008bfda292535f5fa745904ff762366727f4322d464fcf14a24ca8505a2549182ba703f2cc3c6f77b2647888d14deab6b995c6af141d9b8bc1df32ec40d15a2adf9b528d50f29809e1b8e79c8ce90bf63bfe038ef239a92a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6fbc48e0f7b4308a8784b0028353a83c68d7e575052a66ec0be3a451cd2ee2bb3a37c028bf47323a2a766e7f7b7ba2d09471194b7ebfee138052250f93e4f983d51a7e664b1293d6eab062bae97fd21f4db698244ede4b02d201c47c5ac1eed3827c7812fc1b2a553c7109e6b7a9e671a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h851ce58972e5388152ff83c67e31e9fb013ec2ca4f1331b04491468b803bd2f9a571ca3fabe29db2c02adb8046155089ebe6f9b370cbe1bfb50cb41932fe5310fd33712fae19232e0ca92131ca0341e15f4ccb1b965c54d27ac20aa5221f8039afddac7cf435f2d5bf44e72c498564858;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5cb7658e5f0e093b0b282e40632589e145a53b8c7c726a14e8b50f4c3ef4a5b5e323c4ce7c12c64bec6d584107367a2993f1b156fa7065787d15f1c355ee24df17d8ae194d2ead2d2ba96b80e24b4eb6228dfc32b5d61240e3844fd8aa62a8c8d9821ec45a3d9ea06e392f236a44f512;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47e14231306f01bef99df5f6dceb79ad8289e35b657a4fa7c624c0e26afee57851484dadee0b597bcfcb1e78c14ac960c1d60d5571e49d1db03d786e1b710d8ac53b3ad2715b5bdf9c08f660d746b45e0e427b3ee6ea8718ee8168d202fca7f7adb391143a8e73da3c7e90571bb0778a2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h397651efc050bda757045e6e3eabdcc24a05ddac66988ba8f773650dc7f9a076ff402ae2d5b1ad53485485f75dac96dc056398279faf2f0c2dca3b0e8ab9381f7f019c2649fa25a01c7701e104841bf8020a5fedaf4aacf73607e377df2c55327b6b8ee14961a5b545f9f906e93b565d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c499d1339fe7236fa1d8495576806bdf11a170b89c179ccfa4d20c583262ccd1ae05b9f548e00be33108871ed7cef30d7a29175523b053a7432aa89691e233f272ec9e2686ebaf7b0a83f95902b2082f0a43baad3178eec075a82f3aa43d874b98d729030d894d19a6f567f7e617fadc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h675e5c9e40f26a8bd8cdb66995af9023fbed14d8eea548ec6c4719063d6b0e35e3cbab696ba2f514a3fc28433971343e69fbe5984db524c2bcb040c1e36ee91c22a157bb8f893a573d938863388bad6d90f12db521f2988c1df7a7738cd696357b02e67f081a7269020ab99744f8c6bf3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94cb05acdb168e1da91c3f8d96c14ab707bd28648b927f44afeeb1c32bbe52fef2a775280f045d41a5ef555c8a6b2fd9afabe729090de920b6b2d5935205e7edc574c5358a9837101dca9445cf7a584d4e769a509e93e15b90332d16943bf4a20d82b9cd04e65da1b00002c8b8ea34ca6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc40d70160e676297b3d2cd6acf149e796b99a578470970aa0a5d78a17b8bc1baff8120d14908bfaa7a746ded6387005b105ae0393e6c1a535413ce690efdaba1b1049d27141da4c74652fbdb1266e0e4071b82b0c2180e589fd6d313f85ab1d8f5e9acf2986ba33bde61ba9d385c42191;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bca4725ab038faf4538f9a86889131e1064f9e8a64d0e44326b97bd29fd97cf380cfa43a347859a5403ba6a68ec88975a4ad73fdd52f84aee27f8814a6748d9069f5c59df44f8a7f41d6c06cf20f22ba1fdc3b7387e04c37a737ae1cd1a508d725a7efc57a0b7be99f0d0b1a865889e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10538fea1f230a50c02857fc8bbf457706893c3d4b2bec3d599f4bfcf84a2102d7336f39f63a1d4464ee49a04e512b59c520ed947ea2ccccf7f1552f840107fce5b148fd5676a8f140e7988cc686f5a9940d8b9572a599d23a3f7ab9444b38ef8c90ec9ee0ff2eb2897a5b0b415e58553;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccc6aefd94f48eda1fd8ad8fd545ce69cde645e7f441b17331b957c7545bec580b59f3a8097d9c89b50a598b8aafd15a7ebe4ce8fa80e298527e8126cd578134d1a562c27052af92839574c16e24cef8a8a95373fab621b79bb3f210693856de080f0119ff36182929975050aefc2b061;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0517b908e850a293d8b37e6c759c317dc7c00c77250215adadad7fb25d22cf9434ff9d88eaf866ef3f3e8a507bb1e4468407ff5344f6c2c436a58df4e96f2a4a5ff580a08cd8d9436c35dfc266fc514a79a0f903bd82e22bc579975647331ff817e2f9756ec2b1ccb00083dc74f64f80;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70942f2f65550d456ec22677489b3e22e81304121e747cb3a0af57b71b853c56a15e110ea161667ab038c9ce21ca97fa49e4bf55bf60c887839b082c9a41ec48b24ae8fe7f53431c8841c701cd2a1c42d371b49d093fce2d4fd90a6ff7bb6aa2e2ebe032e388fbda00e38471c3a360d27;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b3d4af6b91bab87e2be4a45ccaa87298eb295b0b257bd062a9c8bd81e5a928424f9dec6a390285f6814579887f2b2816f3401c180ac44cd6f99ec3ca8523fac025f92d3b753caa0d6f77998e5defde86755518a69f7186b516f02259a9bf0b2e872c92db499f0f4f1efe94c78320f338;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5176e35b43f451b68b4a20dc6d8b30da05893e3d62d970e68838a87fe707b6d7662e86c9644432da1f2bf7a4f2c3545074b1775d2f1436c3128692869232e53b471e085e7e540b1757a9aa6e96adc819421e466d8bdd9409079c76c571f74f05f1dc34f9a1c930db4e7031b63eaa11b1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27880050b909e1d005ec63ef31340fc040319d5721ad701832c474c68a860528b56f6f5d5ae02f69e2cbe27d118a09f6687b99a56d58fa6159f8aa911f6ae40a0979c9f4aed24662bb00045072ac51474faa8146521b77abebd38998110a578dea852a74601e32e6be64f2032ab6896ca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf866f3a59523785baebbc2711a8f3d0dc1e4b5dccabb77f24c0f9986dd480f5167513915d3c0d06499a0dade7f64112400513a0db72c704f50dadfdc2dc97aa1e12ee6441b23539cb7d71e8cdcbdc869bb52160683d5592221b050c184aeb04804a8e8cbafc98e2e5bd8e5694045ac191;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h257cc81fb0da0fab216f3792103288b01f287b3f2d9168a4fee08013a3bf35faebb8a8a947ddbfd10a7cee1b3cd0542ed0b6bdf8e936d52f42c85258d158fcaaaba451354412689df2a21f55b2fb77896b70ebecc03fe9c92b3d8337098043702f5481570f827088b06e2adcad02977d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h347a29be02c9e615881b15ebaae00105d8b99ba2117f49707a7b01256cadffc8d93f632d213135e4e38dd62a1087e0ad36ca6a9b5f8cfe0714732ac0f939207bffad9e823fcbaf943aa12afd33410f8bd03643a7f64c2b30d6ae494aba950ad276db51226dea8f15102ad7bbfcac06bb6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3e70f4ff8bcf84086e899d1719cfe84400e6ec06b800529056d06558372883cda01cc920a0a474db13a1afaa3030d44993d0c14811b10945d269a083684836ef50ae2aaebb1dcd2e87156105a9e1ffaa4f77c3b38ceb0768f9bd3369e827873462db5e5ef49cd20f109d280b06dcb31e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1959cfdb96af938aee2620aa3bd5a2157066606a74464a3163c322dae32e2894d9c2b3f2ccab0afe6fa9d36e22063207bb826be17c9307b33ce8c002cb5af3f71146824399eb0312ef1b9dc109708b39d35cfb208760deeb0443e34fea257bcc487a114feecbebd8948772978655ffaad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e738fb5b1eca862c759ebbb2f0a41fc8e8ee2f1bb01b38cfa26928f9594d391d686b28256d412ee96c9d46f280e18ea326833255198fbfc963e14fe803d29acde2c2cba86a1739a3290ca4ce62834889be1f367cbc04b6fa915ea44a7cfe02a81a608637761ca89503d9d8382fe18c95;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56a725f9d9a087b45299f062195620ca80a23876bc1b5179462bba745a2c1b3283968633dc74c6070cdac9226b0874cdb360217cea3cbd8cd396c41adba071c735f51104f1ab3a45318f6ff8077d8cf6e02101312850d7ad8322e7c4a93a588c3c2e690cbacac881b7e88c76e749f27fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a88abf7f28b3102d1d77520c1dd5bd3b21a87748c901c7f8d467c7f9bde877d21aea9860a31324f4a9570d201f5cf7b4fd3c17dee3726a9d4256991e800a71121b1613386160a741f566ac0294f50474d2b4537b1273aedd7aa72841cdfcae6ce994a2ab9a5e6407c157814d51eafc7f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8735f45ee3d3f9a18981f26139f1ccb587a66d5c51d9b2c5f469c12a5fe23af2b1053cd9c59e66192cd72d8a6baeacff868d4ae5d2817c9d55a38f208245fe27fb7fb9f3de8d10089e3a13f4e84d7203cc6a8c35c83c9229a208dbfd0d8528cf47dee165dca4a9951b452e49293c91cf6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42d9591d60564167c9cca173bea55d85d4f58386e4cf36af44d559b599b1f2b341d0ad1ec8e0b774abe30ce9e78fb279ec048e8000cceeb029503f0816c3df0a86666ebf654566fb2c2deb775fd9f08c994f645feadd9c0136f94321c56280819d61cd335380773830bb2c3f1153e5347;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34c8702ccf002c964e2ff4fe8a19e779f4c1c8f1501c96a674ebd493f08d48bb80ce473732b9edb5fbe20598f6d3f7138701a8abfbc5da7c17bc218f2fe25face1e3742389d407b34acb192a38004f82effa2973e92359be7455e758f711e512550c3c57de4f604484b3b9ad86c5f7e25;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd92f2e7a52406d8254e7476fd588137fb1043520a8dd0c2a78a52f5bb3c79affd6742a6a783c08cffdb823df782aad4cdc24fb1cfcfd643a8539cfaab94d5436bc2674b19bf0706677f67c63d4d214fa668d4ad8ea8da3eff9b9405bb1d2a13c0f6054642d4f9b1b99ba7d36725291eca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5320b60e3f93b11cfa114e0c23328d0d7e4f901a0cec78f3a6ebd6b4746b1b9a8580724a6db1b2600d4cb0e607ab79a60895d1603dc899385a0d6c73788fda6a00a0660a5846a89d3f4d1c386bdb4057263189c3c89e1ac206923de9322bd6bc812fa1dc1b391ee8a29106c2b776eb00a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce34f5f59660328b1a27ec7616219f63549cf2b44e9e018cc3b64e14fe12b62b7e3f5bdd39621ae8d0da2b499d8f387b430dc76461fbf8bf273a0c65b4ce067777b019b1127f104156210abbb97fd4351f140e6f57d7e64f3a38c2fa71b41e4c83ac53ab5eb5bd61fb8e014ad1b6a3a98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf610022e38ac9abac356b64c9818a6590e523056843177127f257e9fe6b2d965c1f52471f16eb2378a6ae7f5a8937fe360ad283b5873b1b6dca4bee301a7e37e6eb9533d467160b814877161853f440bbcca371933d19d5bf64938146ffe4977fb8bc604338310cbcaf0cb59f7616b007;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9acc34152b526bfe54cf27ae3fd9a85d74c2d3d11d2b3b50447f33ecfd7c3c92c78e2b9783e1a45fc996842ef1b8f8f31f506da898d1045747d6b02389ef2f662c465fa30c6e52acb0571f9db567e24e5ad970362a7a13d4a8380f0a8af30d4e73aa94714e41621148dc02d1a188e98b2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e92b1b0cfe08da149e05d8f7af8e16ae6f600d7368d27bbbcb9f47995dd93bc16bb1ac1b960ac53335453f2db72b14d098fafe6eeb8fcfc238068152e63f843be0e5c0cc5e44251ec458d97117006b0acaba47ff177007512cfa596be9f896c94db6f09c7a293b0dcc0206c9d251f74;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cb87b0422216a28a1b8bda59ab0f7844d54df910328b0feb5abe689876adbc7dce708dd7f037a21f52ceb6855d57a3afb23016e98cab6f774c299a9af0ae97c72f3f97b5b14e6574fcb8417540888aa46474d120419698efb3544a14c33840184ea4c3a8bf34f9ac04ea339a5189db22;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc60f2d962c8514014195f8a4fae824a9d53c881e64ba7382fa9e9a2497911cdfe3ab6c83ef5e80f9123e8b3be4616e38b966c2200b4c3f4fa4ccbd18c2e44ea03045fff6a84e53ecb93b05c485b90c63fa4b3c7cc92617add474059673dea04e68dfc597df106dd21faf44e737abf5847;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ffef621d2cd5a58e704c6ac8ff9cac4f7e5950dcfb50d35d2ec5bf84e888669a7000e4f811fac0d4ca57d97ce5a480acb5f8079522a94dd2dc6a8f33f782fae182094e34bf8f131bad71d8aab5fc152949229042898a1cb1830a91641e69b83971c7d3287feedce4874c4df2bcf29b00;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c6e0a9c19215a26b0e3b273d0d4ac3813397fb26ba5bb79e897b6eb42655f469c23951e611db39fbb9b12abd010c4513c22764a62c087bdc94612e297261c5e22be04d3ebf98e64768bc53bf1f1fc9e24144112241a8d5e2753e0f4f21909917badad192706849e73059a98d94fdbcfd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a9e5eadb95d4ad4f0d2e33720c6f716084060712f52698f4030a5f2556db90b6d374fbaf33a85fe9e85eb3ce685fba617e466ec0947fb050d7545d8b8c4a587e46dc7b91c90dc8899dd08bcc728050571337abeae0ef824934c9a934fb363d942ef34196aac54da4d8ffd93525bc2e46;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd018261b920ecf85f5b7dc38a9009f63ab597331b55d06bcbfd1f771b9d01d7544f25da6b5e221be498345bc2cbea8eec72effd78b045ae138ef1e2ee482d705c216a8d20f4596c33d858e346f00d92d3da13909e6c955531f6426d913b0002892f0be648734c38c64a9b143a41fd846;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h362834112d36637300d2b0498d9be09642d01be804bd09a43758f0a0175c66820fb6ce7bcb786cad14c768fba7d1a1c19d9f677da402b7ecb9b21491204f43ed4d8199d0e248c7f9d8c9965acd35f8c1869276ca18ded09ca82b86d56eff204369f27d350fa653326f9e1b4324cc274b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde07709e09104bb0e5d0d4138dba800c54d3dd79bdfc7b546b129da1affc5650de0cf32848271c794e1d1a3de19ba35d69a7429f9fcaf7d05a1f8bfa3b75718835301fa042cc6eb7a1fcfb38751883988ae4d1bd5e60c0ae46a126475ec3509969a30de346f9ec9c2c1fa177efb735b56;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b7dbe161a214cda4f94258e7a9df6c0e2134b00078e2b9f003f77051031525a612ed01dc1aeb922fdef1799ac97ce951400633a9b4372f4bc15e074e4e7f6ef9f39408bdfdee98b3a5a7d46bfc54f0992d948937cb90733645c43d5c07e4956ba10a87f2c3da2cc98746f09c4d49c741;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80771f2d4a9a57637863ce0add9f022dd3d2c32f2fb5bc179ccf2d00a604e99e520b73702891e07a3a9199e630abf5608f43a24b6387c6d80d87fee275a5a8f068696c9808eb9d62e8fee9548f4865dd9b2e52f6bdf562e4b98acc43c21c1fc784cb57412b8f4b3cfd842dd9c34847e65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4df47f135a25945ed6fb075df6b3e541699a1e52bf3ae7a1c1e2b2a746f59985a4a70c4f797f0166692ff99e4a10e36eeb8a3e787f866e98dc1d48d8018aba21fa8a8720ece59cf0f7d43c6d345f5799e6a6b6b3eb47132272b31c0d0ce79ffab9d56f20d9743da9b68b1af0c7d01ac06;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93f5d063e652f93b3b40b0cd2cbb9ff346d1811d8a7292a9cee567c2f020f32868f37ab3b5a225471a05cbe789a68565a8059f6d58a7bd57c0f1219e3c95ef7b6c0db473ebbd93aec91ed6cabd79b92018e600d2fe533fd681ea751f022d8df8e4fe0ae4da316594fcb24a854f83fdf2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ccbf4edf760100492a437081f949fe88a7de2f8fc03dc2d5ee6873b37458345f34bb311eda219c827d6f51cd2ddc69b590f6fa1018d3dadc2a6ffa665798b6d4493b199dd96654801036354c140399c649b0b85142e9c6ee3c23ba14e878e1788c50b64ebbabbd16852fdc33f5767f93;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75fcba25116d7e575b68f0af8dd1633cd1d9fc3acb90abd3a3f7c1a2dc7189a39274c761c1934cd19f7f08257cebfb9c8361d1d272ff992053f31b679b9e3f69e39753cc0eff327f14154f55a5ec9da3641c824d0af197997acfa02156a1376677d11915b56dbe0516edb8e1c0ff595;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5a86b25bb7bc7ad3dd9da6e3f3d4ea9761c4520b8e3968db072fbefe12e54cb11c054afb85950c90c61574a2ac7accea567a525e9503c359cb609ef97be6d4fd041c2b9cc466815f57b9c151c6daa40271ad1db8993abb87af8e7278140eaef0e18eaaf669eeba2bf34790c1c60aa839;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73580a0e10221c53939fc61c5b209a038e9fc2f2e100117858ef9629dc483fe0bf1610af389a8b99f4723b34eb091f11690ba8baeb4e2c34dd614f382c9277c6e257e2dee83a8444c24c85ce606bae27dbdf13b7958e74b6748d2cd85443b3acd37155ceb3ad0d66ad534d3a50b70286b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b6a2ef9712b10758b0b0fd9ba81b3232ae9465a1986cda7c37926983f24f15add26769ec2695b8f891018273d72ef42d957535df33ac149bebbc692940eaa1bce025d78b391c139cc2710e87c18abd5062ad07e3bb922872170d26e846f19759cf9352f72c01c5d9a41fe2f817b27b8e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc531ace3a1362b699840a3f0dc06bfc196720a4d306a2df03db19dc19c29884a09e0ada4a64f937562211700fa5a462c7b092d5241525b92e3fdd774994c9df8b3f098cc147fd8b35abf3378f1a75406d795c12535d5017bd12dc699f3a0767abf261cf0d4278cc34d0ac3cd75f45490c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb661a98899c2d14533df799d0867110774881cc9031f078c8f42f0dd30d3fd0f3ddad3a5388bb1832f48125b3c64a97812ebe050b1c325905b46aac75709b0e7b3c9cf94319abf68e98390349162f517cd1c263ba75ce4b7a6a2a93d78b55ddf96decc44e2d5f573ef5fcd0027159ff43;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5297aefaeab90508a11a9862e3f5a1b3386891f7e15cab0ecfb0e14b4caba60ec13abd0e748e41f51f332db0124c3fc629e5ab1c8d43f083dab2427f9831eea392034a70d2713315721ebc753b29bf8b5039c0776143603dd26ee291b3ff1c7b08e2b1003828719f2fd349a4899a6659e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4441d033423b1f173fdeb3de8532f04d8d9087c6ea5ce39dab6e5666197c5db82a1795744840157228a64ce6031d0794d179f2cc9ca2fc2012b3cca35233b6752c515f8ede0cd55a53934ee6f1f200eae2ebfcb842eb78c657482fdec3ab7e6cf8f105813d4a7c7220ebdb8c96c930c4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebfd774fcbf85e94480139de9cb04a01316f57d05566cb126302c10f9ea56e70c797fd89e5e9cc91b173fe90cf8950a56b77b2783d25ee51875a3010a84bd341b911e7f77013a792fbe0ee3978eba663935933a1fca544c80258c271cb7ebe1bc746c79cc3cb47a0cca7f803ef610ae66;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f0a70cd5814485533d7177bb52c4331450aa8f6e297ebdaecfe6151538cddc0f361d01ad2ccd75238a7492d49e2355223dddd2fd4bba09bb64de893bae4d2a49508b54b274838a0e8e8f60401738ede96e55a213175a3633f3f835fb82902c5f0e97e51274425b35e9e328bfae138c80;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4363e16b7ea9ebff12873ce64899676db6a667495023b808e9e905d46bf461da5b2dda6487ac876284d59d5bc2529074f5e4b8c87bc972d829217c80ca7ead8a8a0e2d2e5a17883ede21c088ad2094e507621b5636e50d60f4a506e34b1abb1bbe8fb4cbcd6f1e78ec159d1a14531d4a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80a9196ad1f7cf1b728fbdc3ac57894e2aa170d2149fd58c9523bc942d66addfdca2b404ce846ac4afc4d258ccfb9b43c3d1e44b16aed7368edffa845eab49072383a946011e46703a6ca412e635cfe86606524d1aeb338621225adf92c8b3140cf37ff4117dc40456871b6934891fbfc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e9585a298826d70e17301b75d37c5af3923df8b7f8ed3ffcd787ae338c3838da61edde915b48f04b8c7ebb98e943ca294f5e89fa95fd07e98abc73c0820d1436792b9cc2e86b7180c40f82bf2cc527af7b7d286068d3c4f09dc210bd359a001d302ecff8b7e43fa0467aeb692afd8d5f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92b7b927af631f2a158790fa8b6d725f1c04034ec2b4b74e13b5d79ed81b964d25159cfeca688bcb815662f9d1b956eba637b7c5ff421e8363e9f6bf5b02a2378b289471f682afb5982c35fa6f28344300dc741c679807a096e96c93921c11e73ea7fd8eda6e5cf5afdb4ea5f359c3efc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he93373a4a163f47559135862da440477491e135a7487b31ac4875bf101694d8e51cd2936602869193e5bba44bb581b39131243a995ea2f1a4c03dac0180acc9bd63111e826d242983b5725b919111be0610cecb5e3f3bd8d0c7a6d328c0e895e0b73090c4289d7e643026fd5859bb753a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30d50a99b4088b5eeac7a6221afaa5f08f5751a8dd5887a8e6181af54e8ef760459dcbc644263054ab9720f5bc5123e1c7f46647a59946b7bc675845d957e639ab7bfba628b2dd2976bdd5ea635198bd5c22c7a918c3f163430f31adb9fa8bc39d71d845a2877af35ea8bc448698531f9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a00b6fb6b180cf894555ff6f2b43f89847e8462db227cb5ea27995f0c0817bee0e6844c38a819d5cc344ac7f1082a5f01be33c244fd439e048c8c1f7941e3f1031217882f2100d97d7ce7b77842b81e8aa4c04dfec22fb8ac549fd7b6b6e57611d5c686a90d6c86e9b2b78568f23e59e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fae5a4e37c6df19e725348a410f2f05e607136ddc752e4449d83a7e07f54504494489301325b4dcd6c9690d99af60f0c3272d449b90a560025ebba1caa8f94a26bc93a712a4fe3ca49ea8d2492a9dc61fca33151418790772e32602a4bee0b67b1723e98101eca65ccc22e6166c0ef5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ec7437bac923af8a3216355a0b7013487b9b75c7d8dfee8a481e8acb6d50cdc660ddce33b505185364a459fc01263f5debec5a0cc3cbe9f6f7891bdcf07be0ac0f2756abd995823b73db4462cab357f8b9e6b526f3f635b2934a195bd144763c9d52e745c724126ec60f167cdf79cfdf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4fd830148857d01c6474d63c72e56d22486bf141f395459a0f805cd7258ec179ba016f2c7b00870338490945d2e37d1bf82c5515e7f5309cdc0ddfa2733b2121ce496f2a48bfa241f003a0a813a7a2af118ccccac2a489bfb58256eff2cc879810f4d8b54cc3e06033a9189b1382e58b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae1dea8325fa6a1a82e6ead9a49485227aa27dd7455e6bd2bc836aa19a857ed2804fa471daec82a21828353668a02dc0a9b1e03832e096117b9e2074bb7d59dfedbe44ae30742c966d386d1b7a55179c2aefad45446a176ccd89e45f52c96f3580329239d577207eceff589854dd5b1eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h506d1619183e606a394103221782ddbd494f75310a5b319235ab3348e540c9059b072ad6dc9561d77a61e1ec26189c810151272365e5b497d2131f3e4d84349c8f637b4e485bf7ed38e6ac54067a4104cb87daf3f0eb9c92ac9dc1e9328b00f12e26c222244a702f952e97fd5e72a5c38;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedc2e852390c686511248b4e0a63c35d12b1ead66b3baea3f7282c54ca270005e23787df4521f282f0f0910b1c2dac278463d23375b0510858438c14c4a294473f55148e71ad6337e1457d59e2cceea22f19cfe3a653ddfd2df123f5c08a7612362dc7edc1637faafb432a566f5211bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heee474e0b16cce200ec69465288902df258354ae2c7eefb2f92ec6e9667fa36c709b82908a292a0fd01ddd22f5eb5293fc8214eb4626ac18eaea7530e8873974705b71e49354c80568a2ccc785e80d9ab6c400e6692806032847cea1bc3c979c97790ce77bdbf10b96f7f75d0c0a3f098;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heccc1a413e3d00c297a2f25a409079cb5d8c0c4185cff848b9dcad39ac439b6e345510f9692ad156413f142dc61ecf1819331255665feab2f7e8ff7c1cfb4993843e64885e540874db823cee8ce3584653abde65c00c2dfc12903edc59bbe58d4798ea608194e8336a366b2199e5796ce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc89b2a7929a3ebacf2211972b77bb6e504fb9b0ba7f37a46765d692ae712b0c567bbcf6738ed36b2e3bc94f7db1354d82ac20c50b9aa33a09a609bde7944c3457426cb0aa6a86dc1b8514c7283bb419d937a14a406ffc4f6e730f1e87ad71d5f6083b65c42f8d4c1d26518b5911dcef61;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb798e1e14ecbe39b4ab20d304795f870927d354df18ab9e8744f56cc3460e198d2f0b2a972f07da51decb542db3a7eb55bf7f314318baa4a7f0b3ea1fae3a685347396192acc23a66ede1c4cf94f73370d521c3d350894a6cfa24ac2831fbbd3c91797ac51e6d095a5824f0828d0c37d8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h573ba659dd62eed360421e5819708085c3e78558e23021c6b33d39e1681788c4d64649f265cbc35353ab8274d632c46887da0ea11edcb75ec654741a00c47b25f4ee0df1e40083793fe879eb3a515f21454bef43e0945b13664b6d5d1557fa2f5105e5b4722016a160955fc9f090cef40;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72a3403fe7cbcfb3b6cfd968f736968abf176bdca861d69a594e9c4afe027d0c9948931e960fbdbc51cd0427767fec47628c8af4510d4d9f80b382257c73ea730f37ff4e2464cf13909c80cde772182878e94c8085b5a9f68386bdd89402b5a79974515b34820763d2010ca73822d9e9a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf73b70c1c1d9bbfb96eadd5ad41a53afeaa0b1b659b4cc7c1eebaee55d3c05cdd86f42cbdb6e31095f7d5db211b8c792b5882a18938f6b04aabf1fbfa3f69b15a72a55c51e711f0c4b9cc150facdbc0bdacdb067b9ba4a742182748b8d3aed223cfa215b5a8f1c2fc1de349108eb8665;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1589bd9d20a1cb943183df4934d0b203b10532145dd070257d0aa573d7e8499d98ce016e9a6c20fe6cd464fb767ff659fcffab8c26d1054229db49c8d59f479967ebb82412cb4eac1d6763aa0f7011a46ac5c041c832f7934a14e110f6b421aa655f1c491343070e7f50f324bf6f12a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5bcb2d679fce16f56d81a46fa7d7b3be765223a99df0d474a3c4bd6e940988b27ac00eb703a6be4c4d4fae2c2c5399db5d1d37da65958019d98e87288ac395633e28399cf9df4a2675dbf891f372fb5dc3bf68b21cee2276d9d35a5b89135d898bb49b5a29b243ebd7e92449030b7c473;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3edb8d2851fe38143f9288f9b9ab817b04d33aa1371eeb2390e8cde0576c81c519db2818ffce8b9d2fc56410497276ae872a26ccf6e46cd5e372d64d0b904cf8ee76e433fa534cf1bf2e5ea0e64e7026edb4cb377ff0c2ab8862ab6b4adccb91887aeb238ace50317d7fc40def13c172;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76ea4ffe71ca98b0cad221045e2a7a0f2581d3a20f588e011650a7a79a96291427a47cf25271755bc2734f86e21f3dfc9fc159995b44c637c39e81620a79f09004e530ccd1e948eb0484e1f010f3c3cf41084f1eb654af3c2272d2bce2c3d3c6cd8312c2eca77c367a99504ba38d125a7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57d6d8fe96ad7eb4285a79b0f8051576388c466d4b882d2e3f89bd84f9c80b919285c094958ec0e671960c7a75fb5d57d0ed903b2c6cc54b6b6f96adac26b06a104ef3c95abc6eaede64a9e898371f3b1f41383a3fd9e49c956633edc760427a8d894d09917a905a295292cc8865a3bc1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13d3e6c34c4981cef5691860e0884b009096b8170e93462e0f8aa87cd6ef8c1191e95b7bfe6f46686d8555e0b304d13db22fb72b80a013499f365b18a4b2ef2b1ece432624b49752bda8aac46e96722d8b65805e7069c0bb07e28f50bcf89673a7470ff41fa752502aa3af14a7ee14cc8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hea4f11f5c5ebef71e1e3666345c4e43df707d4991934c11e73f811e60a4ca10a941ec376cb0e17313868677d2baa844cac8a95e387479ce8c5028cb00ef402d6ffcf40dbfd6707bb6594833e0e80afcd1df128445d364d75c2b65f503d9d14e183725d6d94eb43f36d6b11c2271ca4aa1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d75e29cc3dfaae1a9ddcb9143287afa84dfcbe8f976aa2ac51cd3d0d6e9b7fea75e19ffaa11e8561c6659b16ddf6a2bbcdf0c14b7baf0f4d9d0c661896af3a1991100c849cffc99ffdfb28106d0f3ed9c78c82fbb60dc93298324885bd421131dc869420445687d7ceb2fecb3854b60f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59df39ba69863336d9f9705653bc27cb93ba58f4d3c7607fbd0036a65eddd2636e921cd6a8b4fa717c332b560e14b28c748788e60b699d8f7d940f7f2dcada985ea652e43a09014d0d7c32ee05598cf42b1c331a23023edfb435c2273ccd8144584f6759c24e4002f3da645f74af0af30;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f331fbc49832de7af06be81f449e6585b514bab3d2a3356f751b3061a44dc2c6dd7a605c80b04ef4b3e2a6a8b3865be6d9a6f9edbdc1de99ec90f53fa290b183bf80db3780a3aff1c0a6f246344f613a19e5b8b8384f0af7030fea9ffa76048f27fea2727c2b03d8fb695861cbed4638;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1a6eddb465415ee6724c254610dce0efa7c660e0cd1f7c8f9824e84c442db383765b529c350847d92e20bdf6c93e41bd846c7ede5d9d3a33e53c0052d406224c50b1f5f21cf5413adf689fa79194d192c68f7a694830024898d48a921584cc97c0e9af231e78e663524a6ef577c063e8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27e2d95a211872c8372f049e53a69ce1750a5ee1d2824fb4e9d81706e9cd58fdb9c2377fd69451cdee61345c9af39a6f6878d7e5ce8614f75419946c23b21dc3eba95cc69e707b4670617965b78e58f20fb6c58b1ddee7f78686e30db6ad7977e58395be061a4f9107068d62ffa2b7f78;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h622ba64166c67fbc5352f27af33e8a50b8a2ea366fbd84259c99823221c53029b37d5433682ac8ecc44830b807257b69f79ec9c0b3ddece63bb056ef7ca6c707027ac9df8ee1836c1d12cfa0e34e819dea459fef0ef705b2025e1c904ac50be6cd1db993b69e14e95296d221ff2d4512c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h446ba9015b6f61c6e93c0984fae36f332158f7b5b650e03193c3c650a8b396b32e73b923cdbaa8927742199765805c24b1b27130849a73625ca7dc733761d3529427ecb1ddcb0113ffac2c5d513eef5a34f5c53826e2f044b8bc0f6857ccbb35c4dab1fe842fd09586852c2dc4a939c1f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha614cab73fa0dabe29a416e8ea6907cad9836a0a18452698e8cfc104b24146b3ac1101c7a33ef114ea7def529ea8da1e2298457d0835ae403342b9764973e5fb9fd2f4257826b9903a46db3498608511265843a1f472f25e69039818484f87d0d8448ec4c8cd96f6c158c2835883ca328;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef6974ed55ec1bdf81e725a95517a37e5ca164ab5f1214cff73c3e9975b54236577f6a5e4da02c1b0fab2dd72395217f57ecf3321a03a7de32ec418fb11ca56d5f1173fc53cc3410f3bf8e5d100f8d758350aa1e7c7c3ce139483007bc99c1b7c22ede462cdf590c15e7117d9332ef427;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2f52fd1a0cafc91a5d50f65d23f1a9d2f4ac663a1a631d897966e7059f1be8e9ad8bdcb726d52d6eeae33ad64f33c54c0f70f314ab538ef70db05a5492adcca1a92135db408916e05dafcd524fbb700007f7edc096c6498376cc22254c37b632fcb80b82017ae77f21fe389598b7c701;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha05a9746bf2d707764797b771bbe7f2d0de4df1382211123135301d5415da5a15f4b7b76078cd977ac626d22323d1ead8f1fb1fb4ecfc28a4640af0503f4c8fad3c71d37a53dfb729612a204f111cd506161ec4aacec725b232b61a8841766b250b68b5b73742aa1315611291c3ab2158;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc0d5590cf1b16d628d24ea9fea32f61767d118fe3a11921b12b3c758b3ab93596f03c9f8b72f8ef2bc8377f95244c438ba919681e6ed9ef692869bd2344bb2ee0078d3909050494046c1448ea83c0e2b09c39ce1306deacda73f9aada3655ba44e8a041bee78d3892a564c3482d973108;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f0b2fa91b5f20a3bbf21ce8eafeea46c532ae40faa896081edcc0973145d4420ed01b6021f6043cc525913ecd42143cf24472a9bde4afbd45de64c74d60fa43820dc6d480f312b74fd5859e03ed46be6dee4fdeacf405c10d6ce9fd030a6d5ccb0b4a627c1864dad50ec978e7e6aee68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hefa4a8d5b0df96ef91f0c25f732ec71a80f516ab12903ec17b3e49af47c46f34629ef568e5dd61e530980f053e3a3d39367b7aa5a167e02875118c847d946a06a8b9db85f2b57f03f414a36db34cd810bed00a62d52c334b46e77c144453190c90306e4b9edcfaec79ee22ef98a0981fb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2da717cbbf231451ca535f8e27d4ec1803c6c793ce6fef88eb52d93521169f1f7d75637093ae105d73d8843f3d51aa75f50c72f430d5b2674a451548ef2f1604451a01c127c4ea7433b2087e2aed844126feaa290097b9e72c92ac65515be93ef883258d29cdb183d30892036619c5635;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7817348ca7f4b50e742d67d7953c14fe9177f5828cdcefe84fa66105e438622760b141717c350656d53685c90617e292200a7c1039b16f0979927a20e259522c0dcf1bee12146f16b2b84a774d0487f5e5b0f91c90000b5d636aae4e2ff28fa69ae79d8cbf873952a193bd0e4031ca43;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4aa431c4a5616c598a67941d14252a0dd57bc08bc6111ab5449d7e4def3efe7b64254b8c5c231d9a2c9ae11f5505fc68a8657a444acdc005e6a1448342c81bd55429faade3e848efb4195596b020115095d1782ba4c9580f2082f966f91bf189d91589f9ed992e8a79328b2924f579fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd695c4df8d024fdd39e4fd14623041b9578403adacdf549b59f7e06678c95670e7b3704d272f4a2480350d5ac7dde1bd7a85850237617bd6a3e84ce4611e4e6ec2daff8541942b039f9379521628beeaec24160b3e944068e10914e3481c9bec9fffd45c72463dfd0a1573e2fea005ddf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93018b6eea8cf704b0e960a7169c58d610d0b6b6ee1bbdd4ca0110c8142d50db3b1aea7e199d32e592e5ebb8130955e5ddea7397d23d2ce386792062e040a508af2d2774b959eee8b36226e26acb84881b6a0eeb0250f1e02cf7d43139bf2aaffb90388b8d9c8430e57a95dd72a88eb1c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he411b45f5feae834cd7bc50f0123684f4bdcc42c8692ae24c71efbd583783e2cebc57677c078ab077167bfcf8b0d135cab398f2fdb86668ac036e4682493f0f517ea60a1955a99149aaed8635e88446d66e9132b93f810850b086510b2a69152c302e192b29953369aebf01b78a93f46c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58699aefedb3768f3b614cc4c6332dbfc7ec1512f8195cea1e458a0883adc13f2b678f581125e90fe349c04e04163a95af431f655cf935071b12bdf16258651022e71913b3b019c0ae237b6c665a55df134e6ad245957adf725f5ab1117c451a2ccc3183c045d8d90236186372a91a83c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27f4efcdc2baaaae6fd3ccc96a14f289fb2eabe2a5e1be440221f5093560c19e93a461a9eb8f9501510ca26b1fd3b37472a9eca8d2c6fb57212ba6db0071bdb376257d1142a91539214d9b6c4fb65c1e2e95c8d917633e2bf82fa14efcadf6dbd9b48b1733505917e0d0a12c2cf9c9892;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ab8febb9ccfd109e03039cf5319b953bb2fb7e1bc600b49c61590ecd4481a5225a6813461f4786431aaef55e8272b08871a1c32eba9a28a5435ff63a07a20f09cc118d07a3df9d7183f657422cd40ada3724ec32e9536834eb831a7c10e12056d5fb598496b3c2cf01ebb3146ce880cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d0df29994e81dc188cfe6d277158fa0d03814bd25b62568b2ea1393760a46384910fb785941de9267db93528412ffde603beda6fa60af602e975501f8abfb816a67a10a6d114a1fcafd0481df5723fd2d724e10217b15fa1794e2ee881a0881bd598e73c2af299d6b848bfdd44ef0b6e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h407df2b7be80a657d1dc8d98ad360e4ea2ce7390d452da8234abcc535a91649bc850849da3ff066d5918b7de9c04d052d7fecfe17e215de834ddd291aeee27f66c993393b59decc886563fb9813a786fa2fd18c1261e12d4d06797aa03f303d1b0e5bf41615918e064d8e2714f9743f2a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf95cd082cc697840d19acdc4d8e3289f435c6414f86bab3c6c64c3243d485fd7bbcdb65f52b10363d0b89ac705a41664c9dd4c3bdfe752378d1eaf358feb7643ae0cf64793711e22cc6a38c564966b3942c8ca1d4774bdb6bbcdfab1ae0dcdcbb977d94705d8337c4e65a130523fb2dc8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43c103e789e2f68128de918b69ab720cc153c86ecc9a0b9726e0c1253bbc4ca6c64a59141efc34b950c6f9fd634f0bf30ec025c841664811cb714cff76752ae7be1a0528ea6894c1a6262d326f90df36d06d4fed9fa3e7c94a68542cce8e6a496a69c183d3db553fa16bc426240362239;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h941413185b3390e96b4567238c6852d9cc2a6d5028490efa3850a8f34cf4d5f0a1f83f43de64018b2d79f92ca2ba170380cf6f86f885eb55001346f3a07a44ed9e3eb5355561249bd9eafe4ab1e5bd18c21b98e2b09addcf507eeeb71a66b72d38985d43bd84a480dc00c93a18f1633e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce7a06a6c10bb719e9097e8be51bf62d2846455886f23cb424962cdf62c0dde5476a9b9d9e845cbb8f3c53485430d1c3d59ee3776bdd2d4ca34355dc3285fee2372fdeb41714607ff3e9bea6b2b6a4a5424fcb439e0100927f35b3cbad4407fd2ea481948a732f7767041b5f19a4ec0c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3be1f2d4901dd6e72b700ffb961ef305a06b52c7df0bafba087709f8b1c82067d05b1a4515be8a24bb637e4076b521bcb1b82a63854fb937b1ace15310671f825ed01387015f61313293dd40b139d8e8a6f7f1661ad89d28675a0b7d38d6fcda059e8a34b74816a8ef868c93dd769ecdd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf893c9b530e03732ca78f175f0b42f4056a92756210e2b822cab69a2d17a2a231861e85381f7fa156e9330a6b507df54d09a3a4849e11cb8447e3595d41a2f536e9692e22353b11973ae6706cf92cdc95a322c7dc660245aa7c1178b12e30be611c2cd6b5b71a4136731505c2fbf311c7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9608a66298e5786efd68ff92901e760119ea6d75eaabdc8cb37bb270f0663430b69fce8e21966b1f915a51d7cc975661a24a768751a800880933b86d420d01284f5d23b447616f9082669d441580bbac43bbc32ff7006862e61d18eb1a5b434a57816c4cc8aa7eedfc842f2c00fba1b6d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38160af2c6d3bd105623a75fca601e37cb3f22d154f206118b3f77beb8ab01d99b8c92f708000db42de722d9dc56758ac10beb6416b48c90a607b6d0b610887bd8d679edec13f85b29d0b149a430c0372d66fd73b968bb63693f56f551edcd7ed9759fb2a4f4d75527e4fcc718991ef45;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff38303048d30c3b31dac663f9dce0a190ea943a64beb076a41444f8250684bd8c25e684204d19aa0fa1038d7109f385664af71f53350805dcf11099b6230561d83de5bdfa2fc2916f8ffe8199922d4096c96397358191dfe2ea4baac9d5f5e1cfcf50dc73a4633fd7b4bb3f0b76dbc5b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb83e04a87f2df64ef2f13b866a50351f2eef781d3e8d6fadaab7f10c2418aea8d71af7b3e40af9d4ae1705f815c760e1129801d404b559fc3e81001558549f46e3de7ed83fb0235196c8ec189aee022d709f9690b23f8daa1fb95fbc29c1c9d320bcd97b6a0110a1641f03e8d3dbd40ab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9337ca729a23bf317865c11283e82679c67d8577d507d47a498ab990b4dcd0b11f75f74c115df9d42ac2e46db71df5bb3e07afd4ee0c00fc7ba7269dc9ab3d8e2fa4d86444ac6361558586d665c7f5df3dfe0cc43c8b49c367faef8c81c0cae64be2937609f9ba1a6540cd6e5e7ca7f8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86072f17ec4a815109211b412fff68ab37c8d16a38f6e005526cb96fc443a1e0f6ce3e8cc05668206d604ba378d112a552c629b447303b4f9bb445646276e70c141b7165548d2f55d4bd3ad042452ea5ddff37cb10857de21c621b8b968cbd7a51366218269141f19d6f2adc56a2e85b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4a6fde395b7d16f142fe0338cee72dcd08b21f1b7fc5446a13a55350709c4b006cdf3a9d999574cad440039e79102549b47b03a2296e014b12a1ac11c1f1f683162e4aaf47439aa27d0ea3dbabd938b210cd0841a965b4d326fcd3ba3aa54d83d295444e44aad34affe04f149af49bc9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd049c2f45acf0bb860e10a604963c3a7fe36923b56424e4d8c8cd22b8fa1c304f7601e22856c8dacc52a5d600f711773e504a56a264976e720bd32bac118b97a8641647fb7823717d6564431abcdf692f7d12b61448afd91fb5a44a6680fa9361fe3c75b55973dfb743bdf0632aa8c6bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab6309debcca318134cec6a0d727d73d42ed6655d5a076a8c93f7b81a3d8e913baece862b9ef7ca20280998f32f6d931b8ef3c48d48a1a50d2f78249342455b472726e19dea4d3ec981739208d24e0ffde35459df513e274c34f7f05be3aa44430189fe5ba2bff256bb92aa5831c42b0c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42cc7354001b939a8ef38992c40b1bef547794751b7432e5755f623e3ea6d621759f41192f24cc0ff21ff0ea0c4c338f0ffa2724adbc68599bd90f68839621c65537f1e5fd96891c2d7612bff9eddb461a9a04efe2f52def29f2e8a80cc64b75992ffa22bfe1eedf0b6a64a62904fdce4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63f46f73e0f5ff82f28ec4c8ce582d87aad9d0eb9b7a458bb4d2d7bd2a72858b89156a04578eabc54c5850bbb5269703aa3b653cac7498b59a10ec2b6d6c638d97e2b23dfa7bda8cccd1a43c72ab70f77bb470506daad4b6d3e16e6f8d26bc286aac04792bab969e893a2cbd54fb632db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7517fc193b6b0a150eba9126b70fa8911a8201b5cdce27d9ee39e0d40784a611674bd157114e600e9429566886d7e0e2dcbd94ac4dc7aae75a5fb361dcf5e45f27c58ced6f6c55c6c7108fa374090599bfc9b06a689c559002daa2357ce3dbcbd8d0e0e6946a5bd1e73bd31482fab038;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54e76f4b58a5fcc53149aa6dfd404b673f2e9bc66cf51c6ad218a9ac21f4f1d60eb009b4fdd29938de1a1e91b9d4841530112ac7db0fef562001d330045c203290f5fa7696c2d2925610c84daf59855893976fb306418896daa9ba48ea67ba0260ca9b23b43b995d374abea7722a01013;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b1383430905d7745b43a957e4d395afae27c933e1a56119c647ff8dede4571e35e024b39e761f26aa5c71eaddf1fc2b498378766d5de6143793716bb7005185206332c3fbff08c0e010d89112677b8a419d908c5b8525e31244619f26fa415d09dd4eca8d45faf1da476975f5decc83b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfd62b3f23bf3d7e599d34a7b606885292476688fb73a89358d53240f1a9c2673085fce2854807870b94ba800bbaa1f94fbb405a2d09da4f500efc94298dea4e430e74bc04612910e4e3c465addd539dfa2bc27f8fa35241f6a9101a2cf92c33873dcf9a606b9e2c278b7ebcac960781;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf393e86018db2151221508bbd38db850aa14096c62e55ec928bd8972d8ad20103433f7e911463f11cfb039543f77d44cc838eced4c19ef2ba7bd2802c76e961e09a24814efcba582036ecc2659b494dd2af838dc7f91d0e2be43d9c1eb78e7d2918a2e7cdc5345bb794db3ea9d85095a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b471f2b2a523f4b1c08299133ca6e3239b012cc40a90571d87ab8880f7bf99c050d1d32969f714444aad394a744d98e05a29de13389a557decd6722db82f85c49d14167322015f54a2716c7c2a00bc99bfd85e2f27fef38e5185cee2995ea0fdb0e41b1d001b4bc7dfa4f895eda468e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8a7f9c4d40d425673132955b830ce68da9c1f62f0d5ff9b4bfc172552a76d7b7d75581bbd90eb176f473ca66c7475a9529844439daa0dd8e85c148c3df93ece75b2de56d0e00aeeb411b90c50d783f58016e8da1ee131981811ffdfec4142562af0d053fb4aa327b2854a22c41e9a5b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9c01d556ec36d90ac02901545e2dc33fe0bbdbfc0f9b08c9d1848040abffad40e2faf3c5b8527720b2811d497b6bad0ebe4c974767e25a817aa85c8ad6771ccfb9d8e0a672ff16593b2f96cc17d350d9d2f64b4576cb648bfbc956ae96fd4f554fe0b220e38dced56b399fef5358101c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf93ddac9f663987f512a771ed28a7552f5dbda711424245854275d9769d4da5afa0f3f883097e40ebf7648a659e92bf55f0947b21e5576656152fc2027204076c3207e76f3bf59714625392ce7543f166d94342446db5a8f9be7febad41f11dd45a3993d8c68c154bd9c4a69c914dbcd7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h880550f3944fa673b9b5a5037827c74f0d9cbc148789d1df5e3e6da5dac98db501bb8c0a28b39b8dfe3a012ae83c0265bb23b78f69292e7f268f7d1c9c24c24c763e6c70b9addb04ba36336613cac783e7726d8a88a65ec1cdf238b7040c3cb6c6d96543cac4eb4c6bd6daa3721174347;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30cc40991793b2f8f211b7fa2dc558b7fb9d4167c1f22df6bd8948a418b8918e2817b618b05392a357580ea61288bc0be57bf5523626a35462dc4f352498a6b6975e7488194c9324ed828f16f6e8f4cc4be9901d67f9aa8fdc30934224832afd6c331cfabe40c6bf5468414c0b6321ac7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d1d1087515dda118e31e649287184ae2c89f55532917aa3431e8feeac16406d5fbbb9be48411367d4401307068e4848e5683a7f317a5834b21dd52899caa2811670d6a8fcc38eba78a08b7ff9479bd4f8091aedbb342da6be1bb5cc11a0ed272d7a045a37ed8fa0727cc541c27e80b18;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha42335a2ba63a534f9561354f5c071fcf05b3e7cb0ce4f167c521037fe2f0eae4b7258bfe72e85926cddd8255e4e2ffcbbce64e9ebcd2bb3553cee2123db65dc28048ac60bfe5d338d4018ef5bc876481299d51b9421229185c80faed7c163d62a6a579a0c6ddfef6d31c16b79217b164;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha734a05690f4bbb21a85b7ae5f864235f7d30d0444b614c20d58f0a5b9711ef38d9603fd195929ef0851ec460d1e6c945eb4113b8f05d2c191a5241133e3cb64df8e1d6058f08c15d2d653ff969162c9d2ddc3b3016762aaae46acc08a8cad18ea33bcd5c6108dbc562b7b06a45bdbfd2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f3c4f54177119bd563a44a569844098a27fa8b2e85b2718d1c6fe0d3a0b1452024e8b49741cbe3d977f928a5fe5e8e6d6433a2aedb6c4f4c9063349d891f49d366b64973563f63ec861945f46002edfc540229c621daba80b3bc4284f6fb3e37678d9a49babe8d658bbeda05356aa613;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha66fbb8e51bcbd8d725fe16bd75c17694fc12711884049b6758ba244853b489a4529b9d817d0860968bb7780bdce85e2c957aa41401a6ebbc32a6a7006e4dfe15f1018a9773af3bc9d2167bfdbce9685423116c3b1c3501a810d9b66fd9205460ac18ef4772cf7ca2d3be9164f1c725e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb7fbf7c4cbf9f4c4a93e31dc25c3568d7a63cca1bc830fe29103506a1dfd5550669d22937a02da91c92e8c12687184543f183dc122e71277842f3030ab6b333b4b03f7806d5af75d8622aa053e81babe6f4620bb124ade7a893007b6b6848c66e56b52be7622765dc3b604ce9c98f753;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d52aaeb3c7c17b571c5d376385448cca6b983484a92faa9603afa7829f82e9261993742771e4418a43d8e214ed07eeaa45c7a38b4d2464e564cae0010c5290cf2509bb416bc201811d99b990a7a022e08f53e8ae933bc285d56379722d8e3d8035670297d0e727a95479360d4a313ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha157775ac626b0d6a3c3452bd956e18b23db471db82710fcb93f9eaf1a1104d093d34881e47011fd2d0b7a14a86a32b887e6f2d31034b1730b0a365264c0abc2b1c562b95ada1c75039cd85a2f0ec836efb4f060dc2b4dd78ad78a50b311c86c946ae17ab9e7b551c2d3f9b5b09594d63;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ca53aa2392b408cdeffda6220cf88fb33681a8de92e190481d15fc84adfea3cab0332a2089f9ce0db3558155ef767b5c8ad4dee3af094be8ac5fd1ebf1207d3e67923e56c998bd51eb3420960431f58c43cacae34fcc7d6863db3cc2ebf6ece3e4a986be0f8eef2931e321654b74b18;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he22b88a428879c3f02d7622a145379c6a2424fe064092220f69b2f63e16fc3e83ba103acf1fa7bea404c3c6fa95863d94facdd7c012ca8114c4b8d5bea984f3916b332ebca3625e55cfe8587efa6d7e3e6e099c413ddbf8b19f9a0ad32715a1835fb4838bfc62c36afafa20a2141ad74e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3057ceb23ae251c1983e9c2255166c7db6dc78d61e708113a2f636e44bb8a8c6dbf555e8bdea39a37c31277ab0e49f4e5d4f28af552d1ff08d04f63ff50a246e9beaf0ebe087cdd4db1c7f205e5799ada6016febd7719ef9ce7dd0439dffc150c319b863e2b6c8c8ccf5b544b97532ac2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33b99b9aa41d029f37235ce5dbab8e2d2326a542c31ad90cc479d8523da58817677b2fac0355f078dd21846667106401c6f6af7199a6040f338a74aca7c35fd447f9fb288a546ccb181fe5eba0c73b2f101e6be80b9eabe66bf2c18683571734df617cf8a82ed9bf3c6fa92b685e4f03a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4ac3654c06b0ffd3541e6d12d6b6490e62199e0990982f73a86e3434a181f848bcc774789db2ec12ade2116b884a1af99c15112d373222f7fc13c35cc2e821a767a33bbc572abbc53fb49d5aa59f23b097c0c746f8a7053dfcac054ef997cec9ebc95166ac4dbbd820074535eee3c792;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc50a453b494a0568f36048555ce7da6d3c351e08ea449767df07b53634bcd6c960e4517c5a019c1d2779b2a4d97a1aec38db1fc0e8bd79e06529a3401f0269b93dfb8d789e96f9a5a8d9a21647d91b1826712ca6ad21c11f5dab7b7ebfc4becf7840e5f3b1409d87a0bd0fe7349f06984;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11aabecb04f1bc6b299ca666ddf39b83b3e094d11fd9d18cb518cfb9c5e578c84e1aa1907ae8a40089cc552c4d8b8111b5508baf54fd6f01b1370e0e65cf92816e367a020e971c7c639ee84e12e9c066e24418fec8bdaa7a3c7d0c6bfe72e5365e150907cf40459649ca753b3394b3ad8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3150491169a18d41cc3a9c118b3d870374804b339bc69f293ce5ac78c3ce8153f68d88aa8e4854d7fe0da4dcfb48a3692b70e7a0e14ee057845210cd845dbbfbe597036c35c9b0e3fd6bf7a1b37d1ee9ed861e45c9faad51d57cb53b3713ffa87fa4a9a0ef3204c42dd244c258f0ca57;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43387afa8242a0a824cc290af7ef43886a0269a3aa6178e0636f08b6d8fea8adb14e84a7c2158c113458ba6e1af50feac7502404c45eee22d5cfacc80985a0564b91d882bd5e59e5ad7c3476e16abb494e3f86c01952381858cb100c0b252a86aa0a8b72b6b9583250988bf9b9bc75992;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h396fdcf6f66c3d6cdfbc717726d9aa4ad811f104b8b47a0a599ae6bc3251d88fb85bd49d98b45c3a0c602548e4721a591f7d4b7bcaf4d26604dbb4aaaab6bb4a47c9b34d65c878b21046e379bea12319bfa16be620d3721aa15c2959bb30a1326bc3c6f325ef861fb3b8444feb76ed2d2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h566266757d6c51fcf124d147c7ea056a02bdade0ce281e03292c11222df343f24810e0e3be95aeb2f59c850a6d642ef0e1d519ea926b39dcb14dd08f6cc69e3d07c4e05c73cca219cd3a06ba13ef41063427cc7c2294b601795f411447ce206bb01432c231b20268d557d0d0faf05039b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36430a82d7fee55092138b20d897049cdb3815b6a0ad1d545eaa754dd4c9a574fc209a0209ac1517474830f7bd73956aa41eca44a1ca5af316633dcd36ea6e8105592296ad7273a2aa9c87888a7ef8d39e49754928e27f469df33f22e97d086c54fb9b6720c036a18ed38c5a9a2c8db03;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb230c8775f619ef33b5c113b2b4670a543c8c5fa5ae753e244bdcbb25e4188ffa6a2d325db1dc0a235d4a33fe065977a80b6d54c0389e30d9a8210233beab53403f63d971b716d17833570d5e55771d94a513432ac18fc421f8b4e8c1deb6b6ec447bb0b11e3e1b644eedf5c133bfbbf3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a02a6a5baf70773cb98bfe87eed2bd3b5fec0c307464c1c5a95cface295b3e178191476d85d9f3caa97105e192f15f6d99feb7558edfb78c858a66d4b9a2ae7b28360155759053b67fb1378c47b31ede2c8424e361cf25ed497c534b5bbf9fec91661d8583328684528ee6c12b8eb16c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb78681793d66c5dbf23bb4095899af90ccc80c242fd70c45322859537f969b498e387e941c24deccfc20976257fc843f239548d9593727f0b3a2985345e1e3e1026992b7dbed84317d0754919066ad52b35a114ea3a084d3aa1e39af8e53e2f297f1d8a9d0f7917258d0f9f9aa2a1b16d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ba65d3a84afa461f05d6d800846d48a481cd3c2255d0776869dc6be8bdfbd2efa1250e504c750970ad535c50d1743f0044f856f85a58753e977932052cae5a283b7f548225e0a08fbef0b5ab68035fefce61fd5cfa4e0b089dddb9fb0be56847fb0bb379bce9fa7cf4c9c9fd66f8a4a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42c781771c58769d5720d3ec0b01ada5bbf2745e10db799faeed9c6f4e63c67f4da260e972b8783366219c72217a80fb3594dcbba5a157ef5b9ce42c045dcbc85569f7c5fc86be9ce3d34e18c19c04bbfd1fc84b4f5c4dcbf8a16a76f2548b2df2ddec0029fd4d97b977021e94119239f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b59652c3405c11f070850388ea851f1effb3b9107fdab92ef1a00b6134ba9fd96cf9d738270c2b1361480c6ca909aa98467ccc9c5b165878c46ec026b6076c764b9669adab15187c83916a3c41f10b5c06cc9de3da7779f2373d524b41eeda91e2317f68482eee2a807be2aaf653750;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1285d6b6fe052b288762173dc7e24840055ee82b1a847c179f64f7be537bf032df25ca8c53b54c26fd92eafc3208db070363934b6f4600c69d12901ddf4fd717701e5d4c68084e71fe2a7d2b3b200f1c3ea10dbda638d85f1f0f799e16de3b809df63f79505680eb23b71d0e2014c236d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec662616acaa59b7cc981222804d6317d2afc3d5ae7bfd555f21660ed67aadef7fa8356b9c26005f11f0c610f84ba91c20d8523d79dcaa6b7ca2b9e8bdcbeb1cda1401098accf280c4071ac166f18b69698448a2a1c1ad13f3bad94290ba5f26a63966cc683351aeec7135d7b519f4f30;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h501f75d65aa05792d745436361870b0243f2e2110b51454917c2490a7c6d9639cdbba6c11a8fe63475053f77eb5b45f4a2b02c882c35ec50b936128fa30258257e6b82f4c04e5df41231d49ecb5c205127e8b70418fc396de6f3953a9fb4b595c27bc2627e00a5c498cc77cb29323cec0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7656fb516e05ea65bd4534bed0f8ccc1db3f38b613361689585fb7e93b0624d756a6a4430a33e8c3c4ff46f5e87392f424fecb3e97bca1ad89e542fb912f1cb3910f1eb09473e674365c9571fbafbada52608591b7e351d15f934c148a0c0fe6589447b83db26938970f1030a5b0e0760;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h223bc3c554bc56ce289ca4d94014070d4e4329302c350a1c518873f80ac34180ec4312e9e238810cce4d7b5f839279ca278d1dd20fba2903530cfc25af5679fbe9f9ef74611d237e81bc9e1e20646758f0ee67a9bcaa46c7566d18d18a7c81e15843b1ce9017cdcc23027745d8ec03d2e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46de741847f134c826ad886ff3188e065710e70ddfd382ea562515d126dac5767ea0162baff24842f20cc0b8b021549f182a14ff053195cb7e6d7eec59d5ae6a65786b8cd0bcb07f42a487b05f520128a590c8760e2f1e53134f758847c3fb3d19924a0fd52ce241e0bdccf58e27f4ef8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7d17a9a9962c32fe8dda5c70ab0adc39ae08268343481752513749aa299e232ba6e0e1cf592ff5089801be102d1a17a8f3ad7c18977c64ad8eb11a3823d0d73a76a428131e684fab0eec5df916a1498e2873caa0cce6acc21db789c84ae23aa1191bd2fed729a7963815326c418e338a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h576d738d06668551b54bba98a305bcc73d3a7bae62d7927dc15b300246ff93be17ea256f28ca669ac53e854366f805c725fe51126cf85fd4c2eccf99610c3b9f60c095f5834702295567689a16c922eb23aa944ede7a9b6502c6e98a71ad244bb15967d30eca1caeae5aa08f32ff77ac6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6adc0ba306817beb0f9a7d7ac90e502f22c6cb7ff04d01c9edbe8654b95fecb6250e8230b446b278a4384144f730432014250140bd0a1a5be0224b705522f7af8594b05e37c18a8baca9d075dce5195a059e4a95cc9884ce27b823e81458a3ab453dd248bdce1c8c849667de9f16d1e43;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecbdd6b48e7aabf63e3ecc782d2406ce82f3f3cc6d38ab168aa572db64f3ce4c1402ad23b212df5c09fcb055a656bd43fd051c5ecee14c457042d88f9f0acdfb95ae5fcb67544ee18764bbe9143be85c13d20a516408bc68174558a0f6947a5397ff8d68ef2250368686d55aeb751201c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfb314ad9b5ddde6d6c9201359b92c4e87b00ac52561a2e05464ca226c92464a7624ca2488f29c5b6410d89852eabadd52e4f130ed159c1229569c7aba86110558a34defed4392d35619e88dbe0f8d42b2acb66f6d9ebf0a48eee915cb695d7d2435ba08084099ce5f0c909567d724f30;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9a50163441ae0b2cad3b68ed9799f8d5d048ce26d5225445fdef879a2cece6286a8611bb6082eda011dcc46fd8ffde09f87f7985f0e02c24ba3f15ff9dd4132852ea020c698292b00df580994caac7fd5317603f531baf719eb40c0dee63a0c0c3d1120e7187dc8f5948821a5af786f7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21f505cfddf4bca3b9acef2a2d30e43c8e724bd9c5a70cc0d2a6398ec508dc901be8a8220c3dddf0f8090adec2ec7b1c4aef77c60e770e2f581ed7f5bb6c80ccb15317d06405be363bdc73b39948a6eb51083fbff0ef37b268b634a9e16e7900a4efa370d17240d166021a4205c7f886b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfac4f97200939845197d098644b8ca28e1b797ad47e77aed58eb5c09e59be620fe8a3adcb0a0a30d52797af97c637a4457c3674fc1782eb783fed115377c96a7edd7ebf408179718b9d04600f1c1a80fbcfe71723800f495d57c32bf90f49b825f69c483029c0f92b9f3dd0e0c7fc632d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a5ac976779d931999bfd43ac2cbda2b6f4462fad96d2f8877efa29c54b8e9a5c6fed7f8c1339178f1e83fd59fa2b2ac4e19c5c81f4e1b494f8fe0e9c9722fcf0c5abe485f709ca8c5add3353d754c607b9539a766d86705f9aff992a76a7ebe14ace707e73c758ef1472d8cf71886488;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbae7750f124a4a40ee4623a871c0185a6fa05143cb5f25e2be27ed19e8f6a7de6a86f88a4d56ac66710c141085e9f325929fa4de2b7592273d7b1ce1124687a50e5178aa594a895affcda4817a5871d7416cc7614c77de3fb8e924f433a2b7bc01f19936f1f8517d9e4e73a7d8797e2a3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd2aadaa1ff6950c3d8c08a229bbcecb1934ef4e6037b957493fe26f287a6f1888b3c3a226cd5a19370e8f7b335bc0b7e98e9476845dc3920d4db363a709eee3ce4e11e4d0dd60cd9bfff4fb1a9aeccd851891190b58eb9d7bb5b3ab5ffbc0bf6e4d63cc6e341e0fe398297e4336a495b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbaabd522e91ab71b300f5b881125d994a95c34ee273d9e2924f7bc23b8977864991b74da4fb69e4e5dc2b60bbe658a9421bba19d7e0e5d5aaaa2aa150fa4e8f20423c316507f50efdf7f3736694111b4894623f11bb437d86bef3e0b5f747bf12bf03324bf72b5d548cdcdea7b136f5fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc148b4cba9d943586ec36a703a132a92d4ef73d36e46c2fcccb8e9d95c9eddf2faeda4f71f8ef6b071c27a5027a3fbccbf3b8866591bf0c2149ecec00c39ecc2e5b33d24ece54f31b76d161123062c9b9a0277dfeab2a8afc78c6397d1cc0bd5a20a76fa3d0abdd78a0c62d02570e7fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac5ad4232887ed0116b7a469b1d6b35f2e3f93a22147455928f5b49c19669a7fe484c315e33e322a4a4eeb3326d88a6fa8824315c8a5fed67797765cf94d1997782569641ae7cc3f4b06118f9c20a5d9f9d17f57e6165eb172954b09a08ebe9c46c66d41ea6b722c25070d54ae1fbb491;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f6c7f40841fd824a9d7807da95fb18ae42b893aac48f1abcd73c3b41ccac9d84eb3575b3b4a0f57dde5a31140579a5e1dd2f1e2467d00a8acb3e8c3d3fcaf2ffb783a80239527603a0d0848f042607637b88bf8a35382f702f294c013e17db833645bcfae270e5097dbab33631764bec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h387eda2f7cb07744c4aceacd6c63a3f641dc6291a472a2399c3b8f49775be6f437421776fcd37116b0fbec7a2b8f419dc1af569ca82932fc3d0715980cba7cf731e5e854abf05d15caf1d0aa96e1700295747b56b84cc5f9055de821613cb1b422c35357dc3ef1975738d7e00894d79e6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70d0757335c9927f417f73021c8591be31ea1b05d6ca24df55305299ec1daea8510aeba27d46ecced4b0ff5373d89627d29262e4aebc8896b0378fa1884119f2a7b14d968ca521e653e2189ec23c183bc4a64434797e492f59414840993d53570cd1d5bb2fea80a3a35d9f4587a16b02e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33f4d7b6061c03030f0be2340ff83d276da8495cb5b4368e036a8f87cdaf9c7ad3a9ba6844a12fb7c5935b3ad4ef20b6de586812c36e22a009fe78eac6055ed5925d42185e2bcef91a573ea3def4e37b1f213d4285e319c258a59be58c1d81c38ed40fb6129d9d0590bc687442c62ed57;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3bef6ed7533c672308905fa5ede89fdeefd1c58abc05262bfb9c3ce34632c7ef234fd27a4f6614936dc1d8268d86ae0a30c260f1e8d1572babc10b69628fa4b70568faf437edcd258d8cf9333acfd5cb973c746e85998148d894d92acf7322aa81166392135be16f3a764a04d835251d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c336f374a8d739ce7ebd3412a6e4df851cb09399e80a481c6b93ba823d88ac85c150e9f8668619d12c4f935676a8b476bc241fba0df621c72b204394012342359ef47c1bc497f49c952563a1ffb47facc43995aaea255f95e2dd7d9ac1952782e34002c36a537707326720e1c75d1bf6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h878de7bcd9e087a84bdc33df12e1c1c30860e9302f5b7a8b0f54a2917c862df3362767ce1f10f9cb22d9a605bc686605f98d24652b138bc8260dfdae954c7477cf931c4f803a9f32858567f5b498636c4babb4283178267db9f2af3edb0fa9bcde97ba75697ee0878283d78f2606fdd88;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa95a1c7100a65631c19b458b5359fde48a2849fb69727af98fb6654ce776a509c77875d277a2a7ef9592129516e31767c72234aef62cd7524ab7a396eeeb565976d71401a2b3fb49aef2274225679e4a781ba25ef788c7eb6fe0e62842160bdd7815e3f4c38e9e481f5019268eeed696;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd5141c8509087ebdb2c144f777dc76508ebb4d105ef0b4561bb23c4e4f277e6c514f2850440cbe0839e5e7e4908c93b3cd7cd35cd2dffa3312ddcf10b6acc2eecfb3540a1438c486c73a126a3f0d024593f26e53342974603f31eaca0a66cc0e12894195e7b0b2617d48e425d388d585;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h728da592b282e93b1ebdc160417ce87776c617a8bd7bc40c086a40b32babba85cefa296a9ab81747b3d40db7fdffd6f4d9653a930f29599c832272fea85f80ee771b7dd84ce4308ee2e0ffad150f47b1e2c33fa272ae69f3eb731da22e8441aac1391f899cdc9de9673b84a6f0dbccaba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3769c8396dc8a5b663496d3da36c49bd6581c8d3ea0dc8efd8dc4052703c9c89ba30162fe2a7b57e58e63e3c7fc63fedfca83288423a91eab849f0b0f031a024a755e11c994e739c3b33956811513aa5a1870bae05b2ff188158382eaac177f61409cec3d77a2a062af323aa610624120;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93cb3f5a3fb228aff797246e0afc71235d684699fc64dddf786542b88f0375055292df38f99381f8d564f378ae2d616da2c4c63442950179edd7c59138d326241c1b87a1ac6fec0c0f9da210dccee8a3031bfb1573f727665bee56f87a3747a5276eed9161afe1272da613523d7103b64;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f7808a1b75d905717401337706b37c3ec7ba84ee4955a83a955afafc1e1e6272f1fad7a6079700a50c97b762b7fb48339b8db85d3778a98821d6a75fbd8cee12f99cb0ad8b7288a839736892109f904fc2880f7b149d249a4ed99cbe3c714b419d9df5a89700471c36a1945ffd181148;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52a0321ab194b9556dd3d5be071933c258beea97a6873725ce1c5e3117a3ecdec037a4f4d9ed1310f4d180147b08d57ec893cedb100b75e68262df2d3b00df2af962e2bdd901659d2019a95f75653de1062463f59b6cc2f0c25074d11d3f59fabcb1e3dad247fbefb5bcb3847664948ee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1b802f26315771d540a6710d1906e5ad93b13748e8bba526dfe630aa9c18fb46866c80a0a5c42826ae8b8b4e2f40ee007d49cedce259bf7cb6c334d9615cd856fb2c4987fc067b87c2bac2fc259fa1b9e9f637f621294b4a094de0044a3d05de4e1ea2cf3eeb279dcd6a209c77eb2ec5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d614c670f4a71c8b55d2495b8bcf04e820f4f0fa3f5fc610fc20ca8ea7a6b5538d14f0e91ae9485e8187fd47baba4c2d86d5075235d458e2c8f24fcd029bb9856b6b724cad16b5955a4b5b199d6e6ffa80ff1d796056a0985470645d18df9f7ebe6b1f7974872874f8c34136a913e6ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d5846d9c9421d1b52abc8adf52b5ff0907c6b53f349f9b13e8bc8d8e64d3c24982a169fa71caafd285ddb8d84873ca8e7606114faa89effa6af8ddbb75b17897ff7517fa44b0734665f14f9cc3d3475c7c7342fccd57d1b04316d26b43f18152c0bd87d43c4a340fee27a1792fff8482;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c5cf1fb5e6b582a96be8b1b4ff06cfa067fe35d1956115611c950b7731afa850d27882454dc04a816864fcdd00d88d57ae155cd8bc0e13d09e5446b37e63238a216200341061535698934daa09a42fcae574aaca2ef7c7fd455b1644ecf1b2e4928dd4c4378b2e9d609ed1726a7f507c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd42980ed9bb80300e17859c174127d488347e9c14475f2eabd37b51ce7a16ab80f3db0bfc6c44f6abfed58babf785e9112e889aca5fcdb50c34059dee9213816ef142f326c23da7d6bf2a675e7354b16b865e4524c1c1aaaad805b1354a507383fe0fc276bae0bdb1809004397432617c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3185da8ebec5fa9d8f6c85b892371b42cb8c45ceb55371e8309b32e1b63c2ce477aee45192e6509b1fd4b9c3beba50f41de77d73e4caf9483e3e23707c10d325d09b160477aa83730636ca28b22b447b1752f96ca2541747191d31c32d8699f6756f20e8e35a35779f7fb68def7afe99;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b7f79bb952a451f563bca129fd1aeb9b09a0f539d4e5dc0168a1dc64e88147014478ad18465a0c15202446dea037f689f71f495c042f82a92247eb0a0ba1a9941cbcf0b1b57ac2266c5b66579ceaa9c7a52ea0eb7f1e1cf0c503fd093fc3af5f73f9179540160a5df15497564e468a0c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2de7c1f477fb588db1a8d23fce8c5021468ba5ab61fdbd4f148b40aeb4b7e2c4aab674c92663355aab9a853fff12e3405459e2c9b5f82a2c54b68ceab72b74925b488bcd272263705bdb5ba34123520f5a0568559d93431bab616d5a32470d8b741eede288444f2585d487a0a39d5e7a1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5afb077989afe0322df39e1a1f9fca111b6b20ea711e4e4ce86c680c2645d6e9cf16499b9528b04cf1cd4831ed57e1908043e62566d517502cd16736764a4525a0359ab13ca28e7b4faac892686ea142adca360bcee085c710370a8456e0783dde29a89294455d29d8ae139f2e25ff8e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63b3237cc099b94c5c365f2c95e7d7299926f12e733e1c5a08ce028c28a4bdd79b998cac40d3ca971dee226893ca3446ced38f5d7e74a013b1df0c60d72d49e91babc553848a935ddfb9b7e2697e6de00b64338f7354930efe3d6456056791598c0d82ad0069123bd633a3e0f2c855cf2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53e53ce595032d48916db991fa1d4943a8392583b15342fb47160d6f43992ade9739b48431c74a0704b691246e6222278b37b4efaf3b4e8d3d96e3db8821df3426c4ce52a46925bddb274906d91f0bd634c6d5d6e4b7082902b3aa1a87845082ad34290561965cd7ec9c62153978b0ec3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf5e5c3ada8999acb1f4007b70cddcaf95f9c2bd8f14973ac6312b9eb3ea63ec67338f4bfa36d087576422fbeb8fdad35ec0ff29000b14d42f335fe96960acc545bdf3a24d72e4c14526d1bb3d330e01e0ee26944d3ba3ff2800f39798b97e982cb5474294db861fb65e2b4c324748770d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26ae7cbff1f391d36bad43408e9c39b9eebacf94cf1185836bf59f46f97df41afa854794c1895661a167214039e9b30cd720125d38e285c42ff501c458a31459529c476676396b8690be8b9f324cd1c7eacbc6f61b2162e1c606880079cced7901b831175d29d084be331c045edfd2394;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7d1ac7ae8561e4320d7b1f4fcad3b078220818f5fa4147c3aa26de5bb919d2cfe1d2b6793727cd7a6901433bf91a84722d3cafc00bc1444c865e25d0f52447e1a40659c53ec998b5f13d5323c415f7f47df17b4a76705e705a9452938f59622a387efac7db73a53a0fe732e16a8f005a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h919bc3d3431176e1caabd66c82df08a251e23f0f2a8a897b1cfe75061b9b519823c375488422719235643fd83fafff7562a19056e774c4c6cb5051b39d75accd2b5f1642c6668235ea0fdc4f1d8a3a1bb929870838a447962c42fbe5b209cca52850852dc8fd104fc8749e32b169ee89e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84f28c2720633c8d51bb8a13e5b208252856cad83e61a2b9fed3ef873997e878dbc010ed1873bf84681268d8daf454cfa141f57f2a544124344ebeb13077e25f99d1e11afa3c6984b6e8f78505f47719167617f3ec28a0091c69f1903aa6043f7ff30ede806ca3d9d58ddb7fa11aef0f7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4be904f67a862256e4e59317e4c89778d081fb4fb678616167cdd0d11dd2a5b4858627b867e2f8b86ee75a7fe4953b06fd7d945779dab38eefa49b17e199a72a9577db994de3d8e8723b018e1e4515ef056d72b7fd91ad17bbf51f1b2d32ad31754ab955518b6a0ce9c81311299dbac78;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b6cf3b13c169fdb0bc06055763027b749ef2382d41d89830bc3a1f98852eaa79394eeeabf4a33e3aae900c31129f59b6571ca962ac55d3bd145bfc26f841cf361560b32e9f893f2b0be9976b3cb8e061c3a7cbe6a3a36c23ffc924714b6e52822a84605e14f80d9b127caced1ebfd852;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1a6fbd8fad107b850adc819196d6fbecf27c9da779ee2ce1584e352782ff5d916f4fba3e816eace8fd8151ade7bc38b39032592703fb282f1787b415f130db1dd8836623dd46a03078c6fc38365a2ad0f4a6aa6a7b78e7ac0529625eb9359976402428e78be542780118f44a1af63ade;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70c507513802cb5f59bca23c2488e03e51130622beab1804f70c9397ab9e91cfd461168c0bfd7c92868bda8259ac25a9d758ff472dd1358e1f56dc4692ca180b237e442daff9bd53bcb82176ba7afae1c9e93fdbe75ef618d8bc29688e249c76faf4fcb58cbbe9487bc62b3b2378469b6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcad362531145343917b69dde5610b24b1b209e7c8b0d7c69353c796287c08b93b2de3b1b67484a56d60a0e3ada87c4393ae9234ce5b190beedf0958af6614b7d940928ea44b0d9e27d2adea49b37e86980b87436bc1f12a3e6c76a4e121f212754fd6716cda42a9477efe7a9ff7d49033;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27089545487bc3ba8a96a83ca1271545719a98f1fcf2ba8b138e161ef97a61897c80eff89c1842062cb0f87fadc19743d750d4aa59fbc1f7b71aed98e1180abe7492f39158198339a122112d2b67b0f291725f99fec4e403d4bea37fe6f29f923ab224d5baec7bbc3b3334401049c6e63;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74985bb4572a6c704573f073b59e7d29dd9234500afbc3032cfd9fb450daadb52fd4422e4c3295663b6b668a11a4b446d38603997189fd06c5c6d0755fb89b66859381ef5c5254fab288681c677409a421583486b6b98de2ed6aa2f5876f72f44f5991d61c12e2bcbf24a01c4452838da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h518da0d3bfc5d4ac2ae2503aeb5e3bb5804324106b32159b9b21b9effe34652a54895170b533d08b6b93d8edc888a9a81da464387e790b9e49b60e1d5d51dd07a837d9a6149dd1cc71b289680285513e2b22881ba35a67960e3b81669149d38619eb23a774e9547b0641661548f29a47b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h273c17b470da09882c9845e63bf14b2b9536fdecdb4cf1885f5b5610770ed75d117a75a5f7a4accd110ad4fd3202d984fea6be39d2977decfecb518aa3398751ad342704b03c034f8dabc0032bf3189af90011e0fbc737b354015677a1f66f7b2a079d6def6d945cc2b3a277adf44d260;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf96a59d44a2e4c23119b9a965ba30d713326b2c6bd9a5773f18af014a86708b69effa61e7fe54c8d9b7eac6bb0ee4c7c08f0f0ea112e34824f8394991497103ff04237a7db203f3b37cdddf6b2e5fde9170f65179ca775690708072de367dc01cd41b7f63640aa4a6ca638ce69b25d64;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h673f42106f92dc75cc374eddef7704640f90cfaf970809ea4d1ba548584dd433080aa865251a1bbb35014a7c8677a3db85baaac0d96002c8def16f3aab300486ca5a6fabef25299d359e79569409172e49f8e70610905058128f33da97e0dcd71d5649b2aa72df27f95a4851248588328;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fc8252dee23b80acda20311d01ab8661973bbe04d26a4fc8cad7c4d45def5e29b2ab3a7b75a8ac7005db5f14b62a6680a35bc643b9db3253109119d8e74d9a4663caf37d68146bed0b221c4ffd734ccec202f9a2f2efadccacb038ea3427c8ed4ef8f5490ed9da87b9b285a8a332115d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52092eda7ea8308a2e197a57fd3c6d0759dcc41ace15e801288993b1bb05d21cfb2cdc0492cd6d337cdf7de2d5f63c82877d5cb434a37cb75e759e9688872cab40644dae908300ee90ec45eb046627997cc1f1f582d3da7565926fe1150976ec423ac6b81396c62de47ba8f0f0b07f7e5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdc21d24017bd0d22244e89db103b48b250dd22e92658bd43db5dfd2724cdb48b5a53e24e9d131c556abfc67638ede5332c535b50800b563a6715fb752fbce6fba0534caca4d7d2cd02a5114ca442ec3884b498508106ba4e14d9cd4c9c7cb87b83ebbc5bae1c48974e3f0e47e671c9c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3aaecf52411be9d991651450896923c60530652666ef3a8e8863b5f39417ddb2ad1f65944da0be13609f71802a70138f665c71209844fafdef51f8e3ef9155155ca222e647008d036eeb80efa1ba18636eda5aecfd929d719b80de1ecba14e4235f0261cafc80dcf01f0573ed0c983597;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0839944a3afa052ebdacd927b0212669154c236755873ca45cda785764a737070e71f2c05368ac3302ce42d0a5aeb8c9196a2e6b25811689372de3d944a7093bbff135e776f61199782008a9621ed64ef312fe7e0f5425c7c8d94cfea09340ed98e7b0aa4fce7cdda1b64a117380942a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9369122928e89962a0cb7cd64938bf691380b2c9682b3b8755aa2317f281cdc5a479da752519f047add3aa39c4b70926a9196df9302e8d7882e9247724222f5f10a13e001fb526b381bfcf59eeff25e0fe768c36477556877a267d31a14d2ac3270a264d6730894bcce6a6d8f07eb0898;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88dd801a423adbbe993d1863215aed7dc0811c3ed8913f4362d37631d1a8643fd3acff6e1036f1037ad15d69c8a1f34d743521f8aa37a0abc9626b391ae9a93d93a12937a6d461638fb5e67a781328eaaaebd5063907a91e3648859476daa0d3000034b7065d7ba6104aeb1b34ad443cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h213ea3e1e531613d0df609e20ae689adab417976281dde2762dbec5e7a4152ee0669864e3d795534e285ada490f70a5ec6e27ed1a45f1956eca9562f42c479c229caa87e379b1474b88c81841cf9202bfb94df2c63dc9918d3ba99aa823065de1c0098d8ed344af539d17b1ce8fe36aac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h234769948a1f20dc553c0531a2fcffd289f502edc14a90b8edd1b6161e89db5b6c2b2eaa2c7946d2827db35c6caeb160ee7f0fae1a066cab8a23cb2c77d894dc68556c1bc69727017333559722e1e515a6f73f92b3e90fbd158f46f5cf2354a433305370bc267c6b9f56eb5fe35cb4dd3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c2a30de7639c66fffedb447fa56c655d1ebd76b122d3b29a28a71588b5177618b629f0fd9698ea91364d41303c24db3e4e587ea17ff5276148101a5682a7d345562abecb002395ead5473ce1e4e4f7aed1a43fca59df3c59c7c215ee3a2bd33c429e6c12b2c83a812e44ac5b36b8d924;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'habf9187190ae3cb38caa89f7ba394eeca509ce7d392763da5a8bee8a11bf60c0951f82c6402e9f1bc31a9ea01c1877ca9c54145a7e3ad2d9208c20d99f42836c3ea1a5d1318e594650d189bb20f51dda59d7e3021aa6b3301633032c217643ea320e0ebefe85d5bce8b05c286766108bf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf31769688c34c3b4a25716dd1325bebc2ff499facf2faf8c34363bb19a1a260e9287f1afe6efafb5512c810937fd731b4f778560adc4f0ffcf935009ff61dad9992480644ac553683f20dddacda8b078e99247a965a0d520d6aa5f5658eef59d6591ee9c179b0d51ba97a57dcc42d8c66;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ec632d9f4de97e717fa89359470c63d9fe73da7f97226904e476487c038acca5ecba2b44623c70a84b8e0002b868a220085252ad5df3a565b327d39b996fbb50dc3c2896c6bbbf61dfef742f3e294d54a936112066c11ff98d41346701abd3bb50c0851101f25c5dc00aeafc93aacef1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc5fa6dca4b7a278d37a80617081e1a7dce64736d2de8c14929395d0faaf3c82fced1be3d9ac9850e4c56accbbb9b36d473e1226b617638dab2e25d2cfd7548120a8b27ce7ccd9aa459dcc25a91730371736a2757219d2bfeab5bb0b4b4cce7a43bae483b66444cd7edc87f4b54ce9e58;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7bcded6faa034825242768da12d8a62908e52dfd2eafc52cced33512315085adfa6265ac346f2923137f87df3ea3bcf025d369fc06dca90facf6bb2aefaceebf473910375969a1ff24bace4fcb73028b50ca1bef8421882add224b49e899eed35f09c2f58c4d5f4a65dffa65cf65d2644;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h354d98c06148cbfc1898766c388d89c980035bd34fa705b94222122ef660111ca36411279cb5c841b348d0f4eed71e5153b07b8a4e5ed11f9c59b4284ac50a894ba098f19a29e914f887918dcdfe14dafb2a8cc240089c4dd85b45bf22177bb3ef7770ff0823a1757b0e40830b3cd5a02;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6859fa9500cbd56843433517df5ad52a797e019ce4079263fb4f5362cd9cfebe08cc63a55a53a807e27737e9542a5b16990115b5572d21bc615a2e4c8d0ae846e5602d9d5d0e514e4d3490d95993477f0f2d13bdcb50b7e6ac35cd98d670294f9dd368c5ba9683e525585a6ac2b667185;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5eece0cd188aa5d0d6a166994310614a31c431510bb0db647d7da0c0f4ad59eeeb5ba63ca435eb39cf6039af32b845996b45697c7950ba0171266dd568113ba4f98bc2fbd027db286c6159102d25f67b5cac2d4b7f89bd6efca1bab63e5981916256457461de76fbbe6fa49ee6b045ed7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7cc7fcccc4edbf098559147adb5da0d2c73cfc1a3f4f50fa3356e01a412ddd8e016b8bf9941487f9a6ecb253d161733aa56843f55c80380af905997bc2569344b33f035783b069cde73a743a3ffa45be60948e06fd4f333effdef5388b62a946dc2b0618ca01bfc1eb8058cd15ab7507;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9be7d4ceccb7807c8c50d0fde6f587b2b39fbc9aa8530a005a3d4767db24a0d4dd6c5354e02ee7a2e26fe2551746d7be7a4add5d9a27c8ca76b85ed9721d3b0355cf523b76be4b29aee767a0ee83f0f6b62d59b28493f5de9548eb14d7e0e79354efde1abfa3b083ce0268579eda0f06;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49fae68cd544edafe32f7f0697fd32aa5fc6d0868eeb7653288ded5c1f3ae848b3b5f6c96099897d686a64cd9ee2399879a7b1571539d4660c41247f3185d478ec4ee3b1a2d6c912aea79418e9c4a73ada7c02c6da6f68933caaebf2cf202a81c431884100a97435935373479eceba98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c6b0e0413460a2d282a8bc19691ce7bd04c310f395cdb2091a27f47d996bdf99082fbfc4ab35f25aa32a80ceb852dff0555e6ff2fb608a27b74d9a03a606fe3a2e2181b6da1bdcf7cdd2fd5297bf08d46accc378fb79e94f7210f63d39c0bfa5f361253f22bbdab5889b5a540d3ecfb5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbc58c1e657742c446118b5951aa1d1b3902345218bdd6d5937ad007784ca49686c9ab576676ee32f0bf5548e073f0e73a70d8c9e10d8c2efc166d4ffaf04c42ac9ae2233fbc1c14c4a9ba87d69886ef17fe28d7f4c2015f3fb25a0e78511072526307b3437d40924d714f433e4dc7155;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h36515d72484bc88cc351dff1d75c7af6aa3d1b3f15b7817fae2eb38fa0cfe0345efc2c308546d5dabcf6026d48400785b7c8b9efc9aab355db400eb6872d9960544683fca33fd39f49aa597a712d8275291d544a17e8ac313ed30caf5223c0507577136e64f1d3efc7d781ad96c21bb25;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h925ededfc1c5ab96ef797a1c03f7ac0b7ba63e1e7b4ef019f8a8b43fde4bc218e6baf5be040dd57c98d54842433a2cedbf629fd942e401dd9c254916eeb8788bf899749556f1628dc0d999d9c3091ed38d5e0099c53a19d840f378fa868f0d612ebc5a585a1afb95771c7ebe5a4b42301;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e03f3902a2ed25c4a2c8e03b34d833ab8a76b53ab11a71dc5164b9f23950de992e823d9e9546dcd38cd2974f3cfd4828d4f762c8daeafc12a3ec6c3021a7a0ad4d8b632be2c31a79666f0d47365637809a88622bfa4de89813e4c59ee9cd0346cfb51278a717e2ba38fb05e60c347c5c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h294e6742d763dd4f73aea68093f631e41b06d0755a1b6d6041b94b3911ce8b518efeb44762c9f03aae45a7deca3a156ec238d45938959acb4aeccaf623a09138ff8228cea5f9d2c039d0b0fdaf02b69ad679781abdcd3b4716435a53911573fa3c12822f38ef6292a75a637e0f8282fb2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h174a16493ea7979e909d2a0e849b986227b5bbed8a617dd7b7bd57a2a63e2de4ce06a4ba41e78786c21e54a6d4e8d1992b72212a65179191d104a7de6ccdeb6952f3f9ac443c269cb0e43ff16f39fe494efa931e10a7b04574c3f46b9ac198c05efd8c3027839de831d729e42f39f4611;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a199367bcd66f3a745587498f32b61ab06e440ea0c30d9a43ef464e7655085ea3eb8984ee0eb552b26bf9987132b58fe4bbc83d48e45aa4ae21f3ac60fcdbc5be319d56fa69a1e830925027651d1e349152859f1595d3a8ee1f86dcb307be3772e24b2cbcbdb6b9522fd7bed062b544c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27f231fa11d9f46ba95ee2123126e426743b6b1b9317af71f8f113cbf68be824a91fbe2c2ba20408b9ba9fbc7aed99d16d8a0fb4d0801aec7e917e34fb550ae203f9e00ef8e9b2af95ad231b2923ebeae7b4479200b2b6ca6f3762e7245dbae2a058703e0f4b727c9ea9a6725c9527f4d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f953d7dcec794ec360e029449258e5d3bfed3d032b2cef4a95a2ef40e95ed0b03e690948542069ae8de0bb7a49f2ec9b6f880052ee691c63758956a7d35c1cbc3ba39443113ca8592dfd8bcb3426bc8a93d8a8cc1e73ceedf0c6631ace638d254194d2d9713f99d6bd6bde1c5f0818e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e6b145285a41e7b6f783f627ffe6c9cdffb518733b9d4bf41be894f3ebaa7a89510f7ccd4332cd911544b929262a39ed22a3ad489634db6c27bd23b05a50124842940209238a9fe5e14363463c4ae2b14f9eb9c193091da95262e6cea760937949c78a16d437b02b7a34689dd9aa588c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1956d2ad93caf2fbe157b481c8fdc69388a21fb6aad620ad5251022f28ece8e50683617aae6424116d8e3217f32788169109c57deb6795fc61633a121aa27ff2c77e38d9ac2da9b361d760e25749355ee78539d819e11455f548a5597abf658f7421d5a5f4f1b1439d5dc2830b3aa539;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf70f6f4cbbd53fdfcf0e0f0239d7f861c2dd9228c9496d014f64cd301edf5f1b7166dcbdfcf6e0e6cc81b4548df7216006692bf5a3cb26bd069871924343bbfd6f5547e8476a7560d79e1f17e547c79a42e09d28270af26a7ca04f205f3b8abe22c6c7ca385c814223a23ecf54c165bf9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha61d140c75a94c572d6742c2fe1023180939c02b5214eaa19250a89896a86a34e360a625a56754944db53ee86082cd180ce6f28eb402a1161ee89bc2f5f059a0f22d7cafe8826103903fcfc6331ab2b5d52455239769d1e389aed1d9dee003af89710f4a56f3f31a2bfa11771227ecedb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d6c9a28a2e76f04a31859e2778ee9c238a6264aab29b30e0cf068173d364d25e26497b802033c2e1086c70f150140d1cfe914843b4293e825d59e64a90cad7eff5f22f0f47b3fc329244449cb538064c92756d2c3740e86e1c1840b18b2c56da503055827ceae89f51231657e25706f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28f53b0aa7abe68ac730ee53b7642fdf021802cd0527a650b8a1a66c6fd348cbe9a4423f7e35374a9aa6d89095e594530fa44bc03b70a612dc7ce3e5b6a74c95390a73c709425e8d664044781cc9d1e20267f02d8acf3fbbf68a0f0bdab6be074b7e7379084c280fab4e5b1feb4c1b4fd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ff57a0fdebc40d620743a7dc7aaaca7401f460dd3403b10a0c055062a11b13c3d179f46eee8660fb86bd23e31a81ea46caa6463d013d4c8ab7300b655e33a0c931b3e03fea540cca2dccfe52286d25cc54b8776a2997e0ad2e96a9b0a8a3c4de4aeea704ed3bac8e69c1e283bc6cc5b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8280344998ce8e0bdc0a035312830d3445fdb1d94dd51680f327cc6589ae25b5bbec96cb1bb70b84c86112a35c2861e7a7a9c785e079bdb2594e85e57b2b4f4e81f9429e59ea57d6313aa20fe2ce74c01c60dfdbbb437d27ec4ca1ee8061da124a77a059dd9fc19fc30d92dfe0651d12;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8dada59f28a3d5f26f3aa22d021a5fd573e7aa44141b5524bc7710ba511662efc4e6ed336a7bad6ba1a1703aaa223d6b49125dbf549cafc3c78e132c17bc755f29da6f3b469c7e1e62c98e0ba0ac58c6495fbf4e762533497faa8ad06a46e6da9e5ef3702a69febd39811b471859c1d88;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h675a7ea26094a7acab49852d2f4366ccab51d9caf4ac4cbe01e2ebbc79da0548ad7ce0f512ba1973025069e2be47793ee91053b9abe68019b8b2dd9ab25c590a6b39f76a92f0981598993069088b31407928a63807d13b12bc1971b9cac44e7066300e50cc9049651171030f0116d7c24;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88aeef32d3b50fb89cec8a09c3b2743fe2b00ab138c9e26870ec38267da864d75cc1c61b4a78857ef1995ae983ea24ad0b589a6f14f27188511f0ba49743b5c057f5dad8c82931b31491f73ea9e2a767a216e6c236255c556f99c2ae94971def492a100e1c71dc65ebc42cbab410df814;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf366924f048af43853fd73954a3fd16a7fba79a5a57703a5897503bf73d4ccd105d8b100df4fc265cb52179b7ad5650aeda803bc16dab3750519bfd27c958ed249f6c27edc79bb3a3a5b957999cd67db3dce2bdbd1a47c58d1ebab01a870f52bc1971f73c5bf916ceb6a4613997ea6bf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20428171cb57ad6de2d12bb76dd240a6aaba5e12e0e37f96597383af14db03778eb0104ab30de123d5f518e1acf47efedd7ab0c39e00ecbd808cb7fa8e66ca3f61ded9d1df9a8a0bcc7137cd947d91e09e9da6275456aacc3ba4d18bc0bfc7ca453fb81c50c7f90ba0908dafbe3f6d4e8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7dcc4b8ac8f4b8dac10e173d87c2fce75dc3eeeeab021be3dda1d5898740301336964a185024e66f0d4742a991071f15ea316784ab9dd3f51dc34559a5220833676a539ac1de46326fcfef986cc83713f2f476e15c319ba6ffa9c6a874b1d309c6dbbbab76d671b737084628b5d88ea00;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h338e6a7190e141af1c26440aeabf06a96c7ba73ac5dbb03799b09e4822cbfc956f9d55f52e8fe642986819732aea6145642089aaccccaac44c87cb835910d45d38de7180ee4fd5fdf2237cee24e788f5fb4eb7576951c339424376b633d9df88505ffd9ce6a33fe0255205b5bef809985;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd3b623509aae026910830d7c6c61e215759765a9fff1ba783f8071ae1cdea4527d0a08b4e1b6029aa840c5513b7183480abd9fcee5c92e6f6f11cf996516334477591bb44cb2bad02498dce3fc57d4bc2a4ee24612214537e11fae414682776663a9ffed53aac337ef5d747593dff6ea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f41bd35d30938ead623da0b9637a33c6837e9698e5f96132f0dd444af97380133c1cfeaac93cadbae462049ffd05cc37bea790629364cc8de4321b7009d47ef79b366f4496dd504cd5b243acf9cb0ee99955ec8fadefcef4061731b65400d10683890ca96e7f1362ad47ec38395b0a21;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1d2c02cbee563f28514f75b3e16b4af38c538ddb29fac8336333fe186dc006787372d3315f0e229ed90c352af32da26ac287cbc729d9210f128c348bda5d828d2b1c31ce3a49776ebf48fd2a2f5c5164a67a3a247a600e3d3040be3c005efd2bbf9db690b78d8935c6b1a4b831699d63;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79639a239343ce50614d773f70feedde869094d9e3148e89755859e917ee18c2cc93c918a68f981857b2b81fedb819ce555dd4b12d8792b8dce8bf8531879a3e789749d603942352b2c5da4a7b8cdb5ea59b2a3a6d231a7f6eaa94e9d0ea7827f3d194ceddb05478081b2b1e121e4e2ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h461a503f0c7bcccf5b086a7aa1cf0a5ebb44549f4a1ab87e8559d87bb6cdbbe9233646e21b898a6af5cea8e82e7d87ce66a72e26bc23b3700e77ec1f49e69badd2dcb0e35aa0d67c6c7a3396fba2f0a3af95d046f46445c2b01167b6405de6ae36709addc361d124047e4996a8322da4a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb60996dc37bc3e6f9458b6a8f98382c6a9c4ac398a01bcb9b8df424e1df9d7fb9e6720311c4fb5f962206077295aa15b297b5c411c91687935949f6b73e7aa2b8193885311b5187be88ed7d62f9e5327e4770912c07be46e9a0923430741b7cfd8e80010bc652fff546985c8a5cebdacb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3cf42af7fc15443d9b11bb54b8668e794112eb4b7950662017a2d35c4ea09623a8a9b4b20c427de22403c1ddbf86ec601e641beb943e0e94a241a78cc024fa1dc7c038e2cf67edef8891539457198ea9b11b31f849b6c5d535c9bfb9a6164a8c32709dc9b0abb8f5b5b95f29de03d695;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47cd2a2b14ddaa40a733e41a1f6ec0b01e4e46acf61e2d52cfc0901eb299363dc0bff1662459368b91d69c255308bcf7e88cf111ff6558a08e80b98c8bad26f3de2c343857538b14cd38b5c4e184bc981365817c8aa508dfb29eb699c323d1e93a18a1327f7e87ec1889471cf1166d8df;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd15390586a72e7f0312790f47e62abe21a31040abd632f49c862e44e1f5bb7a7438aecdb3dd38b2854c89f6cfe493fd594c8569284bdf9fc2a1ec1a54ac1751fc4a40c5dbd5f07818ed102165082d911bbefdfa69ade4f4e507ad8c107221c951e60777bfb6c64a112be80f90b575e24;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h747781a012793b1f4e7a8a86b2027ce3897a8b28bc3c374085ab97c75c67524d5cb702d93c641a7eb45647f916c257bf3937257786481cfa327ec146812a3108705e12fbb98db731e39d1408f64a15bb07f308595ec09c14b436b6199be9474b2ecab751badf81049d902fb194d4ef16b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c386247d08fef14c63075faee69f029d22c78599dce30dbb44c87efc2ee11dc131c2c0edab398e56249488c74a65fb59e0ceddc86831a853e10f801ab86f1c5a7b67ae5927d05564c634ddc20fcbb61323a258855a251e41b478bb122f7bbc11fafc6a609c8e4ecfc3a7dff3f1420d09;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6e69d437a1207955713e2275e24b0d4896085560b838be251351740e5733af774b7e78f910de575bd219e336b38e25be4f02b69f884560bb33fd8776d8e8d6ec128b4b04481acb73e236453a8b6a8b9e0ba87d9326024008b90f2e8026b32d673353c491b4adeb23f84a55a1946b4da1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24421915d3f799e7ebb4a24c292d95ee9d55f20a70b7526b3b460262ccb2a50b73fe524bad8dacc5c2b756df57bc9e606f981c4d6d1e2ffaa2ab7546833f79812fed683f5abbfa0dd8fa195bf90b0b1179b1dec9b1d94366f66b5b57e1027384dd3991536c0305c93bf6266da489643b0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6632d7a675fe26fc73d5502a9a508987adacaef5ec2719077a484390ddfcfa20903a4273fb7d32451f9e63910c35080b51eeb4c691af98aa0f116633e254d149344341ebaf1a67849b2bfe17afd4091b033095b8e40689f2e3f4a05649f62594cb3c4def5fc7da8c6b205085b75671bde;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc23cc9ee1bfdf4680ddbe644cd7158a6871fa8c476b361d548d31be9b2c4f2bbe0822f20f559be78ddbbf1c7cfeb538a33b6544ef0796adadb106dc6d4b72759fda0b440068444e18c0c2d2b326b8feb5a0f405f4ad8b77cc0e21d03d613f6c531d356fa9b2391bea93a81c7bc361935;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16c7b8e383fad79334e83cb1472ebab2060460a240d3b1b982615ec45c496319c11ea46c79358e8aeb6a0b55dbe07abc1e19988ad1bf2c4d1f2448cc480b6d80897c631f9a10169eddea45bb0b2cf85898afc1def96e92ff0beacdea584587985e388b69363f5eb784a3be5628e0c7ca3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb775be3ec2fa75c5c7ae92339d7be7a874a5da7b704936566c1c5c402cc1dfeb9555117b4913416ef2ac069ec98962fe3356cd0bf73ee308e983af76b3a61cac818612b521829a2f0625754151961e339be043562f58e3ebadd9732aae57389d3fea9efe1faa67742ed55e4f3eb070ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcaab1887abba5b6c117f8388418f944a40132eba579a63c8b8f00791134c9e740ff30d3b247df9c4e781abfd47c374198e76c5d0488562760d94e825da6d74818dd40a2ba9346cc35e5cf2122c5a6acf63ea4d051aed897b44475078b93462da2214c82e426bb42fa3b57122da8abf2b4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf16786c96260cf34d4d457bef33a00fa405bb307d8dd12077b66f89fd938a5b1a42f39a2ab55e9501c7385f48546738e0ea217fbf16c2c5d3618968a0d624f56fde69705c463d5f7be633fcbc7ce631b11892b018ebfb1a34599db75f3167502d09b0837aac042d722ba51ec0f4ae41c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e6a0464add2924819fcac5a56a141d95263196e62bb8776c8532002be92c2adfb1a5c901e3e7b77ed69941e183b9cbee4f56885873c96e35f36a607ff5b1112c0fec9b91bedf71950a5c9d4cbbe2f437ebb8acd4abe393d1fecd9534d5453964418f112b3aea18d120e2fcffcdc15561;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64e83363d8f6e847861da5db7c8bea815a9880aa94d441f30e7a0c264f958708f771c6d4c0e1f7155f170698e5429612e4017fb5f08b273d5d62d06dd955082d73dbe4ec34a7ce8bbecb9e7e65a1fffc6718f14ecf8ad759b31b4015d599be759ccc36e72ea4902ad88a679c183fe33ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f5559fc4af647c5d768d6f7f88da0869956437ba06644b353deadc57aee32c1f4c7aedcc70a8274e7443af93e0948e0505112f5d63807852af5f473a3668c059f955500e2bc5d6393834d41c620c6bdd3f8d019c72a328fa1726dd81302eede2c1aeba48b0510ea12b769aa035cc89e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h145e21f4f88f39aa9463c7e9844002c383def2e8fd79f4e492ab5b62e63c8e041eb3ab0c46b14145bb5e254933d7595cc9030e275205e3080edff9fac365015594b80a252c915f7a8731279a1bf54dc3c8db79912abfd6a45cd477f08e08157caa25d0c4473ec6f800935298d433fecd6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd792404c04666071dfb0c21185326a602e0fa9f7178e629b890aca3c49fbf5255597b6b84358be578c86226480d65f6419e03f78f48b1d0bc75997b5eb35535c7fb21a760420ed7187ffd9a35e143705135e9868bafdbfefda9b69601f956b86b587a91c66174f3a0f1d55d4facfd766e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf72e0bd675260cc81ae0cb404af1d8cfa7d0ef8009be49a9d42aa129f18ba0cda907ffa44f22a035df3171a46abc6587d76b07be7bdc2b82d83994709d946e6254548feac20263765dd2bbd57acbb466162dc37f61d5431fb3993f4412708ffdb0102edf4e81f1341ec416c5438ddddf5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h812a30dbe7231dbae72254fc6cd42f63a1bf9279b6c69cb6bf8a79540083a3398674f8a20b60da147457622687ae087d84b4a8d54f9a07dadfc46d742e086266818470db528ba86a71e13ab06c8078bee01c5950fb1345f55fdd6da16aac800013d3f816f3c02125afbc12339173e36e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25f9d9784ed050d3eff3d8f4ef3b08defaa4c24a8f472c598c18a70f88d099c7c11c42a2636de19c2de5b051cf56d500430ea0e9dde49b9b473485e9135f8288c6b02fe85a5b9bb5c51a153356d0d8586a6e9cc108f08560b5b1c38e56a8d219f652adbd743a76a38ebe890b2b4ea63b0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd93c391cd16e2bd0aedfdd29f6e276e1783efdc002d452e6e83dba821b47c7b40e95e02bb96b182f9965767d0954643f2b543725018db402ddb0a6b72e52d58b9b83a85a7b9b80cceafc4fb24467c340ce1f8b64bdb9765213912c92b37c92d5bb983c52c6346693a1925502ebdbbd9cd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2615f28ea49ccd2888dc66e40627059e96830e930cf8bb079e25a166cf47be763abab0111464bba1966f11d5c02f9b818f208921ef90b8c328c7569993d099a10aafe72bd47884fe1812602c1f98be85b0fa9124ea78b1da5bbc1be434444ae87d78b21fb25c0214702e1ecbc9db03b65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90432c14986d207ef2f9cb6ebd8443d016cbc1e23feec17fa7e615a63aebd767f583f7f4f160f7396bafd21246cad1324d6e7e4149c4efe3aff1dcbc195160eb8c541d98455e34dd5453983dcaf681df2b692bf3352f5255a1633fbb1b41d9cd1e189d828025051d552f04a7dcfbd9ed4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he88da18dbfce6737ac76313f673a9582d931295b13b4e5d573594a980f1fc9db0d9e3483c90ae46d5717352b524f045260778548f55ae12d925c92a6e79ba4a12dab14f99e69c891687692c4c9ec4fd2c6154e60a1aedf496e8ede77a44cd5f6e173f6645442b66951bd974d29386511b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc608254969dc2e5a9ce09b40d9a0a1c231db9b6247d98e0e73b55e025dc34e0840a7d50060af5c6cdbe804d9348b6ebf23bb6d8dba7887cc1bbb841eeffb95167d147bd7908bcd326eae326ee59f420a931992db15b3b2c2683e30b781371639b3fde697526f264c5919b63fc9c7b18fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1a27017074cb282343e25d6c93238377dd831422c2ee717b13ce5cbe2a6f6fa6b99d1cdc51cd27fd8390563b5a69db3080dc93881767e77930524b50b04f448900960acd33251d14985c6944beee6e9419b3d1b357c7b3ae6bc7dd77687dc24204bbe180c28913faa2beae2aa4ffc681;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd44594e40abbcb3a79f7addcb4e6e99ad411b49642ae36b0c3836574e7bcbd986499fc16d3ae166528e2a97fd27ff0fbb5a52e5bda9440e0b64c0d0d02f40f0a24f0f726f6959e6818b921741f53f9a31bd256e4c5b794514ef3a15540cc6b1751f76f32be1a24df9fd3fc200d06a2e9c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7a1981cdadf05533f5502a2d7a984f24efe79250deb95bee88df361a6a6306066d9e8b82a86e39010772c2f1628291790bed56da9165a4e590245fc42fd2dc220c2f21466e90446da31db84b7c99c9473852ab20f55ecfb40c4f58aaa5fda4c997cc361f74b044da42ec4a993444efa2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb60201a05883015839d5beb5f62fc3f95c59c9317d44b612fc580327db9c6bec0d53575a3e3cd640619e303c2e3c41dd39c15a555ff9f3e61150db5029e2387bd2c9fa672a796d7e21e82cc865d25375b51583b5c94e6e961a92e7e9e6f6e6e0e30225c14a0031ddfdb2b71b015dbd0e6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h590fb2d7395e6d1f778db1ef422ce6aa89ab08fc24fac91ce7b2f21b58cb5c72c7085ef95993143b719b9f8f40626a52fdd39777f91eb3fb063d2e6bd51966809dd30f78f7196d23e6c163406fc2971c9f9c16281113adbad8532832983803d489d4c2c8d1f98d8739f2a332a9731eea9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e6823e872a5a7e78cba7105fc219d77257f1cd2c03470a2c04fe69c0895882ef817e0964c4ca2c3aee368dc776dc2f5011fff4aab2605452a4e9b839302fbea8f0614f7c94a4f03b24a2dd3795ef0e49153408607477d4c5ae19412b89f73cb63f94fe9321f5fd89f56dd6d486f80aee;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7af28e2e8876fcd5e81862145c434a05c1216a96b994a35145ac9bf79f640e8505bc0a79af46357ae0c8fee57381ded9df97089479a758691446c08644d140c7eda0cbcbc38cc4ad9f7336712510717aabc316c4ad9f722703808db5f951afb683e4c27439b427589b06105829593f412;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf792e3ec7b58aa647662a8f8ae3789204ef747a4836149becfdfb313f74053ee4bd478ad3adeb72dd08546c9a20c7a9b60723ec9afd18d000a99a3bd826bff280f23f30c39d77f2346e7329d522fa18a291e0479ffe7314e2cb233fa7d2f04ce71361599695d15f056422633424dbf22;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98372394d0cdbc35517132041996b4cb82be7bc43ea4f8c8d46a44fdcf68288aafc7c8840800f5fb8ccfe840b5f2c13b603dff5620b2a2fe750fab26fb77df1b303d9d81f33830c845a9cfb21dc8e1df4bc0fb311ccbbcf9b3fc99f552cac61ab30fc076eb3b6c4215b6654b985c8279;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccc3a3917fed0d71f8d7de6653d7b9023eb57a5173269f497ecb648492dd82b5d940e1e374ace300278573404b397289bf50c7db7ed0b999ee1cc71fec1f6b033877046378c2a8baa2fdea997beb15e0245415f6438c7d446a06163d06e9a72c3a362119158829283381e1b86a42fd8b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e3cd6b4caa84bd182a6c6d804c11e5d9026e09befd3c1868794f2ff647f4b44bb01a6e94374966df8babb30e724fbc585b0be0c72794c9eabcdc5e471b7ffc73ce00548e9bde2b186646b1f832710266fd900bca94fbaecf11be1e5a837ca1fe0c0494749fcac437c51ccc29ec8ac7af;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf2218f789a40658195343ca6c045cc92a843d66e7704109de127b3243b02ad5b5d71fc1d4f023095576c9ecb23fdfa8f7097fa71e498abea436ac26afd7951387aaa53fe703ef20ebbbcf93186583d6df0341299c8a40818fcedeacfc8253d558e80f17c0e67ec1d842ffd76564a4a1b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha91a34316787dc7f8dde6c7f571a98620af4edf43a8675ff9b97a0b3bc015672c2d420ea7012c0863e62f20df9b4ad6e6fbec5167d19f7c1fcff86e4bee9476e5d0ac063ce76819ae00a657bdc3263135beb0a4ae3548bf9769edfa9afa0d3547dbf5851339dd7f03f28ba0985532ec17;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18a5489c14571f9c4d6caa942118e2f0495d9359ccc3bed33a7a158eefe878672fde66d881c191203d456a0d5b91b82fa50d54dc88b2ff8f7d313255a7bd3986645467edbf77c49db355f8adfaad9b7149db40a624a05c9956e93c21ab3504fed670f680808a4ecda94c44e3a7be12a48;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf3c87207a568bb9f66757211e8e1dd37bf7e52015491aa16c4e93b10aa182a0d8519fd681c2a4310cc69fabaf314f265f64e06ba32c7cae8c3c100831202bb379cd8703cc91bf5281ce97f8969c1479a71ed3fd555cfae6b5f028d671aa67aacf851a6581864185045a5b8086c7a18c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ba27251fe3ddc46a38fe5107fea1ec58cac044e1862eca3030403e5d70b4f3c5a08fffcd1bc4cccd899180453e6e78a7370eb5fe13761c93c89ad03d0795a2348cd38dc879dcd80d8a83c58e3737fbac9821e94720ed184496233835ceae102cd7287df105e6a8ebb918ed49261d0106;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdcd5ae1bc33b92b8ac904b250d693f49da43ee9d27c6b33d259c6c9da37589ec4c644e00e2a9b0f580aa4e6942e2918adb810fead53a2d4eba76d068a3099ff57eedbb70509ea31bb1d64a0acc3758d236a6f1fdf7c9541badc80c326c0732a9e29b8d74b6753dd57a78caf11071d2485;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he52cded796945b2dc2349b9da4219473088bc7f501c1927477c466b4a838ed2d7e4a9fe7f0bf057f2c7396d4fc702ce01017af2ab855057352ebfa5202ae2e2541226b6bca8136a796e5aba78e62763d2bd8a98dadb12017cc6a7ce12c4f6cc5df995abde29cf4ddc40c13497103e569b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43c176f033df8b592d4f34e7cbbe192b65b2de2f49a272dc44d11a7f51ddfe83e554e13817d1d4c4d6dc0695e0923b480e70cfb5d82aff48b2a7e6613bfe08a3803dcf746ab22df951056524163d676e9573d21499d13dfb10a49247d8a1bada5d32985461321c0da71211b11536c11e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbd3f686a5815af8d8b7c41184a38a817ab1b7293d57008379d70ada534a351739cf88c788b834319b6b0b6e2d29f19dd0c5f0429c98ed2d7a1b614d8d4f39f0b93aeaf2408ed1b9d372e3a3fb74e665556155d9b1d77179ef9a4484e85d4594106fe694fbb11911c983f1c8ca2134954;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69a1925607056c410016ec015638371e74c0d0c43cb6d730f54a3e04c095ac9f161bceda61691b87e782a356b22d7c8f8c28f8c4078cd420c7b3da07ccfef30f321b2d9f6375c9ae23c201ab8c344fb1ae7e67166c5d790f00a743c7a488687188ab0af2030d8b5e7c4d981584891f2ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd3560326add6e03f9af521a87a4e571ae91b27a31fdbb04fbfeefd57ac7761a54dd50adfbef121d795b953a4fa5be430fef4bdf74376c757bad3ca1690ccb822cb4e3128977ebe074c8ecfefe6550b51da7351aceff0a7bfc1bfd3af1485d9079cdd9076703a246be29c60017007bd69;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h369903b92e9b542fb12d96675ea97cb1120e1ce44cd8de29d0d3b641711c57346170cd194afc04a8863a26ce74bbe0d32ec9a251cfed187eb629425d8b2e69cb674beb7dfd99e3f15c32fb8471046e00c40099254755ce206f3091953de0b329773a599cd41dad4b212b2cdb61e8b5f60;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23d8553c9b76ba0738e4821023a521fc741b6238cbb75497711298f4860e43f59837cbd6b63210ac5b7e6e38ae61b129211d0a6a7f228b38e376356bf13f97a398011a5b13d3f6d793b591ac82d8c224403abea80667c3021fa7132f7dba805fd47e6cd9e932d87411522b5cf8593385b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf12547c61340b6aa51ede92b80c37924130f6816a42757f3e56b06dae529f1307be9e2404d774636d7a82b321cf242810cf64ce1e58a253e585a0a9d2c30225591d4a8b5feecef754a224dbf01cf67cf3115894d2fe68761f0e45175af839c2fc4827d4fabfd2cd652462d67a2d650a8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca9a8a50beecfc9ac0482efb0c071643a15294e988ed91d3395d0c3e4868f9c4eb8e96f753642b8fccc559d0a44c1888db8b1925f63265f0959ed04d9c092899d78995ce20f3f63655f67a6409710b41a30b8a10677d19fea8c9d5c55696cae889b79ea9fe58720bdfc9b09ba857a7804;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff069b62662ec33001acdfe2bbe446796874b63836e5ed63575a9e405b18c631ba156fe9c8d4321ab543baf957cbf3fc10e8e6c0b4e4e9f866a36b72a043a7c1298276848769195f779b77d425b9dc5c4bed2cec50d4cabef8577e48e2ef587c2571b4203dfc13f22a43e7dfaf82dc010;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha59efa32e3051723198cd00b91203bebcfebc0a0b5187adce0f0293f8729ed1ef153097923f5f94cda09ccc2f444aa5713dc31cd8733ec27fde77e85d02beb6ce343146833f379e9acc045f4158ea4ec7f1bdbf8b5d38868945229010dea2eae82fd73ab524871204b992c980287b2ef1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bcaf0945668b32875e13130aba3f1fbb68765c5e58fd1a7ae59f1f43908c96f7d69b227df01944e25f9eb1134e4de1309ce83d0111a439d58b872a538e4eccad1604e30b7e7a0fe173ca3bf1220d7e257164279b26140e70375dbfa109fcfcfcca545e34ebadcbda89ffdaa7fd23109e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6c291cdc37160d9a2380f3bb6247f92641709dcc6ec107a783b7fc323669e3b54be1754d8715ed08ecb283349a4315fed27567fe4ae6344758124ecbd90c32f04fc3285475417e26467d95312336e4b4b1a254b553dcf30eb07104537fec9011dad51c7048559aa86ef760bd9baa843b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10650d81467ce90b7270a68f65e24bec0fc7bec753411d850b5170527be4bb4e3b5ad532f83a8394d7b5a389400838dbe12dc7bd29b98e62a9a323ab75c7e75828a3228ede3d85a03102d61196384228eea208579d0d137d7d6406e22c8d64012416098c6c726dc02ac66c7c5549b662;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71ea2cfad00e3d68665d0f5fa7dd65389a271ccaef61b4887e9187fecee168db3b6acc9c25fcf48e98d771f9dbf3da070eda060d900530c0e88ca2918edfd0bb997a07808f7c8eee715bb5c463b7207bbacaff96d645a95407ede28e4abbc8ade4af05116f2596795fea86f3c85154eba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58838ed9581b4fc494f36867471e4f499292f1ab84d10ff75b225254b0d0ba43680901371bd52477e46462c943430dbbe30b80186c828cb480d602cc47f42681541db8669a9ad0a2fc633e7e312e5b13ebb9f80daedbf5ace071a3785c620bcc6c635021ec1d5865f6d69cc3670772969;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd6381e71d4da13285afae2249ae838f0db668cac014aaa5d5ff6e8ee1c824dbced55723ab1f3293f73e7de4a52db532b60387dda10ec65173afdbae09fee8a6e118493a0e4d3b09c7b0e09b88f1372d8c0227dc5e3b13ae41d83f570aadf453fb4f6f6925c9559f536d62495ee2fa279;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h571b4db0d1be2880932c9e4df6868fd883af43c02966bfc92cfbcb13449725e027b2e98da61701febd64b3672c259471d032a5ad7299aa1d4b922e2f4375233986574a4a7116d72702f1b5151c9692b25fed6e0539aa24d444caceea4194b746faf20babe9c28d16773c1feca004ab8bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64d82960a2bd133c3d62734449a2d1b35d2748944407a37a3cb55252c9d24a3363d63d1c820428303b519c25eb951de78566cd9e868fb51469ff2265e5e8555065408f92377b283214c84f823c055593ab845dcb92a43fce152ee6217d0408e2c3800c862ea52bfa3c49dc8b196dd22ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4d3cd5c64f4399f9a8d44a6e33a560e4fcf0171ff8f3bd1114113d3e611a1f61dbc42f29a90a4fa2b031ff0af50db421b0fa6439e976c32882432d5f71cb437fe58d2e269c9876ee2f669e7c48bab7d5536b440da6b862d6f98166f1b81d4dd2620993b3c3eb4c200a8562bb991d9d96;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha05d71e4cd3b2980e2a6b4cd9b026371f60499539ea0f321a3b68a11006fdfe2c290cb549cfea3c8699832fa1b324c4e82b9f764f5f3e2e53857f994f7c50d4ea1c4129862fdd5cef8c645821b20375540a28e7dee9cb02ff4c22cbd69fbfd315bcbb7ea5b092ff060a9b15f4e6419bcb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd91b8e79a55949d3ee7a3597b07e3dd5c0dc66c68768416766f4307ef7f84722e5be79e86de4d834aaa514f7a0c113168eafb64d76248eab3936a426ef75683e82b13b62d370950be4770b89c8fe303eae7d0dc428c6f5ac5d93cae5577eec327d515d5458d9b3b2ca93bfbf51e9e573e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f232b56f832b3abedd02983d9927e032505a90c14e167e3d53b5da3aaee45a44b61a7ae61c72986994acedc186d0dd53cf9ad09c7830dba239910def2b9c06aade16ae6ac86dc5f8a85356f48042abccd58c59062f3d63346cab1c3a932d8de9ebf04732013224da421cc8b0ae80a84a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99bc54fd2049cbbde848cf649ce1c271ffc9895f43c17e9bfa8afc8ecb370c6937934d539ea4252b523a0d06fbe8acf1b2c4346f301a4fc33a11e2ad3fd924db373a89064f53dfa54dec699524e0ae5675532a7236eac9099309a6a7f70c818cff79cb5443fb25788adf5b1bf263902f2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h201d7f4931cf1ca80ecb31fbfd07805ebfe23160bb14a6a4093c08b438323e90a232d9a73fcaa1a6defd1056b365bb2abc14d969f724f3278232db91040c7e0159ecc4e77555c543d9b1fb7e0fb72c4922d632ad713163d66b1587600083cbc797cb498b95703c852e0c766377dfb969e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8140883c62c11cf4724404a45ed12ca4111d42235192ab149981c724681a135803c957b5a4034343738174fc91999b1a481530745f06ebc67270958df4c102f40348269027146cc797d6a2a8cb87b0515d478da434380a6b541f58d37d0dd8eb4f0c85fabe8db0d50637ef53758fb4c9b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he793f956be1d85ecc43aaa7acb127e41eb92aa4d0fb3788d62318eed61985363f50ebc04dbc0c43e79ee0b316bc5c03fa983dc5c5dcefad4bf09315cb484be8be267b8ae3fec570ef22757911a19f48b48f8f65b8e7b6b169721f60e59b2068f1b981a6144f75e00eaacd1e5315afa98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6215d262572256bf1d5c48a6cbb100f550e8fc85f22a573f9250da1efd1f7cdf9c5713ca2c5b52cb5b5be822e676c6c27eb219e3f09932af03bb17c3f0bc2fef9447cb5cddd34a6235d7717874b1208d4ec98c7fb1f3b552f6108ab76438e27945ade170bcf4e499dbc8a79b31bc69360;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4146776c1726fb10b081a82abb05a28f6662dd33ebb77ac0e6b69580b1769a1387e5508af93ba3b44806f4bcea900e36a807f6338baf2daaefdcf816526b98a4d6ff50ebd77840b43cdabebd98a47c22060482160a71afc136ad93a38003d2d7c3a24a35c5f1fa5b141152569ce7b8081;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7ea914aa3156d68167b8dbfb1a472d6c28b6ace2f7ad50d1d4f7de2a5ae56063acc3c92c942f8bba356238137884e439a745ec0d4ae0a3200c9c272a34c7024efbedc0273e392814eda72591f73d29fdc18b281f1376861fc794c3a6438765f8475917db54dd9797a17d448808ee5e4d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc21810795031308dfbff58d055585edd4b987e55b36c42dfe7ff20066c211236c3c7953cef3bc13b9f497efad6c89ec2a0ae14fb145664046b43c9313827ac734980c6d120a4d3379845be2c9003a618f44fab554bbc49d208580b918f5ae2bb83eb8211ed7155987d5f9a9d6c13bcb83;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99ff12a7f252ba74ada42d47bdebd460a6e29c4b8c368eca848f81078ad4dd28eeba6c94b1292cbdcf904ae46dcccdab3ecb6a6f434e6ddcc5288bc85b7318c65c347796380b7921ff22cd0c0fc2807da02fa33cfc9a0a639c925b0f9f3c40d2de74af0c716178033399e6e3e3e4d5563;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cd218a5c160e10ca4a1562e8e92752948e0bd531500c0123ef00cfdeb3f218c8d5d376aec2f213e023bda7032d879b097a3bccd0ecb9b62eb6f06fea51c13664af5fd0015da7ae05b4eb43a4caf5ba636110023e6b3f72703a1ce372a6a716f88b0aad4123676f439038f268047a8ea6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf8f4c9336ee1b5b30afa09ae788b10502af0ac5257050325bd337d5c362d64c519c1a9f4b16621d267e0cfb942e386362b91da40391bc05ce9a9a78f4558f77c19c235d4866927af2c575c03bed32161ab06919a374790573cf2d507913f92dfa63e86b80e433381e45e9b4d1e849156;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90bce22efdc0727ef527eec4117991b3986ba5c4d9421d5606e5570f933169090e5ef2e729e25258a207e171972b03f0e48f6e25e5c00864d7f2da86c685d2644955b4b3b5f7be13785456bcc67865c05d89733cea86b34659d759169d39dc7ecb708f1eb2d9fabd003affe35ea4f36e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14098551e815281b9be4cdf618624d605348943d69acb45e082dc2ce274033ea0c67ef18147614d108114f389f5b5a8be70a1a1431589300b333c18c521476bbfde569c351d6eff9b648254e706ddbc44d02cf63d2dec6c3d6d885faf4e842ae2ab8875661595e6b45b0ec657f65de770;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f8255edcf376c25eb62019d6158dab59296f7b9101a2669024f839bb4d7d2107514c905b924f9078b1ce53533b5c4f517d7d9ae6ff55e6da3ecfed412c2658fd1c2cb41c840b2a520268409ceeec92d415df561ee3e16a53acec0d688939fe10de33b976f97597a314adf6edeb9a5a30;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc49c92046fb20b9eaa277723527db583a91c311f39159bd4ea28aea4c1177cf1376b7eb55ea2711bbebcb8f17d73bd6aac950ddddae1dcc4f416a55f87bc201adf148a865f932ec5b88643dbb01aad917837ae551e9a79ffc29fb5330ee6165ebac0432e5a02c80098e5d2c2540025284;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfae13d79357f24ffa492419964d9b3c9004158378b85c20b7aa560d9a6b3f9103233b0766a8aa19c1067535aee9f8988f9c0a00a3f57de126e5f351481e036dfeda431d927bb7ab527d6a4b2ce76e088d1bcfe01f2af53ec753001e0fc89c38159fd506778304ac9315e64566588eb50;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h294097419128c02ba84d5990d287859970723592e878e9f63a5c97761d589423e0c31dbceaabaa2be18533d835caa8a74a9c791f900aced96048ef5561160c637897f07bb06fdc4bcdb7745a68995d0e8356ac6c96863bc17608c5c48eee4d1109206533422f54138fcdf1f370d9f574a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7ef67b30a65a587bf695bfb0aedd84d943c52870b929db129e75d20ce0811aa9885b75d914b1b4e574710658eb7f04057509c665ebf53ebc2cca8540a50874ba0ded7249c6db0e959ebfbd3d016905411e8bdd69965feb652e86451fd8074f216137ec749363b863b0dcf64fdd2f22cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5459028608b6b958b2e05fd7aaa78d989d10db14bce1a7e266e2cc68e2215266465122667edc97737a20a37bbe930c8f00be5dd8658d47c598189c5024860045c663b9bdcfc2df948e2caa320647f3efdc12f124711db36d9d39f25f04cec1c27ff8bcea055d9f88b2968307b23787045;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h184233d661ef1ff3affdadbc4dea567e22437f56daad9ac355de464e21b2b018af4d53aafc590e0dfc4b2aaa987e95634350aec5d7e8d278f572133edeef0a113c1a1e5c6e84ced7f6fc2f047a5c93aa269080c05fabb547f685783bf902f9b183551b914a53c038b6ac28cab14c6d1ce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee25caeec7e80b97b7444684e442161de38617672aad3fd363edeb8d0c4bef8f6264dc6b224f35a5f7733010acab785ee9548f1a58491ca5d15eed94d1fe166cd308d8b2a6eebbf3d01c6ce15af4814109aaf074897d1262a810a4d0e0ca5c8e4db2df3be3739503df6a6e0444345d21f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6956cce32758f4a2f9952fc7c29d99898744ae5979180030c9322f75422ba6545677cb12f4463616225d2f8d662c55b5c21cfbbe1c7182c018794a1b9455f2521ef7188699c75ef80b1d6311f2db00aee80834fef3051fe959decd78eb27f4afc7c87de3ee22c9406ba29d3bcae9365bd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h572d72acc9ff455aea4514190d588279de00fa6e240a908ea6c2b67e402311265ef29484f175031b2a775b80b33d46609c6a6329fc9a467f12725f7dd9bafd5635b2a8305e5bbac110d8da6ea87cf973253cd12fdfa8814a3f831aae5dea29a4792115d43a37f525cb179c5472a5c73c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5005fbc9db532fdf1250e96eaa6bcc0cc0f1311c6c050aae885594efc01a42a9133a3996d4a64d823f1b6796efd9c99bb135887031c9d49de41772537ded25b9621a6d4fee256874c411fe66d8bf3de573721fd12e52372a45ae2a8d18aa0a99080c86cf52df07da085e04ec3fb93bd6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef04974adb7e0975e0291a3998b181343b6d43021bbf1580dae440fc749a35c97b484380dc22b299b73e7c39b6631b863dc227d249a5ec862b842de34e15e6ce2a5760e181ae7fae3733d8b4f868eedc7c4a36d87aaadb6eb63ef5053a19f1110a8dc677a3709c727770cac33b62ad90;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80cf7651b53ebe2a0628d1cecc25acdaafb19e67628772170a4d32a8382f96130a8085cc4245aab6247a29b2066ae9fcdb9896da699d3efb57b0e2dbc58effc2b3b1c974dac3634809af77294284f2fe541cb84ee91a3433f1c64116224b2182f6b85d0670de7ae73ca08e09c18343eaf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6eb29183b081637988377803f1cf90163cf202e4e674d0f70e3c1cf6b84bcf773903031fb2eb3279a379b543a1691549198c5ec2102ab8d1f6123e2ec877b32d658cf28a7764c9ee14220a3cbd7ba2195e3a6db6ac24ef2a322b384c9eb2508fcfdf4cba6d70fc5c2c8373dae6fc9037e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e962175f6d0b861702030b7d8ff1adf3c76b964075d760a4664099ffe55052d4852f73ca49e0b0d1a078745daa8bf37d5c2f0b4210be28622dc77969eedf1c178b78377aa25670f40862df1141c8cb6fcbf97a55980082002eb26003233ee51f64bafd040eb11aa550543853b9f0bad1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6f0d833d3d52c86b21d6bb9e9fd5efa1c065f6775c0ac4cc2493689505e2ae60ae4f43911a45a2209fdefb719633148ff31291787ceeacb6c90b88aa443735723800b514aecde1789b1580e029c617a64fefc1bde162666a5fdfc50495f5658bd8dc3be229473eaabf48e10c228a9553;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66628630401aeffe2d2a98878519f8ead138ab0a14ad91199b8b5b5417b20e273a96a5a2fd00163f115692b7ad0b591437d500dee5c9fde4957132c309e17488508db60a5c6f2dedf14f75f1309a77040f30ed788274c8ed67186972e9757053600617e1aaf9383ce393a8a3e94b1629;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb8606b97ff6e6daa00f62ed28e4c57ba1e3adec12e25a81a017b4706ace78e7ab10fbcd00f606d42b5d8159e9b005888b3191d31674e3a2da05e9aa97c890846784ec75e4a7759d806cb78a562618e3023ff0f67f967a3aef50aff8adf1ced9b6bf6cefb27897e0e6ae85bfe804fbac5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec23ee24e8a433696d6306e2700c3472de2cb25690d3fb5cf14cc74a03ba31f0ebb619e4cf68fba1feaf87693f2dc90b08a7864b047e08a537f1916a78c640ad3ead38c11d10508105492a00d91278d7105793eaa2232cedd3e84db45c7ba3ea2028147ef5491fccc50f9d36f691af497;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22e972312e95c76042bf5ae873fa566a66ab550503ecfd7d1e523c4dbe542d43bdfd5dd89624f60d9915fffa9b1be5cf6110ca53793f7e060324619b3f1448eac263267c09a463fca10a334e59a4bb01893b130db3f6a4d700439a9d9d6de350be527ff9eb258fbb111bde9f7424b91fb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94bb715ee041fdae6b1d3cee6b5a42db0e0ef15ee861fe7cc265a4742c469647cdbcca39addf4c77b62718e8d476a1fbbcd6f36dfa81855ec09df0e4cc016a828f2d50688cb511901715d8bd687b018c5f298d62e7e380504575fd63d5e6ed48e4ecb44ca792b8befc11abe845a315cb9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h600b516a0bca980a38bce17e0396eb13284f567b1bf2e2def2584b5eb53eb1066c96f3d714e9e5675c009070fc3e9f1a62c25335d793963e0fd46ca4914bebbfafbccfe3c6187a4aa67e0ed0f4456bfb4b598f8c36327169a979ec46c3d6f058a1b4f74adcf71f630b35b92e4a98c6034;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4ef3664c66b18fc89c6bfac350a8cea1611b495b25504afd1ef8eeb7d359857b118afe0c65027a298e05b96b0b41f19ce12c5bb241fae0ca916eada47bad3c9dc9aa04c6af2e393f0e2403729cfa7ae56a4e0129dc2e4b48d15700548a016ad32688b7aad7a5976253761b0e6b62397d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4b76a5814538b43af3dd6e2eb5fca53c3eba8ad965a08c16cca1dd8db1f673e2958ab09a11c9356bea75d071d70a8558cffb04bb6358d6457ac19ef785377be07e3c906018b34881cdb701f95e7edea5924df694f487cfee89225c344ba4fab71fe42c7ff7bf422b2ef9270e1f9f4332;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7173548f01ba250c73d7bbd5faec0489b9ab911bbd945f19d0a2ca1966b76ad85efc3654220a3ffdd0f461f70da3a5d18d73bb42acfb5ed400561e1ea3ada8955b8cf4dc6a36dafa7458985454e68f67ffb7a5651dd4d501afcd0ef93f4d78fdce70f66171f8cc4a282ebf3e3675ec329;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h196db51887deb41838ac23bbd627bbf7dd946a691507c93a947328a1a51ee76daaca091bea9a7fb93c5acc8227eb2484d6035fd1a944ca7dce8cbacd14ed7666e7ecb898f94069849dd25d72346eb62ea8fe94127ffc42eac46f6a2729fe49d15dbf308beb91fbe4b80c826688d43dca7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95fe3c0665e7ca3f0eb50cdb52f65c22f9c102cc037dd53a2df6bf5d641e4a98db1ee48569345b2581ef1c0b71c38aa262a6408e1dc450f7e150186cde741e82ee4d3096c1d14c001ae7f55cbd7cee0abe3e8a0962a6fd2d32ad73c6cbf55aa01ed4d480b7a5ab033cd515565abff35d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57133d91d920bd3f242f5acc6c124251126434b0eb772c1ab51a19cf6c4ba406e3950a6e7e92522c525e1cfac6471a44d8c8afb1bc3d662fc41dfe52599886e840a3809fe88c218820a44ff8cf0a80b208f6293dd126df283ada6e54d0a989932cf1976a1f1ac25c4f582a3c9eea7fbb1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b65a367baf3d78797c84ff16e2a6301b1ca47b3be2fbafd4c8a88b1f5cbe9d192de928b45760287f9ce91e4609408e39f01cfa4d58c781052f7c1e43b96a6d87fe7c4c7b716f201eaeef3376001338b32c05b06352ace0285c0c0bc7405b40001a2916faba8036c14e0b0ed7a91a307a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c4e0ee9028598444414195fe678f2de4b5d2a03a44498b59c768b206da7243dc03b14f212bd982dd714b452997216b30c5b41f713a6adcd6590df5629f4e1c64ce10d28cd0f396fc4ea28d4e63aef00b3a04b07a8b13c23c4b4fa28f79a3b248f34ba33f5681dfa172ec3037b0878754;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87919ed48dbb948c645ffbf8a6878310ff14f17b89d8717273e161ef8b364fe58e0660e20503b9336782c3cdf38ad8aaed340f015b1c893c78b4e836c273990ba43ecb16dd806cd1afacc63ca0afd42ae2ba899b28a0e402a9a7008b204ac1f9ea5fb764167d3bb66941dd28d05b495d0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed4c9dc8f8d57f16e4493813e44a8e7e40e4b93b8fe2184d5fc9670368e3bb8654f103dccc28a7ddf73d027c4f6237277e63e8aa470086fe5db54b0f6ed1b6003fec97a39d4590f9a8678f219b03bf8ec0502e9d06aa4b5e04ed5ac8d7ce476b6e15dbfc490ec8a0998557c82efcfdf21;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d43bb3dc68125cbe7717d656c03a7a48264b815145ab67023e3c2c33c769747207ff6253f16c7925319fc79c0b96c52c3a20b6793fdca46633c44c0efb219c919a3f06dcfd6b9255086840de25e83281dfeef40851493c32c7d7d7324ad72292dc5a23fadf344a34e30fa0fc75e1c63e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfdea970dc4ba729a2514be7b517018da935439219f0d710f152daa9e9c0319e2e3463d4fe9fe4759aaad9585a560327afedf0e027819a34de60f3249b72f02e1c8de6443d633e781d18754bc2d5724fb35f5fc7a7e8509bc8a1946baa4cf77f0ff345e899bfdf007df8004434d5b4e3c6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf21c951b54ed38a42fecd2e6796826af0c7a51aa45b1433a0a962fb6d9e23cbd6b0694c5234af9a8906c6749935a4cce2c1c778da18668c1d166eb5552362a4fdd46ad0497a549dfe379fec3a4bea0b15447109fcb1bab7184c030a28f7d7fc0b35e133e74b1ca8802b123ebf4b859fd4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c2482fddfff98fb3e0127784dc21453176307401a2853ff618347a039524471910c209051ae0fa722d169553c910f7f2a7194b0bc8b0e4d98b6719e9c00b70001ee63000da254ac3daaad7672875d3c22852bd3b9daabe97d3de23b571cb39c00e7d02ba385491a919e717606b9876ca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5395a314faefcd8c3953ea3b1bc3d567639d3f4032fb0d92dd85de9933040b3f54519d77af3dc95047fdbcbeed27bd3cc5d5718b1e8cbf472140a1cd8cf2a5b19ad5e6a63cd756902740a62157b1fc5774c7a43820af3547812edcbc514c9b419abbb8b677e1344f7a054a7e2ba27f29d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbec4c5986dbe1e3e8dfcfa2b18fc840f21de7b65198e94a08dcbc9673d904722ab86e069976d0754973118f9b7d02318eb2bfe4f164369837aa5def8b63440b74e6eaf175b09def72eaa4d16e57cbc91f614cc5c6def79961266f80ef6c840edd38366551605584837ea829778b3554;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69c93e7eaff7337aa6a87d0177a24830a421119385dce478fb3895405e27575bcd1cbd927eea49a412828c55e14c4833821e96c9c0c06b69973cfde2c263068d6325255fc48f29c9eaf767c715ef62eea2d9e16855349d6b45eba59cec77081f91fe5342dc50c26680327d9d58a2fd5e7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c08700537092dc7d6a8b572521e7cc2415947264c9084191c498a3199568276ac8faa896a9767c26ad52e55dfd0e876ae6f10aef78ca7ec9a39cdddce497cd00b1a3101becdd1b87e6a67efe2f645f4ec4492be2ee706fda1c94f76562ec421a43d38f10c3a445fa94d214c1281d52a0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hafffe5114a3c316ab15f854957d23094fe4883f5f84b03c39c22cf9059acb4de7e0b7481f1bca557dda0487dc7930fb0992b133185afca3a04bfbf052bfed66bbaca16ffc6327c21b5bcd6f9cdf89d5d1f813c940f94c2b1a4470e0f0a5b5efb09ee02c927e3dc08929888a645f8ddd60;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74482fc309d5b2c3e3a6cb1e816ce38c7efd7dc4291bdb8ff35bbff2d518eb7924732fd57ebf5764cbc2bbbe418e2447550c49a0013040090a80fda7c658fadb9879513302147590653d63c510b0a4a1b7cc17b81551d3fbbecff8b9cffedbc3c4b851e1db0337c74ac5b37228f0e4984;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h611bb0e656580d9680f6350bcfad2ed957b631e4a3fbf64f82923761d2eaf2cb68abb3e936933cf0daa61059807bf28b68801129635e97a92dc9a1e1ef360d81c5c262248ac8f6393a00c11f966c9da0280a4198a80dbe503b4bebe80e616eb38a5cf0debb8fd44b93224ad27149789b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5226433b47802000d87132a2fdf07e969dc8fd625ce153be058b14b82338fb6ced5fb843aaf7f452556352b28eb4ae83faac3d86811c8a0cef8707f525397c91313eceef6e1f5bb991c786fa8211a11c2150940aaaa7a38efd2e104711ad6a18191e20e6cb0e1555b481b229f647336d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa03248f731330fa89b0b91880705a24d9dba30cf6cc52cfbbd95bf747aeb74d93dab58ab969527a3e675180e5280dd064935b8f66ad946f765f9d8cd68a76c273457d7614281e9c9cb7ff6a53ed137baad9556e3baa2b26cd8e8aac38809520964d5c23e97f5ce2ee52fae0f57ba43c5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b085c82bf4005d5d5e0f7a17b1df243e4b518258c96fa1f92a2b9584c193c5a1ce406490cb40f6a69f72310360402b13d25787eff3aa582252a6e34fab4dcc6f49720c6a307ad0f061ba61add93e7a3514c3a5e7be061f7ea0201e386d31a1b22143b3f4aa9cafdeefe9bc38f703394f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4f0cbc6c9890a9c42fac6dff102f3f232d9e572a5b00ef83be8c6ab74232ebb46dcbf0c98ac7c3c3123f4238e4c6af759e7b2f240f5dacf52beee6773075ba53d798ad3ff70ec7b2d65dd02cf0e818e410c213de1c299c4837d39677ec80cb52e776db7231470494fc4e264b987603cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h856400bc4bd6d053c74f8304d151c2ab5136ed6935ec63a4a83705216e35504079c4e1b62c852f09d2a32afbae77cabfce2595ee3ff52de156c81459a3d687daa08d8c59460d29fee02ffdba540f5b8c65d33a7530e8e1050f65e9aa91479986c385da1774d416b86043dca834e8a4f7c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22256442fef3e33c0b35bb21e840a1c7403e7782c6ff93542fd04de389856509f4269b39c55ceaf78f2ba78d463a146b13327ce87643166a4b4dde8aea2cdbe3ca892a9acc800dbcbc3f5bf289fec8828587e9503023ab917ccad51c3b69b6388a5e896eeda01029eea33e1982de501dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d6f87af83f9b826bfa50a7f471152bcc246be0d59fe8412f091730d461a4f076246b5f0d4e0d49d5203d0cb99ceff56e8dd5cb276d28a1a8ec47df993bc0285bc5baa592a0da52f578f370e7be341c8b61eb570197e17d7d5c4e25fce8eda6e3a7c10cba49730dc9cca9d30af3a73b36;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had1b0f7a576686d03644c2602a66960b304482a218d48fa269fc3cb7929a00686abdeedc0206a2650aa7ffa120461dae84f2c27c77bd4d188fe9e2c0517b62c72fe274178636ef3357b050a6ba5eff228f7f5a012f79deaf07a532b7bb8cc5a17bde3bbe8264b10a95ab7acb981c43446;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8fbc5ddcb8103eabdb95ef979ea4448e746c7b7ce58a573fe19190b8888d2caaa8f6579babfc3d272623270cc024b62e9e31d8acaecbba450417b033fd3ca3602f0e48edaf1e49bef0ed9c81e2ce55e79c1d73961dfcc8b6754e9f2930be26890e7c811c20081f8cd5ee05ce00b710c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6be45b1e33e4d5fa0db809940b4d19d0867fecd143773afaa95507942efba3b671d4cc2d828e7a9237401dc11fd39fb98a9ee6a6eebe8a43d4d5aa4349173441fe34c751ef2a3fa0f9ee1e16261014e002154806f9de42896650dff64c4a743a7508f65d0735111cc2a4963c68afdfa62;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8479695c3f8c71cae0c583528bcaae676bc632ceca92c318a414531a9e56452bc8e2c9569025ab40e36cdefb0c500e177f8ad92c62c5086ad7e9c727140cd451bb4431a90de4a129ca991ace734f96810ccd936561fa5d8d28a306fe5e487048982ee240d27781d544e1e2b4616d2ec74;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d42c43c0cf4894b0250bacdf853c65d8a862dba96b95928bea74ece952f0b933fc1154ea2305279f996dec2b6840db51fba76db2310b998cc41d4411b33f2bb2e45a5d765b6c3462f2643fc9280a7e7117a06e8260fc724ea3dcaa57c11ba66aad11c1c61ff14d3e92170cbcc5be9f29;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha70c0ef743c62aba7fd30755857b9df68eb20c6993a97ad6c595f46bf95b95b388089647fdc5f505afed189ab1145b08b60c52b78e5e3e9f314b29c1af6f72d3bd69235b4bb0d51e455b2f9f85825929987a2d5917b2a7204181288a8163e3dc523bbc7327412d38211d5a20f6f6806c7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he094ca4d6ebfd7e670cff9750f50bc0119eacb6aea494103493c895e4cb03a3dbf561b51c5245ab930004830fd5008484604a6da86927d7d4200d1d29b1ac465707ed451fca5857e737916252adc0057e97f51ed0181d67c97dcb399bc80f07d99437248d879c4cab9dd0ca460f71981e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5068d509bdb9faa3824f3d294ad6930ce52976f5d5b981a996bbc9fc4e3f67a244cbfd7a40861fce9d0a968d57e7f7b6d6844fab4f026205658c8378119f066772bd8471c6d6f9a3f4391fab9a1d3cb7d0c4407a6b1c296e0d55a46ae2e1bc53cb9744b62b66b1b4fdb16bdfe47414344;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfce76c4bd7ba6e092fc78becea3fefdccb5ef62aee61a3347cba83e3da237c0657aea913fae2c1e9b045069a7ec807ef4f5b1deb6504403dce3e4922cb8753b551a22555fca867df3e8c72d5de37b002af70cf8a13e53b6f9d45e64f12c8d1df72d0a1c7fca54df0c3c663d9eb298b93;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4703ccf5ab8ae3b8b69fa5795e1db99184f9f54e855188cdb9011c62f4189699b5ff55c154d54a041ced192caec69b8ceb0cb67998ac594cef9e2c812e273f7d9e06c95c097c29e0d57ed64c31a939ee9dcd06437156cc818b348d2fe69cbd91b433e94d2b76c545663c0fb8cde43e5ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54513c77c74af4abead09a31bfa179abe6954949042dc75ebffe66ad799639b27bb29abd891159ae0f3317e449b3a55688b75098d4dc67165645fc1e21f03e83d304a65656993eb25702f58e2ceb81738ce421e899fbc617d8badee608f667a78ad5368e8127cc42229d3f39d97803d5a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h494971725dd0a073075ba65956389887eee262761d6a20f435df9272b5337ea5227635b31458a068835f06b5a7310ffa40d9ba3aaefae77de481fc4275f2e8be939ae37771f0224df3de98fa944ec6054cc2c658801c7239de89b07ed5d13d170f6a5eb8ab6a61c7df85624327c101d53;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a863b24a0cc131cafeedf7e2a748cdc82276b6dd7934bddf2c580a719452db856e46edac0b639d52b6d5917de33f471215d53f8256c1c176a8e84eded1edbb3de41dd92c3a9ed1d2cffc2ff74f789591683363f560277e680912832441f00d6df1db9f3bbeff7a89398cb651c02846b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd472a779cbd3fff71c1e11c3cd8b8813b95d1e26d4e0730a8e4c3d35a38de2cb221d281d54d40f2b053fc217b2fa0348ad6b63fcf74f5a21f111edca76d584d861386d544c3c281e0a35c7f2f25d336a04242761cabb6d45ddaadf0ec2fee7abbd4a8236f1bd9f7aed618db212f8df95;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7f2ab94e4602dd44f686c735a1c069430c75fc329edd30555d0c5feb8e6bf9d536b655385c9f75b8d8df7074763b3684062324d91960ca9c457d5e5f26839ffcf57064907f9514c7baeea9fca6ba732315711c728fbba12b713cb7707c359d836278022a769cfe0d7460207696db6a54;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he99ed2c9c74f6bc38ad7be42056e8e26be44102da912a96327cf3ce2c586f3ec54aea648d92b66d3bb9e809bdb91037f9212d692ce374524b56d9a89e51da39c3ff019d66ac65480377dbb5247a9b347c8905368a7d30caac9b8b694f973813a5ca553db6582a91480bb5b1937b593962;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb40802e910f5e9ffdc6dcf1bacd657ea2933e7664737f8bb3b62f4ec745b0a699f17a9e9baacac8852f67af9a6d18a3ac69ac18f9dc1b1980aeede9368b13b702d1c88a057b4f85bfe91eaf2a02ffb955b50c0a48a040d03e91ec3245188887c3f71dd6691b0c22e5db3f25ddd0d0ddd1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d81cf9f7e17f80d09b63a35d27f4e1298cdfe205350a1bafd1e7d499a8220f461e299902d88acb3b97ba6c77f468472cff11bca687b92ae026c7e91a8bb6928e55dbbcaf49a2aee3d2dfa0c649ea7849ecec6a815cba37588560f4350cee233296a08b1130ec03d2f5a0a8749a902a0c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43f23ea77ff01f7ddbc42ed07cbd6b542453ca1212e244a5cccc6464e94f9efcb5d7dc57e5e71e5fbcf2aa039e641679ea7185bb23cbebc5f90b3f84c7b7fbb922ca31e2fcc150d16b782ee62acac69c99f8057219bfea1c3c9e05b74c8339a2713e76cdbf74424cabddff3d7a1ed155f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he055328ef265ac0e745e8991ad7f892e385be20afd34e28b3f888beb8bd8bf432973a8c620c2d03e5d416b2f436b96e51bff13d3b1897183a796dfc32dd26ed65d47ba675723588a98beb8caf366ffadb7c19b3174d0e21914b710e24900dcef6b235c4b16f10f1c0b5ce167ed9f19035;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95c59c6afe3df8f2602e63359d8643d732ac7e5edc7c67c068e2529e484798b9971bc84fd2e92d9608183c1bdab81672c17ce9460321eebaadc382c0f20e8a53f3cf77beda77dfa20ccad05a66c2a3a5d6c259095beea797f9c7a7bf0b6505b60deccbeb872502bd8f061929790cc5d05;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3d5f964f66c57f5d38aa4eb89d1347c9b27470d8afa89fc93ed7d427216ca69830bb7cd3980e8684fba33bc1fe5d64383476735aab1d8806cb3357fe532cfacb71ff728a42c718cae95566b0d15ae65be83ca81f0a47c0380a691ffadedae88f128dd5be12c7f9bad3ca00fdfa711145;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd5799ae441b62c81a74187f947f2702cbd1dfb4bf148b0d1c6fe4879a180c6731e690a2ff0061b4fe8168ed9cb7eaf142962bca53bf276c663cf287ba175a6a7babae6eb9aaac7273de8413ec1ab1440093178e8d1e801e88cc6a168a72671702b24115dda713a5c21532a33e54a731;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h447529dccbe3e525c071a8bac91fd57eadf82896f71c740efb57824a778d82470730a810be0618c0ca16b9105dbc555d2b76a7956cc576b6c6c8fce17cee57a5772b887a5a7ed2185af34d247cf048f90b79590ff238950fa33f891e7ea1db5b5f6ed35560c8372587e58cc99516d3c51;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hefabd2f21bd4a2179b6eff3bbadb0398a3872764a1d93d7d2518561184e2f24675f51c5f285deeee0767f2e5eca92bc026cf70862d86b29d3295b3dd6c5f0e5fae0f2180f5afce0ab16bfb853568506bd0fb333fe43c45eb42ab126117d766b38edccb482aaea6b6dea937f6c5305d530;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89a99a4df24cda85c2498aa35b52c4687cbd6271796f270b21d642d80bbb56ef4c13068af03767282b295233636b379064303f91c008bcab5530c34b03139395702846e947304ac2e9b7320d98cc1f3b169927efefecda6576a2b9ac3ea42a2124294156f0cf59dee8809097a7209caf2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed62903170c2b202fedc687d1d96601d8efb36308bdf28d897784e7977375c77014d54f1bf7f619a0b6cd40be04219953805984def197b9c8f23962b56cbc4322988d0f9f36b168afd7ec5410d6460f4c1c8f18742e7b266f081b0cd8b360b44c5e6e5b09f0740d11b2b13f573776b3f7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfb69c27007faba171575b14083329de8e9a32f4f3671b701a4bf3cca7dfaed61a5705176c6b8f9862f7c5d376b93cc40a2586d93f47951379859992d2038aa2cd4df39fa87ba07e3dbb1d8741ef52191733201bd1a5b6437778e1c368c2e83adb7e84b78cb9b3317a10feaa615732b9d;
        #1
        $finish();
    end
endmodule
