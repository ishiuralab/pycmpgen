module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [18:0] src20;
    reg [17:0] src21;
    reg [16:0] src22;
    reg [15:0] src23;
    reg [14:0] src24;
    reg [13:0] src25;
    reg [12:0] src26;
    reg [11:0] src27;
    reg [10:0] src28;
    reg [9:0] src29;
    reg [8:0] src30;
    reg [7:0] src31;
    reg [6:0] src32;
    reg [5:0] src33;
    reg [4:0] src34;
    reg [3:0] src35;
    reg [2:0] src36;
    reg [1:0] src37;
    reg [0:0] src38;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [39:0] srcsum;
    wire [39:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3])<<35) + ((src36[0] + src36[1] + src36[2])<<36) + ((src37[0] + src37[1])<<37) + ((src38[0])<<38);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hceb2c8dce775de0f877ec3d2b1a96f3c7cb575a8d1c36450162dad9474edc891c14daca8ec53a06ec8fd114bbd397b82c89d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce1e0eeb127a730997cb6c909f07c6872a5567220e10659826082f870f4585647136d9e0633ad285b7278059b7dc31b6afc9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bc50abfff19cdb027c4793a38014e8f7bf1f16d42999b20ab77717d49579a8ff6e1a60dbd8b3572b1431f1b21aececf351f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha240a8aad50b18c6a60470e45ecb3ee08cf168f331f36dc536ace08f22bdfb3e48d733deeb1ee1322a90b6af69a89e20bbc9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28642c9f7e8e01b9db5d141ef925678fb63398064384e0e8a673969403a109400c784c82453207bff3f177842fc14599bcc7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a08e91bedd235b7657519a43f46f271812d0b78b41d3821b87998fd8ece2ad6c5204db15f64b78fa6b1cbe1894ed7db454f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdaeef60394678a21986e360941241c5aecbbfa0e7a0be2c1f1bd09b2ea9826efbd98daca727f5cf2c8ec4bc6c7ff2f703eed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63d98a3b931cc5387265d9424e805a4c3183b2ea0dc585e69ec9c18e9df0aa89db00f0c9c440523a3ad5732e524a179755be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdad3865bd7b139cf6c1c2729049a7945f8ce2335ee0cadd324613280fbd299d607db0d9efe742364e649304246a182f50efb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff5a264e2a76698eca53e079701671e348ef11bdfcca760bd38eed3bad4d39f9d5750cbbae24eae755125fca8ee82d2b35e8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82c13c6aec2bdebdb5fb85471d15dcb5c37f8974fa4eaf76ba14e1d130a7a0d0e510f54348293560bbc17c93b5521588b300;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bbf1bf21db56e4fa38cfa1060885ef50f447c4ab3437faa924d839e1b3111a32b0555afbd3fdd1cc16ff05648b888a55d1a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20b0140e679e36454cad72af47cecb5b3932e263efe5ab8398c826061061d75b4687aa98af2d133a2ba31b3ffb9170a8a3b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3260dd8a725edeca38e12e7921a876afb285e68113cb2cd64893bc2843c2c30b06decac53ae3b0d9330455a5aa97745d6863;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f5366876493ac7c0c34905e9d17fe9e74b5b0c94fbfea8f51d28c5ec647339d64e2df6975cc6b1e5e14cd492293644074c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51bb63565518c83ac8bd656de90bd8022c6eabcceb8f786cb9d20d175fd9ebf0ff53d74ef19f0168598458ed82f606d6942;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1b3a259cfa896009e74b2e1e52ede73d31a1b7a1aa216b23872de6b2d9649566c61d5b7093c47675d4c64778108e4616a74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2233cdaf4c806c887f02ce1e61ce01a126fb0385217b57fe42a095d0e16fa98a20b3323825055b17cd7add49a42b2708ffe2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he55e5cf76f3835c76c0c8f1ea3cbd44569692116489d2f47617c2ce8f1d7e90a08d08f14c4c2650d9d2113d6b9613db14fdd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f171d21e2553c78c28aaea853ddbf4b69265b45a6e7526018e1ebfd2bdb18b42c0124b736a74bd7513982e50023cc1f1a41;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7ed736e26d7e6f154c1c03447ff6d5f820f079f8cbde0294bbf219980d3286200e0753546a33d96efe63351ea09e24163c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa910988b1204baf73459dece7a3e0d8ff5311b486f50bd7927d0ce16e4e04b643d2fcc3e0ba877052d88647c4053ec4e708;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44378076f1f38af5d72fb9e25d518c7171d4b7f8550bc547fcb4ecfe4f5d39bcd8f063045c4bc7e8582e559eb022117f4e48;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c7fca5150a5974eb9741029561fa61c1d6a4bebb8136b8700a0a2127a31d808673ee069a4bc996e826ed8a52df237949917;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf63025868f8b49b7e5ac3dd194cade9c743e21b634f2ce868edd0c6ce61a9349f625af2571379193cdeff0918f734df2aeb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdac6aa27e801e44f1ee82bba62ba6e6ff5577612d7b5fb78969b2bf55119de0b0e8659b0be8682f8bd0f89db51aade90d16;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb4ce2e900364244418f2d75fc20a688bacb54d465ea647b5e7ceb6e52e5012170e4898e82afc25bb69bb65e64752706c93d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcfd10a548450d23202052a13bc2b70f733d2abdfb7c7b003288cee6988387e855bfb366e79c92b2e469a824274cfb5f5aac6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31799d5d0b9664738e1fd4460ae74fb8576961ca846dde1b4c8a230cfb1d3485a77db5aa186bf36ae1859b4682872f5505b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha884d8f0a880059964b06d82e4b513f7293b5e798dd0cd5cedaa890abb00b7ab85c4ebff9a1316addae9219daf5668053513;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7e68d71a5938079cdfc3b54c915113490070cad1c40e536b693e502c6e795c3232a17f28fbf5084cdeb6d7ecbfe6b6832eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8545084426220d533446389cd4b8a730e319e81ce7d9d4f355cf1db939d50c0db2f084c9b307b56216f280b80d195122ec18;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15cad53bdd1818d3f43f764a489b36ad8d86f0ed23d53495c2758af50e109236c6a459bd1b2ebb8fd4f4ab385e326fd588e8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb6f07592cd5d464671b34639c6b13d164ccbc12fe4a8473efad575c2f3513f0fcda6d07df6f8f15ab7cbf0abb46ac6294d7a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22a96333877d34477d0c842bdc02973c8784ad292b938d44546c894ff2f3348e29cb030ce79ff50b05cc25cd71962f03ac3b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb40d4092397c7b3e9c8a57c8fa32e440da32904a97f15550c76918b77d04a4609cdf3eba57ff676fd4a3631c4529680bef5e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd916a4df4c65cc7838853eb4d7e1403844b12c3010ab3dfdf478720a6246617e26b97923f12bbbed2e8edcb886e86c1cd78;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff076e3b1de56f52868a6f08a2a2e032870c969b9bdbdce6503b55781567517ccc2e766dbc2c746b63832334505d0de92cc8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbae5858789110cb8c3760144bd0384c448ceda789ad488652e09064bd5005186040576fbe930c010d560919e9fa94d8e48f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90e4d56aace6e83997fba921a6ca888b8bb80db1b6f74194af511137e76e0f7b752326a81d919a464648b3475510209cfb23;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he950c2ee924fb69ac6ae6e141adae9759426b37d42d1cf8410f9871d5bf94ad437e8c8a2fcba0886e8f0be29b921e26fd97d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d7e5b1b4aaa6e03c22a6cc3fa634aa74ff39aa1cbd0760952dde4e20418aeded34c47e5074e8ddbbaec65341ed7f3a8f856;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e66154273e82127ebbedf29fcea45054e7965789ddd7960fa3d2c0a789033a06740a192f5b78af7a0112cc8e0f65bda2c21;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8953fb6c97b2950243be682690760b66f6c1e1adeac6415e5014d65c53aa896180173c47cdeb5c4a37d01a14e9fb02f7497f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24df8e6c46294869dd54f74fcc0ff5a0e5bf889f63c9706ec51ea34cba77a3b3226e64aa43c71a6a9a5aceb63ac1c306d85b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13f57c92fe1f7f8f79e28d15f50dd430a1e6c6ed49bb2388d919fcaefd7cc162e8e258eb0e974b244d4b7c0b3b3da6a3dc57;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h896763c0e0e1dde8e3772730dda73f72e215fa168722d57cd2e66be8e9aa2fe9a237f826ef13254d3ba0b221b01905e5853a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h944bbdd775aa48bda7ed207e00de90eca33a1afae7869057f864055f0c3b4ff4328798df9d022b45a870982dab23adde5f2b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b67cbc2254693bd83ca28b0d77b7e0181b744759ad2db4c3c4a63062950330b23da973d85a3d8e60ba88541b4b41a151594;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37aa014ad15a64a22aa2194cc98fa553620f518a6558c9f302864882025a06b2be7c488ef90a2a4728c78cbe167f6015f617;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ce20fec10723c07aaa037a6942b3ce83c189ce692e2affb95493ad87f3d082101e22b03ec36d428f3af89eb1a09b5787a4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76c9a4cfed2abfdda7b6caeff1bc8c5ff63aac3f3aa1c9e177c6de2802f2f6808e92e1613891378bd9adbc2ae298deee2291;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h716c63b6720b44d438c3923ea38d524b34cc65ecdd2717a5285fd2e8681a062e21a90604becd14028fe1c9501a4a073c4c65;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc860ce81b66b519650081a53b6f74db56a71122b74158f8b5ba5bc90385106e0953c8e84db6a9b67b875f0b67cf3d378aaa0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf09f93a89b98dd390278f490103edf31650fbc1be16ce83e2f415b0912539c2a3246bf07d7b1ae74b16fa258496939b1495c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c57ff95e6285e80f29df81c122a9feb39e487fd626d2582b560024aa6a4c894b2229fd40bf110f6b3d26907bcee94558477;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3422a2c21f8b381b36de6a4a265009ab638f72dc15282eaa7d585d98cd9357c21d05bb46d3372d9999e6b027fb6c5b8a4dc9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he434684679950f51a66425487657a38314994ffbc53aa36e5592b238565a1dfcc36cf14405cba7ddcf2e0926ed04d562115a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b92c1d8b7714edc452f2f4a784007f4f8c3fd55c31fa54eb509628acec72af89031f8d574cad1c51a1eb2921662da2f7281;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h473f8e856d837357abedf3179ee0c8450a6919c098d3ec8cb57b5ac3360c8e1f42007323885095fd920a730891fd51edcf46;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h793eeeb496e63c9d371c014db36afe271a939827d6c1b288d1eea5b630b89e0563a463b8f5b224a6007fd966d9a74e14c37c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52edfedfeccca3cec67323683fa8964161d93a209b93191280f71db89bb607ace914fc14f798302d4ff8269fdf29577d9bb9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd01738d7f3375e29139e2fa22d7dd9225650342448cbcc725dc8aab8cd43ebab8ce6bedf8d8c717ffc62e4aa504863bcf6be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4df8325dd47f2b571d63bad113869b2dcd74efcb492c6bdb8245c82effffa59228702075863f7d445331ab0c049a3b7de543;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7aa194c855f7a40a7a7af5498199de86e372647f9da4527289ca904a8f5b836de908f9090958f2c47f46acbda35679328273;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd191deb37d489f70a67b6328c124c488ca74b3561011b2dfcca3f05658081222cf87d19896b21ac94676afd253f343b488df;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7690691981e5935c9d95ad0e1f3887800bd5dfea74b2c7caf1a9b581dda973eec65f0a4e504bd70f5b10e373de7ef04731ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc53f1f1f9176451df33fcc179b54c47b02984b159b0e57a4cb7e5df6fa31c00bf6aedbaf7b95b42fd1e9e73148bed65cc01b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2363938d4b848f1c1738002b5a1c7e4aff96225c1119f01940a20881e1ae0bc8714cbe957f6edc2e8d2ce49ba212924d27d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd705f6b790aa81ed1da49b1764d46f3d6bb5942feaf6bf2f4199f3577e3d25ae03762f425bf316b8b8c5d4db11cc374b526a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2beb498646a6591dd814d47301fe977d6f5e77e7583c7b990b677ba57a6ca784e7c2a9895ce770039c094e628be549f77b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a2c0f9f7d7f9096e4fa985e064a723c0974b20797841461ef9401905a4529999cdac71d394e7576038850aa69ff9e920f2e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc115a207319927b62e1e149d1092a3afd4abf41060e45357a21869f18a0b889ba54c980e9ba25c29444586f882ce8aa9e7a9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h532c669c870a7ff6a95bf253422eb907e05c6f87618dc144b20916d3637c957354e6155dfa293cd74a05bb5bf695c3664ca1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe1b8bfc54f9c98febaf1b22c27ce2e9b7ad85257f19f8cd7bf91eeb72963f24a25ab2e51df4db6a109d5b93e663167f3d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1634df864430491d828133b7e54f535e31521ce0ae6fa160507a8e822bb6424d68b001018db67aa2d93b23a37340480f50ed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2012392e587a4a731a245ac50ae05d2dbc7e155864a8103826801d3a07f067cd4ffbf33449121e0f545459ffa0d105a97a68;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58ed40df2c6370fa7e3561df3587499a68951c3dc26d6c11ff2ed4daae3a65978c37b2513447ad6f9726e4bdce20a4f54e24;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ea717697303d69f18c7ca0b84e8cbe355eef53877eb2d03d433450e82b581bc7611d037525bb301c696edecbc9c526a38ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h227243395dae105f72067f50842fee974531203d93472cf44c6cce16a95f96b5ebe6fa36c62a19ef8e0eff9df00547f686cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h550bae6d2f0cd8bb8c8051d3aa35b59e89247468934bcae66431b1988d58ddbba2847d32b7cdd14c47d4a5f95679d12572bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he53b3d685852284693b5e6aa6fc7c7fc515bf76df01160a9e8572901d58be3ad7d34aa41d511ee21b4502114d277ddd9843a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f3b2bf306eb7ba39571a08c29b0b6d67dfb848fd2b50af565d982bb91678f5e8e569a41fedec6e0ca0a5d208aca4ce0b9b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he93f5a9d01c0dd186803051f635c74e85fdece8d8a40ea210e9bc25a0c4238279780c8cc35963312446c45a142a0fffc7750;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h275f29988bf979fade82e7fb8cd5506f468eb4eb0af5b38f6ee1bf988389e856070bbe97f2418cd4e4634bb8efeca7a69323;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13598c69ea49ab250a734e68e7179d21fb6fddaccac972485ec2dc6ca2f69e5ea28d620a4b29457f294184574124d35972c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d2a92a487f5b1e8ac02f5ed9fbf7496c9b6bc17200afdc96e8c93cc0c48e62ecc52ea81f1c0841dfdd434a58c1c802e312a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f8adfe9fbe583bd8c862ca6a68453b22b11313b268725676f7e3f4e0623efd4fcd646183fa2123f5f05c0ec2f8e312fae4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h893d7e49026b28aa65de8ecf58b3f2bd88418ab6210a32bd67ab0ab8e6689b9d72b95c6ff627ec5519e1ebd72b69297c0a4a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28d6e0c30cebe0e7103421208e223725f3dcb930b5960d43b34e65379a0095a49e0665c537fdc4caa47dccbc3262d287dd20;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h415dd0004c66a365cd3d38d46558b890df16d280439929a4b435727872d0f520cf16a7995ceb4fbe767760463a3853fdc385;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd2d52d953bbff75f63b5776a43b0171cb65b52b2377d57e5e7245378598dce103f7cb996f5d38464277dc8dbeb9a4b4ff8e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1ae6435fe4e21e278c719563729d5f1da7158c238248d56629be469bc4e2dcd98373897b184b40e1c286d699465ee8ae802;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82b3c50e779922f07cb251eb5c6b11385b9c25dcaa658c3dc3be254187de3ad990508345677212215421b5e5f5901e118bf0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he00e378806ca3954a917fcc2bf724aa3e1425048104fb0d5a88aa5de60e1c2cbe1c1587d6651e2fc144eb9b39449509a4e0f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93c209404a5490ed1818c8c1098faafa3ff1d3eea4af07a637cc44b40153d405399ced54219a874f8c5984585dc2de1dad08;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6c7e4e0a83dbe9c56d68d9b0571bb99d85d22c0162859354b8747798fc42d907a56841251d1743b7728aee7d05ea98bf5d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd80b0d089dee46d4781e39e71943dfc2fe545f016b9765a9f26063e1af017ecfc1ae16df214a082e47a5ca647fdcfb110bec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h477ade125759059e922168dd163748e0d0a4a51bc0994f2b52b35ad7a69010a9ef93d8ae855dc031b3d74f6fead7f0f7f2cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h39af3a99dc64faef3dae38ce83874ecc922f6e301288e58d6542015a38a83b0edb159873862be6ac0cd275f99ad1d9aff5ae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2dc8ca4a818160c5f591e37baab7f3b65627ef0af7a94c3dfdd465b54c7a83c08d5ff3a734aa32418a2b5e0bcfe2d0a9010d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf43fbf1d9dacefe069499b40a8efe34b4824f5e0144c2dddef23767d486c42365d1706c01f47d59fa7b6a1f6c331685a118e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31aad952a3485488baa189070a5520fc61379dfff8d8170c6fa2080af12cc5ca4c445823c0fb32e736990a8ce9bba7fde025;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6f6501e58f0e3dfb6769aa8d632cb65c468169bb1f039a08b38ab23c07fbc5c9de196d87765df6445e62cbbcd39feece977;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h349918f991c52cabed356b0654ac5bb7abe83ee34a20ba161e0ac77e39571a5645bc18eaeec85d5f901c2951ab911598f8c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7ea38bae2d3399cce3517b6054b46a091b13edc5934e40057ef817d500b53ce86d919f3f1feada1a4fbe655c606afa918b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6bb2f42a312c966c70bc6a97ccb1c2051774bcceed601d72f51cd6c2eb614b4c3bedd57fb683a40206167d7b6687ce79051a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4ba2a67a71be43d1c313470cb0e09daf8f88e19178e82214c004ada89b43fd78e1a5d1db2bed31b9e6df880c95e403b36ab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h963adac00a70a49a3eca9a730b414c081ebdaaabb4b167c744841d323e6a1793f965bca2bc4e31c563856eb8babba6068d4f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h110f8ec16ad92af215e4704ef6331453adec06565d7175cfb0ca5ecbf9aa3b12c47cfb301fe1c61af97876ee5389854a6cf1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha65be9ef5f3804e5c54d63101ed2be4619a703962a1c29f195b2442112d6e98727d9b9ad9768ca5ce724065dac8f403de1e9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fc9c9582782827c6382c338cace5253c753f6ccf11d998950a6aca82358881390d0b6d1faf86170771f9046def4e1fc8084;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4d9ad6d05f83c7523dc89e1c6c05150c45d54f16a26b7d390ea4395c070ababc80a16d13b0e279f0e16a6e731b80c8f4081;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h79c73af78d95adb9fae7e484e388cf88775d7f150a4eb9a531cd72a81213e3ced66325c5014297f5e3fd45ea9fef79435e35;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcecf1794c181310551f2a55c4b81f6f203d4da2c00adf22bef021ceb4efe6af914b590427b5be4fb09f685a37b9a74cf8dd9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h369c44f89eb4a32da3b43662a99b792f621d358714897c907a04b06db2a028a86c0ce383af01deae20720420d32405c7ec46;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd8c3d54e281b99a68217183f4baff2b6d6503e64dad8ce13d24ad05789b52dfe24614bafc8c7c170f85197a061f0e88c312;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1aff2273e89ef2d216a1aa450e3776d33547d722d6c16d5b0dcd250ddb86fe1e23ba8978d0e7ecad41482bbeeee9e265a6e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b80ff6819be2bac104856fd5eefa6964d1b09bf9a1c9c967a81418555c266ad634c02523c76bc03fb7898732ef045beb9bf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbab607990117c9421859e58438457d6ef5f06e48b54b90cdaba6f59d8f767178ed1f4d6c435635e877828d1e1f4952f4ca16;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf8e3cb667247d3e90609e644d9e9306d283e2706f9669b3903e0d308a6525bbb526f6d968cbe9a3fbe8116636cd1639176d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99c7a5546020fa57eb68ddc947ece0250b4a971dd24bbbf29071da65cd28ce2d41f13564b005a936f4df90dcf5a5b119844b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77ad5e807c51a4d235d46b939157495fb497c33e4060de7522e4fb0ad91df330e86ed2cc07fa4d75cbd0dc6b180c159f7ed7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c4a321a72b5f79cb81d5edf1758d69fa89d9e4fb923a0804ac7bf8aa694fe3d44b36ff05aa122ae517394faeadd94ad639d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9fe05b8c4b0de48408c6353b3db4b34488e38d2f4c81a394e8aea91f796fd8de2c26bfd773233015bf29901483730e68ed3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h732ae73c200059d67506c1d7639e50857e556320bbb5595125f24fa2778a8825fbbd0fdba96e88e005970505bd3d46a320c4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha985ee54a5364eb80bada7d7175700d099b1d94b144207280ed14033056ff17af2c2ae536120c94589d1089170be8ad69165;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ba8586d4c2f2104bb6e5a77c91d157ddb761071cf9d51dd05ed329f182f80d686126da546fdb297fbc755072bc69e3860fd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69c257cb2468b648a799913d84bcdc803ea00fb1f16669ae4425551b8a88a4931b367d7cfc5dc4ee9fa905755152a7bb538;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8775680675327f5267681a7b49f66eb02993697bce5c23ca0f2623a5f71febcbdabc09aa3d88627dfec069911964eeec289;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86e33b8377e47df0f409e94b02f0382ee0e654900dad51b710b696d1704b072e15360fd9baf0086a572fbddcdc3b40a90be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c0cd7125e1dc473ea18e3e6ef1f7e3bf4a8392d841200a0b9d3ebb8e3db08af87fba2a2ee417bc365b06b4535be637224c4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd6a70845417c8a669e4f0a9d271395b65fc26937212726b76b42cfca36540e7fafa00d92a196dc1e404f9470dda9a89ae46;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed20c17135d5a645256c5b8b76257e80a2abb2e09df0642c76ae5fc414a5b1e06116cd71776815a4dba17e83a098e4d6c4ca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62a9d7a1de41163b9c045dd40b6e17aa52732b731b0cc7e61e912517cde9598e542649ad3124d25a5f219d116a5ed602f8b7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h778ab1d18dd35c1827800309716be7513edf877a8f46073cd95b7fd2bbd597b60d46c8562505f76b92fe92628054d6c6d25;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd5f3c46a23eb037ef25082ad78987c54aefcf1e29c38e6ace31cd0778eb14eaee8230ae32bba8b30bc903ca6b670dd47dd0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h636f0275c110bc5125103fc498b6bd69388a96732b6c8bcd66fc2edc149b8aa7cf0bf6cd8b44ce5b6592db1ba483664fb6ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h791f31215b54d08f6eb0444db9067b31b5e3b8e1133f281f8560384f846fef37d7bf55794ba887a1be84bfdde63e4e53196e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h649085751607d395966302685cd659726deb4230eacfb26924485c1271bb88e4435154e32d73671f674a742795cab2bf7d02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7acaf52c6a290ebdebef818efec32db5093f32729ecd5257bab025a5271245abd39572cea26db0ef23eb35e0e6ca1b8dda9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89175ce7b733b700207d15705d4163102a0e686fbdc460a38382340e09390bd706105ffd8c875e499b4c87bfffe5bf07d51c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha875a2e82aea9e9574d69a3927cd85c49adcd729ba324c1e5cb5ef9daf2f3f79939f283aee1ebd233cb0980d9154bb9f8257;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb818478d7b7a3dfc816f05634a4a21be3b4f975dfe6e581894527e70af44d04f4ffb0b3684a5807671735f5cff43f9732265;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8567b0a3026b0b2b2e20f1d62e95d19c8433c0cc9acf460b2ea975a1df4c691b261063460b58e26b1b7af187b374b7c8997;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h702f9f65bcd4d7cd27bec6cb3809fff51ce59d37e94bba4aa732eb335fdbb8d11742d29f012ecfa09b2c5fea25b0c2d9be04;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb9baa5de7a1e9733da30efca2b355555f53a99b12658e12bf8a3461c4e01cbb72c23d921a22dd251747094b34cd5f97994fd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0c22a259f4a97f958e05cd6def6631e95ff3b4bd949edffd11bb8b781f1a9cd14800535a38ecc00aaa8fd1be9e2085c2113;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2dc8f3371b504c7ee945e095944ec0d65304d1f7f2ee0dd56383aebe9f217f94848b6c1964421cb8fad501c0f3b38b4620e7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6963bdbefe5719e2a5366e0d888e54d20ab78ff7b6df42c6d42b699255bafc07308f4f10d82d13d1388f74ce01eaf60e21a0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3877777632909030184d9e0b9516b982cee1f19463ad4f8a1f92f299bdc4707401f635882e3ef78445a8ccfcc7d6b90ac276;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0e7fbbd0bb2e88da6fb9b7cbe0aaea67337268ffd8275e0674c28ba875703c066fe4f4189258be1216076c46649788ea887;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2edd4f0b6557e0ac0bcabc87326525ff2445692466834a294ed01ea075299580583d450f38e3c8c4f8b8257701c1dddef345;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf357229c6fdde8f618b369abc23b8f682e0f966987e7434aa06953ab543d6af18e0ff17a96dd42ff195e0ed91e748067349;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h184f9150d62b8ad9d709f2ad2a912a0afef8c6b2f44f7e865246bb503ad0c5e6f5ee0b035f1109b4494a043504b345efb94e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2333c85d4a6f3f3fa2a2851fff72f7d06e02a31d939f6e910830f2cfdbc93c526b8d9c33d87668e440fd1b0dd49595d3f4d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2ef41ebb89f70e78b4f00973bcb8e34290fe251bb4fb92e7870b2869c65912b3441a59a71f5734f71a85a6b843deeaa0726;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcab508c341be34dcb54a8b0f9a79695dbf598461c7a54db33c47f83d24e21957d52133af7e90afc3f8a6cb5421c79aba8fc2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha63fda086ae1787dee2d324ac31ef5d53d9fbe40330b82cbf16b0c131c1b55fe38a1600f062fa10a0ad424e09e63809d0dda;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bc64544356aee0cac564dedbdb26b95d2a48e98dd16d3709f6b507bc95a82e065b6a67a22fcd4dbed37128138fa0e5b75f4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h874e847f2a80f7b655e4e1844cf39bb853e932998dac55004459f7d584d674cdf6cfaf8e16fffbd1160174a65663bc037c83;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7416d56e5592997ec4f90f19fe19df35343a06cabc86634f2368d420a7d2211aae5dd593a7c9a1573052a411191836ae46d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37ab3dfa384ec3dc99f9340282deffbe55d5b485b092e8a22770b830321cb94dfeb1debef740f4c4d5080aa9f089b39982fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ccc41ac1126ec81271c179d9ffe38ab2a44bc858038f0ac67931c226e9d02e1f176bb25822ab41e0ff30340a669662ac762;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h573f1c76d2e2a7d68bb65f09415a1acaaf1b83af5e5526066dab2eaa6d6a352353175cac4641bd686254d7b00c26d4ecdaa8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h299e50dfe0b7aef75971dfb3a3eadbda711b26e25671e44458dc14942258cef5356900bd069610e51478cfbf4e208100834a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7abc5e0624e277af84dd443570f3192d38ecce769ccba93afc9e4f15c8286f8e0078bcc928fdfbcc634be51fc0152cdd4b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd38b70e5d179c1b773851290813c0c4b03102677409367192214e2a4a63bcc00af9fefd2f61936d67cc8ad04392c87749fdc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h358421e9f1321c79719852e09b4dc615564a25301f8161455f7acb803eb97535a9a4654872bcb619284eb729a6fbdd19df8e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50dcdf1bed0468b97a2a7466fe4d4ce90060ef67573d20dcdde2521ac5e66412865cc482558a89f95af852b1f07e1023fb70;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f4027c5f04270d221ce27890759ab4ddd86dcbf986a070e82a5918b0ce2026b70416d15b3c3cdd34f28df507ea946ad26d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h725a69a68ab56cdfee4faf00e5f4b808e1732cef91809a65f4080f01b309328a4b1ac047e924e51d02db8451423da2578242;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63066dfae5340293c06340e7242e560af84b94df3c661a9e63bfb51ba9832007c9c027d0edf63bff53c94887a55e23443eb5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc31e72e4259eeb60706a2827e603284ff309e70dfd893a0fbca803b6541f134c744d4dca04041de71182bb74a4f07b22be1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h403866315fa9e9758686befea01a96f6b44d54165d4ff15808bc34e8933205aedb7b5fbb20a8f1e737b82cc71d754c2f9eed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1b0c2bbea4bdd39f608f2cba57e2bd84628fb355aadb0ef6d641b2982adf53d4726ddeae3fd9778d408b4f1255cef9ebc46;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4afa0e53b1814da85592efffb3d2fb40efada88af1c1313a2d573936b77c40b0f03df5bedf0160b5f0b75a2c15f9bd5a44a7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ddf8eb313223bbfee0439a260d2b97b335b2b56ed675526636e0b0e9c0a1e5eeb0559ed3b08d375bec5b4738de4ace55bbc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41eb66191613c9a0b09203916a8b2e4cb112f21682916f5648228ae2dc11933a1e4988fb0f2ce3b8afe86909bd32552de551;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53fed4cbea88796003ddcf9966a85e1d31b570f1f9dfa67203f7f9e7e000c00f13f0c6521b4862a1eff795c8d0b2c553c1b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc771132f93cb71bc8d596586a9f95625c0e049b62c9c67ef81ec8427e42396d47288dceccbbf9a0113d0ffd83fd75498460b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfaf84039dbc90b85640ecd2f15650f060099cdee048b4a444a9b12963af307f1db21bd90fa9d7bf5fa9b534c60e0f36f8f1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he32fbebc3821bcb468b6603e037baaa16158a95f9dbdb96e246c590db5219a882cafeb83bd0cc64368039db5d079794a5aab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b291cd2d463fc7ac95dd8a84ba923de656ff00cae74940ec1b71038fedfcbde6981f06d67760e1a3f89d86f9e0e4ed38106;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b8662d16547f16a3df309f0bfc6165ff5248fd6f9109cd3bdb7b56d276fdf2b393b602b9859326e5018e808633c8d5f1860;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h646079fe4b1086788976759166358f5f8c02b33e85121f45b8518e4b461eaf182aca3cc63610234fcbf6ab436090bab1eeed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9b5ccf228428b7d8631b318acfe5da7786ededd527830d35df4d3f7e2eeb78d294dd6804624a06b9e379d4927df73cd4285;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3bb91f05e670047109cf5fa88dbedc5f10e2b139737bf083f676da88483699a2d6869c5ad08aaef97ba8abacbc403b71c8ed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc9f8ee6bf807b203f6860ec763aa6c547de67139cfd8c1613e40fb603df7acac4ef3734c8779797d03fbac10842d45bf39c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83b0fa3e9181c20073c4ca517bacd4ff66418f1afcf893b57b415eec0eadd7114435a23ea9978a2e1c85fcf04b5b012f7fb9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h206827fd1d42e17c1429472e1d097689592b5d9308e10a6bf80d5282e3144e8ff8df5135f95af457ce1ff1e2764dcb4c7700;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70d932458f38e3d7db09e00b069a619024bb9eca5c787f7f6f3761a0f4a4ae22527a39be56a1a3f6399f638fdd7e47198aad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heaea6b4ab92e904c86438d9a8731c1457b67a92ff6516a525a2375b696c45d10605a9a8e99a2f4d9a86ea2f27604affc5312;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1042ed2419e4ac99b85a415c0c0f736144f16ba21d7f1da5ab0563c402c445bf07dc9479b38fc481d036100542bb1d562769;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha549b9e81b63e8d44623869f69b908303e78b943812df274c1a2b46ee8a85be38ff68bd194361d7cc0b983c865c5a6d3f98f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90897fd72ee4fe31beba75bfce642322ff4432ac0b41e710d4d20d1b19996e7cb7a650fbe5cff24ca8fbb9c3dde051ec99ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d2a58df39160cc970ce3e6d280a96e4493791499a4545e97b5dd846b2f87cc86fd70353e2525c5ea1715acc22d7440194ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63dd8016457eadb06014f2068f7f8e960ed2b2b0b8af47249d1e6da423986dc4b9ddfb95c699e2a415649bddfa695a74b5bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94bf03cbf25b3f58b87a08223794e7840941c5392ec6085927501dc0a24883fceecf572336d4793e8e6c868cbcf211262248;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38ab0d288d280ff9fc5a3f693e131c052f07bf37031a8d9d4b8960ccc50982d2cbd004313dc66cc3acbd660625f3ce58e6e6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61774122625bad647713ce075ede2a8e400f2cd77fb972c8c0a5b63017cde32411db21e76ea3cf482ad4c30c78696677d58a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha32495f5527ea5de41023e36a3711b7c9c4a7be813c9c3eb60a8299ce15d993f1f93767c99ce3da84d00b3c56dda2b3f04;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hafbb56e92a0b4d36d7fd72970a6de674f4fe3887b7fad37d96068dd10e33c6ac15d26fa73be1838e8e4faf89e9325b9775f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7705c6262ce5e150cba8a855922338ba32dab606fbc767b835e7b348ddfc2a09af5097f49a69de89a48e85632319018b81e0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ef9d31ce64fd5eb11b3011a73475d213a81c5d96d6cf4bf7e10f6e4edbc12d54c23922976db4efee8770f7a41c7a6f947d5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c070de2ca9a7a2d93c9841661d7dd2dcb8c8ed716833f66286da034e650cf9f8a22b9654356a923728f298d049efd2848fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8712abf866d7a35ca478103c2cbc00858e5808492388050964d407d255cbcdf232b57eda1f811b99bd5a1836214cb4f677ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69f161d060563f5e03c0810589a6c4e049312235397064d087ba2c5478f3a0f0cfcdcd95695cffcbe6b59689602a8d2a450c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcaffbd42cc619f981937e2fcf6d1dcc3a2c1582803a0a94469052e943f73d4c3cc4621183e2846d2f274c9b010696997b90a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf57428d1375c681dd0a1fcddb39268abd0cb4ebc1376ad0ca2f5bceb5761076527fd7c2b2c6cad48e921c17a977e187eabc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0b0e7993f5a745949ebecfc228f314f5cd31da4c2f5ad1de49eef728982cf9a32685e015db3aa6ab535a995011b983bc67f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8940db7a4dd8ccb3cb0d16879e5b5358a5403ae4dbbe387d6c79edf4d1a5fad4d79df475d6943644278d0ec3773bb1dc68b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb13be1958499d54c64a5bf3dc40fc139c7ee8e2ed289937e4862e8c2667ee1f53e560f05f01d3be8c3a316a90b3bbdc54e08;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a7a31a9188a06665af0c4cbfba265af4d4fe19c661ca0b18cb09ea86e09099b540554d30d25e1940e18eb3bcc754bdf70f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3593a043a5cf3c0a8d93076232deab30688b822e284c6ad3e2d23d534a798c660ccb2c7f4d197f9fd0c2db4a76e2ef049fe8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb120b97ad374cd5d058991b47209bcf4e5b7c3d285836a84c954a0ea5cc8bb0e6906b935300e2859266ba62e271c6725e8ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ae545f5006935620104325e484642133846a6cac4265543efe162a045d973f62f08aa4291098f57a2aca42923f4c4408543;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ca42eb3a8b468c60341f3315d85503037e8da1974e025f04da2ce5bbee653c99614f976e51ef587a5853ca2ed79874b419;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18b9db6baa9e8bcf00d17a8ed4adabe87a7cc72a817c9ad58ef0fae54e1fba0647a5bc10c9823b18e5e5179456da72ddccb5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1db73114a846c9edcf3d0174c7759ec2e4132912eeb5038a4eaffaa1b65c9ed30ed6ff4c5defe7f4c62dc8a3de4d395ed7aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e86f5783f1bb1cf5c782806a447cbe9629af86affdc1259c358617037eb7fa596286293b822759cd414361ecafd5d5404b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c4073963d6856a33b9ac2809e1ae46a1df81ec0e9af9260e13926f48c43401ad35bbf8290723fbe86833ebeb3ea0c43bc84;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h307a83f9df629494a9f60965b21e3be3de4c6a7f54c40a2e35104d7a0ba622b05603ff7bf9de54be6ff8819afe8645f74ada;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb152b49713028c4bcf3b43ba1b553009d131d8b427b912a25c871c6755b0c359f91ce00cc87c3ad152f74d9ee0c1d8dac65a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5f7409d0138bccb9eb70a2a2d2dfa62f2797e36e603ca7b3242d64980fa1c0396ed9589dce67ac7151f56f711efbc80cb76;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8391527107ea9f519cec55775b72f2edb460a214f4fa5f1d779d1ef3e9fa1f237bfad8a21334d2d789b51b9e8a4ad07059d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1f763e28a9d6fbd84d0556528257c9822356481233fb0bac85b06335cb2e16cc637f88d1a9370f002b0b1b469c3a8f9178e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8af1c3ad56cce0a157018a0e32f81c83d1fc90c1cf07bed597b8990d9a7eaec74121d890ede6d2de39ffa16b09646cbe6bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h511725e57671362d11a89c550dccadc2e67737ef243338ce36baf377d2287da6473fd4f06de21bd10a04ee79cbf1e0f3d0e4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65c730fa1610e751c894d94b9e63d6f3aec51083a80e784eb5ec004af240b70fe3943ebccc25922993664b13d0f5d9754172;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95dbb471c851ee6e7dcbc5dfa021095c23e5193efab444a78741c1efa889563b57b8eb3cb0351dc2286ae77021962a91dcef;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9fc41a43f9427a15b9e4588d8789af4ee5354533c1d8719acb4a0aa171ea6bb58a6f9a883cf9e0be97a06f25ce783088841;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5df911832407b8aaea1c8dd9557f13daa2d6c7ffeb6b2a1fb6cef0e509261b796265b1bf768e41c7ced4093e36a6c765a3ae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1083f31c810959f43935b1e0e26c3068a057557d69dbf4038ecaa7291847976c4fd0ce5dc45bb7a2f0e71429e31171a2aa51;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb4a8a3ee7f24a5c636d2b6c2e2a600aa772e3ca789140a99583be6d4cdbc5383baa52b60a5f90268b81d20a00d24d924187;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f0cc25014bf32dfa871e3b4c16f88e2fecb4522b1fc9ea3f766fd2cd8d6b731eed29b9db30d14c763fde7d700abdb0e9be6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8c057ba71ca0e8e4aeb66939dc9a8be67167514c408264f54db460443a405bb01c21ee92260b608f3de6872dc90adac5c3c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d0736334b1b6e483e9d3b1a048110b63f36463eaad7c719f47077cfda994307004e705e0873f71eafd71133f3d80723ca53;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4330cafabaa3936d42c55720d21e01d32ef60b19fb6d0b3b16de1275e719fe9f70ae4521a1acfe3a847f728e7a49cec63ca5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84af8bc84abfd1d9a27b3efd6bd7e7f08efdf727729aa2b204259a5067bd464a5625d10ba2827319972b7971c5a5ef29cfa2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef667ee408cba8965c745459dd89f8505c99d479a611cae1ef90fd7e4590fd4ad0647d3da1f48847f5894b77026cdd16f33e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4140845d50b8dd00a412f540ad8a8a179235e56ec07ab6a602e816f9220e30ed706ce0ccfcf6f73e4e2aa1ecdd2a0a2b9c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51183b25283c3999822c906b315e27d70f288d881c48fb6f928d9663021caa257e275753ccf5c7b2929784e4831860d2c941;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fdfe0dea2a594353e3ded8341c6151c819769452a6fd5341fa88f42e66d32ec437f438ac07f48bed46d6003fc211baf2ea2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3332f59fc30d179cf69b0fba0ec13eb8fa88b2a4708e9dfa9b383a8194219b8588591e8f650b5e7109bfb7ae8cf3c28577b3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ecc8992579d4d196d7c955ad48cf46c5e10d8b1cd07d00fd150730f08f8cd3fbaec50964c8a251263654ec583a6443256c3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c5e25cb27feaa9923d41eb8c47bf1adc5683b78120a8d570cf80986f9e86eb1d788e42c012e0eb13ceed5464514fa335ef9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10add20827bc9fc22c16db33b7447f843cfed80def867ff94f3083b8c8dee50186a7978f3148065c69ec2b33a477607fe3e0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9a56b75250e892af12adde655be9f9b7738af9114702eb56006d2f4ed81b17f77588f72174c2efd315fcb54acabaf4e4a75b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h279021d5ba529260bf55954b499b58b6565ee036332d92b0ba7e67607c157c8e8ba740d87b018d1020d02110d38e42c6bf3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h759c43e25725408efa4847efbbd6fb7b103cc5f1b3bc52373f4dfe8fd9417fd5ba6164dea360c54531ea20e12a80aa635674;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd29b7131d8729c025ddaecc845f4377bd57c0364fe1982f7782c613e6976fe8d2d83a123c2dfc7f32a86532cf9a29757045c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bd121bec49cce29b470625c84e440c92ab9acf15a62ac1fc6fca3e510ea30de1344342d8e1c46c0174bf89f1fe8799baf90;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3a7521f2582f2662d54198cdf92d5620e431c72e18801f1b73a53e89e7ce544e933641e87af19297ebeaf2889af14805cb4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24cbc1fe230871f8eb3e5f7569cb97f4f4c7eb66215d43612789885a7936228ea1fc805cd1e1e7f838f074263f766a588966;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd51a718085031b4b2adcbd6b1a6fd675d1a25e59106277394be481e6a39a91ba374f1176302455765d399c6b7ffde9c16597;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf28d2cdf732c69dc8af70a7f519059931c159fab3b7ee8758be9ec504438fc326c2e58368afa4b0efa0153ecb5dd08fcbd39;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8b41033d0f13e77dbf6ce260048aff4fe019373fea92a605f7dcdbf61fbc0f913055b44dbb72592297450bf0ec6e72a5771;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e7225f518a2d6d28f76226b05ed07d6f48c1a7e378689c1a0e350aa116a1198ee0aec7038152025294b920e6b084c15018e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd79eb6d6904e6862311c28bc8aae0faa0f0ce3d96c5fb16620281233a1ccc2fefe912ef0cc0eef344b3a9f3955602f3bf1bc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6da7f168c12fa84b0e2bb4490f0efc30cf3e828257a1f517cae2c07baaee8b76b01bad7dbd2b69e75639c4dfb0b26441d996;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb25e83bdc669180977231d31650a09a2aeb32e5960ff36f89a8c6c4e58ff729e545ceecdf72d7bcf1b8d7dd2696c0c2398f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb70fb7d1097dfacd43e22629252a732c5cfaaf1af4a0e578a5395213fc7c58b1bc6e6f60e885b5f195c14b58877c19efb338;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32566d2890077d71db4c504081a811f19a3b57bfc1a1dd6d111ad4182720fd830cbb6bad34df7e819060f1e710440c523845;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf2bd02abfed9ae7819f6e0a4c3d2e3c80c92bef3094b88810996fca8ea04cd896ced0a192dd0e1ff22f8ef76af5044997a6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h410a930608f5454a925f61eb6ecbaeffbc001a2c9c6dcda15f0759e193a19ba8f75db00cbb5f37e116e42965a7995cf7a175;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf935f1e2ebc07e58bedda41c3e409be1e7670f31fc6a3c67c9e57c0c7905439b445ab88684ba13305117693c9ff243235d0d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h323d67b75ff1e803ce7ae938caeed48e750e90a9f4ea747348cf2a4fe951c98e431e2d6fcd42ad47823bd7de345d4d51ae9e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h836c7fa01f9ee69074871afe3fecf9572b8d8c445934ac1955b10e0099b102e686e0c14fcd07e44913f06cce28daddf5f31f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcbe7da2e5c17cf8de903b025933226148645d85399cdc381e1d48c873ef40509ac23e7328c17bb48142be00e2b07f5ccd9df;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75d6d28842727a70d7d16bfde4d2d6b0b9bb0fec0a1071f3471cf427cf4ad67b3bd506f54ac7a13c7f5b9327927a077363d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha246693432db483c181333386427348630c39e0d6b49b7d2a3552b5a804e36d096a080e0b1bb5d4e57e561120283e70d36f1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a57a38677c34fc243519125ec1ab847d2aca4a79dc145f8154c10a1b55273c573c9ac4eee477d13a08c0eef609bc9e7de62;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2bb2faabfdd861028cfc950c876eadab386eddfa283e7d923a3bdd14d87e0df27d0b81ebd25b105da61aa0e44f91482c2f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc9803ce74d98064ce021527664cdb8b5ff977fe9e3566f6f09c6b5278a46adc4d4ef1be908831496db74775654844b3964;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a24b4bc3843ea96988cf49a30f918c5b71501d287ce6db3954ed71f65ccfb05acc2129926fa1b5f6024c5572d1704c230ab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h465c14c6ed1dba30c940e51f26a7bd1f8ee76b5bc6bc85cd12835c3bc634975ef841718e938c70c31fa746957e66fa0e2afb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf162228afc755d4d274d2144afcb88f9610574fa0242110c8957fbe3a4fc0d0ba8bbb9e0529546b1a81449db35568aa64d3b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ec1689e048a670003563908f84378680b340c8be5e9447d915d658cf9254843ebd76254fc3acccaa9100158adcde0f2664;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf77edafc6bb2ff2e493e6b356c6baabd4977603f613ce9a851f2b47c730753f0e0fcac8da909a96ddf3689a027f8fb5d3b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10c7dc0e5f54e6e745d5e978a3d2384f17d2d514d4f92a4d428cc2ace31901b9a6de333558c6b2d25cd6241dcc77e30f126e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha86f84a96f451777b81daed69aee373094acddd4fb76eb6a6a032def7dc3f222afd21f18e3fecb0adced9867e796b1692d01;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2591d2eefc768529030b78c81e09d7afca55d9806ad7f8ca23770ac31a1df04fd127dd38c3584a81d7b13697909de0bde1a6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha33c783eb658142b8ba17323bec706d7f12f5d368917d98278c2d3a8b7225d0d808f8a12ee3a97a6276f68228e97bbb8ecca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he151478b4c7eb41dcbda0e30ea11604f546c34a730bcc8936e10afe3e6d575becd8993276c34d44891fbf090c93fcb837957;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55f9936ded85f833abf1fb11e758994b6f3cc10b4d1d29a53efd28293e3f1878620b5a712744fe049b4e01eabd80e5296932;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h323f25c8e89c68d4d0ebbcca59d973be83cf3c0e3ed52126377aecb94612aaab9df049c29fc2b32ee959fb04deca3b96d3d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdb2e557e514e7ce52fb2f8517887397ffca49583535a2978f638dcd483042b8bdbf69a15bef9f61083c4dc42313d29ca260;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0e96bb50cd39916b413312e6b013de659c78901cc9a9021f502ee1d409201e2fd3be4d71b77e3fd18c6b8f163e169f09ff8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h525cca409ba75d6b4d7ad3159fa7ddf2bf4c1f85070489da529376de2962af9888d16f9f5977952572ffeb576689fbfd2be7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd383941a77969d9a5a304972134c2231797332f32fa1ffc0beb4296bf85d86ab3f6ce559f1e9c75dc14eea7003d1b94bec6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1898018a72e0f99bb9dd33b0b011a32008a85fa5ec311e7f58562b9250e80a74aecad0163aaef50e11d0612112371c2ebf1a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ee44b76804fcd0fa2838f0895dece8a3d207881d421cb9f0cbf91448173c3b50c296bd28b458c28613ded8e0fa41ef7aed5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb8a5c86875163050c512396eba628e3fdd638f0dcf4277a12cba9faa2b11c6da378e3c16bf34536fe37c50c8884f8a49381;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd11815c1c39bfe84f1c3d0f9ee05bcca3c134e29195f65f877e40cfc45a7bfff53e50ef27fd15e59c1b19cc6157426e69a35;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27e5c80cdc4789957c59fb920a22e0c811a1171310f1b2d6bc42a6827dcc4f98e75d190660e99f5c089bf936cc8d23e496bd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ad5637d35a53f5df61bd2d5547b72388bcf44e35adc0817dda54c435c8b706e8f5b09e2390f4f5ad4f385bbd7920ad036a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13d3394bf545da0766dee9cc0719e7a162f9da426c7225286b938925438aec1dec3097d8de84bd439a97db2e1db235ec7d76;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda9204e556c92890fd9759f1503518aa388225fb9d95fabeee5a3c3b72d685f51abc1e98603219e38b9efd6d65e9571ef39a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7cb49da991cd303468354ec885c697f7497acb28deaed066e1811a5a6aa785415b412011a484e3093fbb3731c4db388736e3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae25932606006723b08f07f14b526a9cabd89295a74ecb3050c09fd016f4b9224b2dc829fe44ed67139c3394008d0ef94e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc90035b7ade390cb9f1ef2fa1074b7e415b0b51c4ec2ac5d8cc81c4ca5f08e1533f2d9dbd0e5c0c5a57ef398ecfbb9cd7168;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebef559818be09130b78b0e9247e7569e7a09ed687afb3c649afaceabd175074b1956dbb90db6dd5bf6fdf06cd6606bbb64e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71fd35caa6b5256de51b26cadd3514021d270ac0483f56b0a21b7e7e98c93180260b4313f6d1f46021826973a87dcdc44208;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebb351c4b7306b79e7fd9a6e1dcbea375f6c3482104f9c52f184ce1e3f60052cb8c4a9c4b8ba8cbfc4ddc02881819f28a6b5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15513c335d42f3f2ba00b60e188bed9f47dab472f172bf0f49d56b11568e6ac1de5bbe000715d7078f4f0812d75fb0f8a651;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97ccb35faf24c6cfee08d41f06131abc500ae3d774f23d7798af481ffa17592dc9a26551b085911dacc31fa23c920784a2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89f3f4e5504e0a4e4dee366e64f55d6ba983fe2c4d6ea5a3187e07a7c8b9e1d6d535f316e2a97d1345ae13186bb1fef360f7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca07c0ccef2932d6f03b657fe974cd4e570fbf27e001fe49c4bd1629af0849e49d43f51c11dc00cd1292b748af2647bc76aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h958f0f7d0eb3bfcdfb28326e7b000fa17d74004e287c13f1eac87334929d4eff286a4f6a0a5c2ca40b508d04b999bab8fa3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cfc9fc76c7990ac346412a4c268ec0bc9e1ac779d2e1209cd1426c69e5c2c86f6597484f558d7fc040fece1806b13cbd7d2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h518b20ab475dad8d689514f0698387285c51d920a76f18cdc412ea0eb4e360e6df388cbf11e59a81f861aeee99cc113a5c9e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a7d1f89ed71bdf205fbeb2df3c1eb90c5c8a13356b31194dbc39b0c86cc3a1483a8927ad5fa3096c9c3e4d6e10f4df4d3e1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h682e15d7dc4e3faeaa4b5e64c17ee9bc26b842d45dc2515747c6c98f3fd1acec6850a4f5264e008536ca05884ed4a8bc1105;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85b3a46482d20a31a08193e30c2a2441684de8c84d4cadce17f7ca7940542b6e32683377c5e1754b949e1e4ea4a459b281c6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2588d0cccdf59f34f6faa440c97b9790a6db5bb3ad4399c4db2c2742abef49edebad3bbd021e8ca7732647f4adc7aeff90dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb688a14508773a6d700b7e71901b3f13eb1fcd31730ecfd7be153d470fa3b42609a4439c41588d0068c33a6b3dd2fa00afc4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heafa3ac127abf64e50c07e413144f08bffebda39c274dd93f8cc6a8b8b223c8f1a0581e335f8ce63f839324ef2c7d6e392eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcac99a0525a04439a876293faf22a7afa729b6a8c0aafd83394f5ef6334796851c85fb8012ce9f7cf3adbae8685826b90408;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2491477c023367e5e37e2fc6dcbe47f6608651f18bf74f34c5faec77d8d47d0f0447573d970caa6bcd32fd4e7903ffc0d8c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9faa81e787cecc4e449298c95c96d5e9ce82589d4bf9f5cb74df45026e3764586ad19278c47deb74d7ea4b9106035911e5b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d74fa4a57a75c4563c70db4fda257659b7415d21cd04c2888d0db3eea01d51d0f3bc7ca9d2bcd11f08d870c5d913deaab8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he02e64ba98e9a747e8db44ac631c91730e0f0ce0ab73e0b33ff32d674d54288b92f3e0b56aebceb65799127ccdf367cf3b75;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95d4fe93dab80dc3ee9c9a40608cc30c24ee19e074b9a37b71bf84249261dabdca58c3537c3e12f104dad05f23df0341df9f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42df44b7d6755bafa5df4249b118206be1c7f1b51ae3ff3687c093627cc80c1df565bb5e866682685aaff4aa4b1519625042;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a6fd3ee003057294aa84297964ff263bc6ad5c8476795d6d78ec49f149a712d3c099c4aa5c2de35f87003614f0d0d48fbb6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2dc371558fd0d78f00bb98848c46cf0c3db6c8c1f3f19aa90d24bd08e9e9c7b90c7b15f460bf13fff8a85ea1fbd461a7a48;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf752a7a72771bf4deaed07b551578fb65e3b59ab03228e4b5163a998b4542ffc9426b2f1f576e399bf4bbdbc1aca66de6cb0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf9b91dfd825d7660b942f4167e16575668444320244c02c477070e797ed5fdc2873c598325ab00afa09299dd17b7bc3f9b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc97639e85457fb04cea0886f4e2a85a60b376970fef2bcdff7de9ac2a368f39f52e383ccc911441633c39fd227dc2a590c37;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6588ec6c9da0b229ded4214de9d380064a941b525a135ba8e05dd3e133663604ac209171dbc80f89826c5e24a59c239e4d5f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a1bac44b6e5a39023cfaa9a81bfc9881dd882ee762725bd076b8b4132d4ded138c4e866819325a509ef31692ad48e595c29;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdeccb568013015c7d2f35b17fd6cfdd10ce92201940febf81b9314474d163fe0201e0c8126827e7dd56f1800481d40bc7aeb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62c3475ed8c13fb41fee8ab10ad925dac67c1654ec3e71073b95ed4094d4a30cafc2e4f750439c350d99511cf63ba0d5c6cf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h939c3b96cb08fc8a3f6bc7282290f8efe5ff5151c06ea88b9b4eb297d91fe61c8bc5fb76c6eefa2f2c925446d3ab47858f8c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha31e901c8cc42b652e581647bca6540b7aa703eb331f1b47f3c7e99fba0b465f1f8cc49d2be746bf62a2338411d220254141;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fd4d3163cf4b70b0b95aded9483b7a0eeb5b6ee14601434b528d371ebf302c386f1ee0b2ed0b9e378946b939f903c6f04eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h570564b258e10300ed3fc85c2dcd6576a10103aa731fa6007d7646085e335b0641bc6d500eca2619f946ab19e9275125725d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7029cf8d0e03bdf878c872ee1e7a03965166cf6a865770ae54f36564f465aa3ba7845f06199c4e305903d82ab4d95155f33;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c9495cce410116db3bec8ccbff15d736cdb42bbadcc31175bbe57e2b36926d2c0d3642f2bc028d912f0457c0871e43a5066;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc88487043f65e17951616992fdd17b8e3df8e179d2aa4a5b693969f58bcc00757756a74f71e117eff7c35f4a8a15f1de6dde;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7aa81588a41df5b59a10c19202f68c0b7f0375b8e538478bd51798c255554a7f5883960347d29ffbf8f668be54c196ff4a0d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc14467db9daa9a1203d5ed88933913d5169844cc27365ffd5b61607f4211c302852ab70c81bdd417f4e6aaf1091eb885a7e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21253d060cad9ebf34627e2e4a1b062c0bdca8ffb82c9a42c3be7bac410fad19b06dc58d74adb1cc0bf39092b7f00994a95a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c1f73a64eaf40997d95bbd502c2d6896e88cd05d1a7b5f2f6dbfd75b814691474b079c75d20a777c2352acbd1afd02719e6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab7515189db432962ce67eb7e0a33bfd81b9953b4f7504d8cbdb33c8f80b04e61f135216ac0d6f3f46392aee0343a8eda62e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8acf2582c90a5290e9141679f35615876a2c4814fd450cc30b0c946a3d148b2b14667407978f3ab3b1018d2ac542fc7e167d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h816bb503bd2c6280fbaf46c07cc65e1a8b69a3ee9b962ca4c5da6c170bf18c05c478f551c3960cc941ad8aae9674422a214b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89199f3e4036196a8f0f1491117b89199b5ce8428b969920bb22ec8a81c9573849c6cc55cae476405a44afc303eb94852081;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hafb182fc77cd9a824c85f9c3502976d2540cba3a41f38e2184f472320e9de1e4e40ba169bb36fc971fdd3ab66b0d52787427;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb80494e1f112b19e7515b9974cda0d0b81ba23fafd30b78a6f0bfd48b03e6768a452d42c2660072eee9055909588fcf03851;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf213893c3c2294adcf406dd33d55a35dd9cdf964aa5cbbe9b07ba73a7d4033c4136d7feb68596638f1f79c778bd8843981d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb3b096bdc453a0e671066f5a9cbe9300667d81b00a35be9bb93904f6f85b3ed82e5af5568dd71843a57b698574a77cdaa95;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58715fefbdc011bc9b76a504cbfe2c668199796843b70eca34c68808b83b32e427fbde635ec8cd49f01acb3122177d03fa2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66f0c6c7e4f405d5396c0d240286c23de7ffa070c7d385a212c4b94cc6ce872e9297429d6b58ef1d165238e203761c456e87;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67b25fd7e4cfc36f81b8ac3d8a29d2c40603ba1d84b12b3cf0d39d274f915309ef01765265163ad24d5e417fd5f658ffd077;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h850926ac70f0ac82effd8bd4a3a50fc71716fc67363a5866dae77368532992260064ef04fb35dd5ba699080dc31cd6a5cbf2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb077af1742027746aba0a827f5dc71f5e141bccedad8dbd5e8ca50b956e0c0209cbc60f0d787d40129119e47ab301d5ccd85;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87597733ce28a75f6aa31ab830a972deacb105e1dc158e75cdb92767978bf60eec6a4fe9950793ed5f6a11a1e0cfb06ed9fb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9cec87bd46ccbf4b33691725fd8713f96c7749252f760f6535f79b8ee249fb05faa50c5fa85013aea2ac0ecf68ea1684eecd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae2e1cfd58ef390d9c8a7944455f9259282960968f900b11cc1e6fa669c98de29842d3db6a619126c7884a39e3a95b90ebee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h503efee975cf4eb13c1787559ea63f2bc6b0378c3e9a431a8463abb40718e805f0334727e4b385ddd2aa7e77e57637d21444;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d31714a3c3b04cd4809d9bc64bc3d1fdbf18f8586342e97548a21333390566563fe7c58d3c049071f5bc26f7cb578c32528;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c659db44c99685d6979d77910becaa0ab4b656e37351fa8cb27ecd6e8a43c12c75a3b178dc0bbf57c75135a74c1678cd1bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6d1f7da220c2fef387e210c13e3e2b1f898c15da35708b3c984940172db71dac820ecf2201221bc8c650c89b8d0cd73a3d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he82a94f09de50d6b082f0d2c5c38f7bfa5213c4c2f0937b08bb9ab25d0d7ca12f194d4307a3367c4c5ebe5809f4c18daf1fe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5e2bf2639f59a394bdec32703b88fb4b8d0163a1baba809e7735539a91ab2c7a543c1c092786e3225bd37cbf6de8758ae41;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a98306caa6888640dc97cd99d9956510238c161a9d92f5562c5a3326657de471cc7277c314172d69374ea74c894d7dfcbc7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h54c557c331b260c9ccb41c46bd2568a4934e9a4c9af04160d411acf79731ba6f27512e68ba7a768cd094148393f173331b36;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb677b0fb9dfa68404a3e96d204134bc0a1910b8b6aab3d083903b74fe5f19f3ebdb3d53f76330d3da091f0c1ee757c5c590;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdffcf96a8e8f84d8f521aa9afa2289ff7940373fdc74535165323e6c9ceaa9144b2fe087c4c67c4589717391e1a7c68751d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c5a12102b1c84040573cc5374ce03e23f5dbc1038ae250ef679a819f1b6fd360cf44e5a116190bb05a17eaad7f2e0c15cb7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ebd884dfea71bf196a2e436c4f35d856cb819ba37075c4d1f1ec9fbe867ec875dec184667fde00483ae90d4eb9b3a492522;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h695fa150c4a3817f847b311557bf978843f6df90def6664be76291acaffb3a1b7f00824a31cd417bc7dfd9501c34af12f6ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe2ce555f2c4f45c8b0b434ea776814edee4ab0b94f9160c15d5a78c536eee3ddd8de52ffa002909b24118ae533bdf4ff22c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd47c33d804e50690e471be26ce37c6adfe00d750d57df26710d7f413e778797539a117541be0765af8837fbc03d1ac56e14;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h653506a8e00e8cf8af71b6f3ea0a355e65e93fc74034e74699929839b7b4318d069beb7edbd56c293467973efb60d832a17a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h147e4472fd499e37930c85bc03a153a4cb26c04396685f5b103838deaa815b9bf1cbb92804a38f35428590f903fdbc0baf07;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc82555832430e33efa057a3738e07721bbb386e36733e812e923b945cbd6e2ab82357f9f7987939b4f955ed0d22332579b57;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ea8dd047bc305ef68e53c2f1e9a89f37658b29d8faf9acd2c9b1c6641632352003d2272a49ac9ba470857e65302c1bff027;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4117ae79f89d378952b737c43a2a5740550828ad940b4b51697465013b7015095a393f73d06c98561412d557f05cd4b0d949;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15632ccb329a44696c232f691bf63a48c456fd19b851434c8a2ffed55ad740d9374689e380a9278b36fe988729cf81526e78;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h194276ae7aa5bbf345825c9edabe9d3aacfdc1730dfddb09d20ede9f8e58486d246d9336a4e3fa5781edbd3e3b3aec0c5277;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heea2ec25ed6537e7f8aee62c93e889a22d7343a9a50b0e1360bbfe4c7d4569d6f92dc9414958f81ddc4bbac32413c900fc1f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e924e6f9001dfd0fc0304149652ce4f5828ec66af6d98a7b740337ba1870cd767f37bcad65d55cf5fda3fc9c4258f22fbb1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9fabd0e15e3fe56b17f80e241be4b7a00eb2fdac493ff3ef3b2749107d968e2b60c88dd9e98eab625d9ca83b7f6863f9a66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3dc084715125ca671204074245cbea187249723b48e735704abe42923fb175a5c4d74d455368e3cb983dcafb8381a60fc09f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bfa561e5c5da1b7671cb7caa0a67352e659ca2894a1f4d79eca303faff8e36d0b23bdd85baa98fa4b1da17e2e42fe568ef2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c112df3cc265e9893897f7a81898ebfc92dc5bce79071d347a35c86f78b2f271a009db2f8ddaefeb32452fbedabea3b726;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8face5b861738680610ebc63abbe8ddeefa9f54fc04a39a0b52bff1a47c0ca44cfbe7b2fe63c702e53f8d99cf0fa26aa904;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5336325b1c1487952ada675967d81075536ab1d00575c89866df8ae58549c5d511ddee030efc007a46fb184b1ea9b8b3c289;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ddfa3843b4b6b87904c02056edeaf2af395208ecb3f846270c25be6a83fe54af413f7157adf6f83bdef45a4d934e68458de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a0e03f82e35a23cf94d72eb4030d6173b1ab4901e326ca082b74846f3614d7b99135a64edf1c4d8e2e5de9304be020c6721;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h42f82b56b625b50a6c9f09440da38c981fe2115ca07e99446b50713cd7971b040999dc84d1fe8aed71c756ef01f76578585a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcca38befc6c4117c4359730a4efbb2c8339b82b8fa4c09cd982124807f7b69538db410eaae084466dcd0f36443e877c7a3fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2a91bc0570420579dca9c6f1d5231e5019b281b375116abed17415374bf32274696ca2222f53403cd62f7b25b2c666f69d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9eee26264ce434c4b071a0e926a361cd517e7e525f4009f8b6f1ccfb7dd30a08b6152e93e94ccbb3f500ac26e43f7f9bf754;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ef976dcc6d9d50af774a4e6d2bb5073eac31b5245b83ba86c5fdbc49c65b4146fe738fc32c1c10d8c91bdc21740681ef99e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h318a785735b317addc1a37291045ed3a1a1ff5873a666d7880b581c3406303b87884857188b9baa71d70861269366b625340;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7cd74b792679bcff68b804cb145de789910a521edacf8eb774d9a4f3f0d0ece13ba8b25336cb29275e96828785d6bfb036ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d8f8703b473be2f2c87baa70f2b45c958c56a1f3df16ae76f4248faf7e19d08a9f0994d7f8314ad3de5b8d8ceaa6a855b79;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h665a75fde78a0539a091fedf404ada39b6988eae69e422cd447649e0cd71f3b00d8f36cf5812ab303edbaae64af335dbbd96;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbda659313fd31ac141f064df1f7a1a2d60f489a504cdbfde715ccc25168ea8f217a8ebb14f39d50570ea32fbb1a01c0743bd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc93bf091ea8615cf1c8152518315eb70754f85694b4b3325c80b07f4c1d2d4ad0157d8342970be040a075150dab310828d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd475297d06019fbac308722428d1299d8bb47c2c5cfb8c0eca9a3273b5586cc1ca8f46f46b8d109e7f0eda85926a9e113f8e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heeece1b5f4ef75e801fcfa01fba4dc558cff8242896516b7f96d3de3902cc6310fdc50f2e71810d2e16a7be8ed27f53be3c2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0d8d36f787cbb6259b4976e239ff67efd1566d5eede067cef07b13dc3c62cd41d1e9beed5826f68485ba32d90ee26f51cb5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5bb89ca9cca181b7b5ad499cd050ef39d6a87321f479deae419114923cb26e6b064be0c4879c3579e89be02428be5fb821db;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8af9f18681538bd19c55dda1b07223a1f879f0f9aa79783645d30089045bf810507b9d9e617467bfe6e71e5253a7df3bf63e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h817a5ffa120bf04c0475e96b400ce89c31ad1123b4e435c74cb6f6b6d5f3ec530d595f8e55a79364991ab5156dc4754d8b32;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8564a4f85d99290a49da98fe8a7af596b9189f5e9d8356a305505a5ba270558964b2512908d74be6d00102c22fab1dba5e0d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4aa7bfddc70cdfe1e927f118be6e36ef26df1bea9a60f876d15959205196773294aada2818f67b5352a65d10f6dbfb71a694;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94de4a89f61244e4617d096d8b98307c8bd07fccd8a38674c3c3b14476b144b886e2bd9dfff0b2dacc292190196f0167db65;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55444aed2d074902d13a9a5ab7facdfb2ac339bf6f14875f89a7da4b04ecc0d6065686eb141005d4aac68b62c9ce07ee33fc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5015241aa2061567d7d6f2bf8904ee3cb048f28f966e196cabc8cddfcd54a963aeb0c067409d802391904b8144026cce687;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56539169aa00577e52123d640a4a35b460d849765e468c791e68a48bd47ef3cf54b98b207635ed3150f7ba5699fa9e6d8f7e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc67d495b89077fe9115d189f2e4f4641a0b60f073827edb18d68df80f34a946a24507369285e9cc09ac89eaf0f05492d79f9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf923c1968a6d1133debe9d24df40c8a8b6e1f4729072585d5b92fbbb8a96a8f78d41f42e01bb6634389b78b3ec3a9f8b2173;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h220cca25fa8d7c2849b34f508ae2adcdb7148cf1703e3167c1e081b0284df02e9197f33ba57a16050d730607cf3f259ee89a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4c2fe5ad3318b3be060db8aa8413ea22536050eda022ade2208042e7fb73b2f5877e28a57b5e3687b8dbb5f5b2928f836a8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2781ddab7ac924134cf291616c93cb1361140b8447e856cec33f405b8dd28658fca427943b727e91bfdbd47daac78bfe22da;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he80f18fc4594fe8db8c71f6706b235190d7ddc9901d8b7fb86ca0db9931012bc7b7ea684283051c08289766498efc4e4fbd2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he16e0f28ec381cc6bdee0912977dc2ed3186b5ec65ae76a5f3dcad4375771009dc4d424a62ba751b222bee7aad4f5b4375e8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h367a45aa5ff07fc3dd2af4de623f8b9da5411495f4cfa0b6ad5cd7d7d347e5afb91e3ae7bf034d5641b86ad7cab516415d02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58d86ff2b99c021e47c147ffa8606ce4d89111c233ed031f12b142a0e2250a0c203ac8dab6e64b07aa74af3e3702dc5ad5bd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb8d2f791d946b78f931eaf74aecd72e77a1f3c6e63db3198864884c5e7f3017261296a3088428f1c27ca6c9f2c28e8633aa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba16bd53a32bc7eba7736b7b44c6f86b7ab88ea8c2689e514612df0e74cfe35d951bbdf9b0ed60f1a77899b65a6f90951399;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b207bb4963c04b34667175363afbb35080e8cd3050a8162b7cb7e8da16a437f6b2a464bd9966eb10a338a28aac4e1743343;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc38133c3b84599b662a554235ee5a2fd7d098143423f51e0546106b4033979deae7396333118c830040df3a750ce0c07d3ef;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h583df9a27e9bfef2e550b778d383151680fd323b88b5c8e59e7d36aaa695b68835220d2da6de38a02238b15f8294062f4263;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec54f7f95b05e174860d331aca086fa2486f4d65f6f4d3f0a2d798f5fc54a14d5d66c86d68c73907607898f58f66c13db6ab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c7c068b8b24b0ab8f1dee9df11035c1fa24d60ffbcbc19a476b254b2c537eef9b7c3089bc02e88e7d9ab21747753809400e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e57c199c19bfac37aa6c95fd461716fdc45eeee8ce478c00c0653f194a8e6b0adf4b3aba9b5e9970a1e75ad640820812e27;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd21136838fd5f241f110155e54de30c560f3b4cddb7afaba4cbfacae06b83e794f85a3e92055494546f33caf34b4bd986176;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdff444ff565a83364908f1f6a8b00d2d3684600bec0c76c1e8e3d65d0f3298df9f577ad795caf7a60140648db23bb842977;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf7a4dbc7a6c499278c73c1a8d90162573bd23ba2915fd841e32c8f89d8566648f9bf985e73b673597e54fe2a4e2bd60acd1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha09bb3a170569611d7c03ac24e6eeb6e3734640aaccebf53b4ac6066e08789775520a051498981372f62f378551bb189e0c2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7877eed5b976453c038aa7edc73a00e2817a1ec5087052940efd74bdd769b67b2a45bdff8968012576984924203419bae59d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b5b7ee5c79a0f8cb23d68679c2330d76b296e98a7d63bdfec56d657b94848cdb76e79a95996c7cfe591dec27d30792f6a14;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22eefe35a511ff0385d6fdb1db1e65bbdf6eafa4754793cb1d0b0ed3f74c21eef11cea1e01bb82975d293d43ab62dbc16e8a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3e469eda4193d7c43189979438fa431901359191a85afa2160aef21e67ac7352dd5a70844d8d29e6f1b9f510a7fee4f8a4c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bba45917127fa326afc936b49071535ff3cfc350259be494524493674257de028b9e08a27c3abfefe916d308e59ce427844;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h877ac367b1e69d4bd662a4d219df6dd53b2e70140baa27b758eb593a2a3e0a6a381eceb2087385ca382c290b45d0ac69f0d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbd4eec5375746cd13509f52590f617301d19f088a81ac6509eb4fcddae6b5cad833df650c494db48819b2e6cd0de9cabeb3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h667952372684ec7907925e2be3918b354e583a55fb7ae908a7179d5218a4c8b8ebafb510b2c9419290e286681d4c14c01406;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had291153120b600b8d7beb8c4ef9bdce31abefd50e0177fc730fed88de876ffab9316bb0edc4a0e4cdc65eec7fab6713ecbd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd31bc7a766d3083dacd778395a754b084cff36dfa867062c5f8ed682dc39dfca5649ba814ad4ead6eb3960bc444f955d14dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55c8ec104b79852ac1838dbb205ee9ab465190f6c9b3aaf69f0475ab6d5d93655caef9527920535c22f24b7897d11f8e1710;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h387047dd5494ac815b005e632a2483d1347dba1c4c92c8f1fd2b62c95fbaf6bb1d34856b6250c4efc2fcde1e0f2918343c0f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h751f4230f861d7663422d12cbbdccc8884c0369c847e1b6dc17242161cc84435ece89914a8ed3a690a4275eceaffb8101c94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf841b9d73bdcf126230f0eb5079749b635d6d532fb535172d9e603c95f6810a56badc68283cb0c33c5cb8afcc02ce91c19ad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4238678aee4631ac33b25fc713c6df3ccc7efeb0ced1104d50ef076508c0a79d23b1260f194f25b86affa6f4826920303a42;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25d6130275842d939050ac1c2f133a858fe353b55944f10b7f542a1ced4faa943cc71da045cbea0a03bffcc3bab42a4e4a43;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb12922a74c67086f808866c3a55da3436ad29e2c16cdd62b2ba4a61fe7c6cda3636fbad461c37cbf78ce0fcea0e45ff00d22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8591e85c11335de8184f41816745deb0f74a8ad14608e70a716b95b58f8f3ebc18d4290180a8be7c54a40a11c936f1a4833;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he010a0d381b94b50b57f122fd3b97a5155ded8e533f708d53a2ee897c440ad1b707ba732cb762effd9e6b006e14cfb70c305;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he670ff0bbf88cff11fcaecf69491e313bf639b7f15ca39bf52a17f7ecd967f1c9415907a3275479261cfa1f3e57314c31939;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc62d633fc96c3bef61ea6c2037bdb68f6c26e46e1d9d67f8e510642c86a2d89066ae5fa8841174aa3e2ff75afec264849ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f51e03fa7046b8eacc13c126fe66690b098db7294874ce111b0777b8887dc71019fa107701cc4300e221a5641238b93d6ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha816be439efb59376ca5bda70b47e0e54240325b012fe98465f3615efaa34793c051f08c9b579ff189e91ea52f54fc1bd265;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha57b6355516d298b09a07888dd4b80f545e6718e23f7e766b33abf7f161af7f8fb4c65827194c9cb7100e64d3646afe3f096;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb31760343f2eda368c902e2def715dca7b638f6bba73c69e5e457fa0b84f87ef96c3e110734aca0bb341146d5b9faf6f6da2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6cba7f13be02b379d7b14b688f13ea85baaf1a1263012815d966aee4d9faa9d8596f7fb7feac49086987f57a6a501d19134;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e8e3abfc47f0036b740f4b25c694eb3df90f73b9901afad3c396f89fb1288ee7a5139916fc0160a9d3b87290ec4097d4ed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd02213f3335f7e96309d6b044704f7da110cf5be3643df4c6a7f7a78a93d8c26f2afd732fe84c77c7ba0e1c6d5d6e9fbe074;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9bb899e8086171f9a15e5b4ecbcbb3c54b2aacfdcab04e1ad4f6708b13735367892b75b50c2228d75d589c43f518100eed5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb806e58f5ad8e1c2862216f74777e48953bd7dccf97021e3450b7c2c786848365b49e14372ed3e346c03f76623436d2b960;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4cf4cb2910bf09d5d226162c3681d24aafdce47c5e375a42b4bdddaf8f213c7b154960615b4af6c50971e0fe54600e8a2c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h839d6b4a5d0601892fdc75973fb615834d063eb480f817f7feb51f99ea4a413cb0d0eb76259c003f284075861ffbad68ec66;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h108e60933f7a09058a2d02213b60ebaa3b49f19095f75b44053063dd531544b3cb52fca58eb5323c64331bb3e87d7f70d212;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1ad9bd99565629d89b1814e93a0b68bd14669f2014d52db8c8f73cdd415bf0d89e47233be45566a10c26f104f24bba557c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bd4bf26eeb961a84a6cd1da9a641c878bf84b707f12c3ce46ba6d44b4e8ccbacb106fcc137ac81ff45fbe324b54add30adf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h518b1f0482beda198e6abe2ffdebbdb79d04ee0c60ccdaaa6eb329e21113b3943c01eb4f9d694cb69dad212c077ef72eb60d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3c8a72ae8d83c4c6f49a5124e0b6036e50eb92b05ad427c8e2f8cc479ff39268e388186b2d89fb773d5ac0e401d9269d1d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8bfb3100618ccc1f107d718caefe3ae2f6da9f71cfd8deca4a7ab51a8985ec40d2fc0a236855baafdf8667bae47fc21663a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd751622d58e0422dc727e0d36a0118c4096ace09720b3de1907ae870c3ac1cb1f0f585b91f8c9deb059cbd4a7294e572c07d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c4b363434d32145353fd8019c2b16fa7e9bedce704bbd5470ca2038c7037e0b6fc3533bf9563216dd2fb135481cb50ec95b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1105fbe96c3c9fc6148e0ec6f83c25d5024abe4b2a52ee07e7753c433ed758ab8d6b587be1be4c12e2d18163903b9cd3546b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h91b3e60acb544b4b7d41a8af951dbabab4f168f7330754b4bcff3aa6810ed5ff289aa5037f3d5bef1c1c805a3acd0734bbf6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f8ebb40c05eca777f56ce42672887e938a0baf49c9acc2b44fbff22dc8a2b0fec22c2d3c5a5452e686ff6a45c9842d532b7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1ec173fc0502b9fb47714a81d63fff53e9315dc1567c7845969f79f9f4a167c616ca81ae79a7073d5d4e9642d0d93e00b82;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a9535e9289f07050bb5ff66c2daaf6339281b12847662223cab4f8a3555386a5dbd832524fda6e1aa7d5a3ff00645d9236c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had50eb370206a405dc38e9288b70079a610fce0e607a424c272e0e5b4ecc8d2b829cc4b968e5225e0ea8f1fbdfa84970b989;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4593de9c61eeda3fe6968dceb47e974728afd11682bb281b873223025b906d322de2a0548c8dbbbee38eec90eca51c97d9c0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h683d8e1d3baf5436b6d5b7937be88dd09875c3ccfff6bc58a30341d0c98b64034c2590b3becf94e62d0c70c4d1a34b97321f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe70a872a64c06e9e47de3441b15cafd440c20479965b10d3b3c2ab02ee5ffab96f4dc3ba3cffbde9da5fb60d9175e2c3524;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9542649d1e1ed396be67ab8891f5e6714d8148f96df3654c856df589431084f1e6081edfe49b70775ce3d9587d8a8d9e5962;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9b9b2ef06895dfbac1d7a23de8a7d05f73e293d2b72ca5b4d30a5de5a5aee5a759e4dec7acc724198a520e156428ca2bc87;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdb7bc95dc6168580dc1b8ba8fbdc0511c9cee2fb782be3ee6c27659685a076f6798504713f3e5aa8c8f822af258a6dac819;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he643d0acf5320c1025904bb4869bcb692d9bb0eb678b2ed39f5658e1a9d83208ffc0bd60477e8ba8702eb794d4b51a8c39ec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he33ec31974bd9711c9a245a5ae9cb572f3987aa95db3e9104adf6ebe419704542239a7cf2be1b92c7389b7471cfb61f578f0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6cc67b9b4846b23c1cd23f9a12110da8b3c0c8efd91aea4bb5a704db67ee737f8cce037204df60726ffc4529d1821b268f24;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c30b6da5f8f4bfbd46dad6b26917a569fbfed365e9b2b471799e0f6978a8ca0b0cf35aa736170604fc61f4816ac2d8cb50f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46c9f69c985d03244969df6d5d0ceb53cd3c227e0e57244216258b2df87200d2d9206f248b81949e4824545f7d6d770ddddc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68a99335c4797c5b7c4a2285c47765ae889c6be0d54aa414b972daf00cb4ca08c3f0ce5c0eb97af69d514fa8b94f80e57b23;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d945e201f6a3f804be6e941221e5f2b98942086f1cfbf65f04f7cec97efe2b2c48e6c89cfc3f9a7da27d95409b9e15a004e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5cd8f8489e2dba6639e754cf9d7a7b539d5b0ed7a648647608bea20a57fa487a4f4f8a17b7fd3e2ce116c3d63d7efeedda4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf05bc298dd126174aae4cfd72c6590174ffa4bcbff4b8b4ed89cda93e66809c2ec367b499e036968903858d9385ac7e96842;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2aa49cc91736410830170522fc5fed1d0bb85d2a0bb746dc95083d658ca50cc8e3770552934ce56d20248bb37039fbf98980;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc950881de008b2e98d8b54d7851f6117d1938e78c50470a977aac92e240c309cf4c96c7d0cf6c33e0d7240bd804f076d2d8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29ba3fcbff2069b91ead3d18bbf9c6df9b326d1cfb7f497c888483b4e29ac6247ec1b4e0db49651e090d79396373c139e4fd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heefe4062a118f6cb8515e44e3876460137a208eee1619565905ad9194f9607ce550b1ae79ac692ab1c673a66ec70dafbd9ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h470dcffc73583b45733e091e5b3777ec479b0f9ecc2ee1ff1d0676fd7d409c5ce682e84cb27fab4078cec73500e1172143eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebf074d6f9c825056cdc8915c577fd30d42eb544062b2d079f65b5c39a786c923acc8b8f8efdf54d117c93ac251ff152fa08;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ad20b9e19c88413016fba65b74d9f3e876b6ebdeefcc728dbc437dbd9a9a299ff0dca59807faf7ab91602c00e7824b574f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5031a91e351fbc2f6568fbe4d217d944fda9c7cb5d4d247c78cde4dec1c0467e10a47d17298b6a26e7660966ceb56d91d099;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82e2b2fa0340f08ee94efbd5851545ae97bcfe45e9718bd39772d8af015b89f92c4517aff8f5df46a1d77f4694f2a26717e5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h809fd6d6db7a994927454be471e75c7d44a024de751d959e24ef08c4ea743adb0efd80e15c4a591e4c02bca4f2db33a7f4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he966e23d530106ee653c3fbffec90fe9fbc579427edf8ba03c0d7cb26d48a67587f72bc27e9a795d3f186550405bda84490;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcba2bdff7504e8c5506da9ebbc9e1b0f7d1fe809b0ddc395e63c1e7285df13a2b01a3df9ff4eb1a225d8c31834c7d26afe0f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a9992946fce1a1548ccb7398be79cc7859800c905d0414c10f3a99e3562d43d60ff31985cf6994aa911695a2173f9848030;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b4b7a46423f5cb57ce9a6338c1932794124a9ddd974a406d662b16c4f3b185f9a54ea10f6a72b0cb1d69bafc5bfbdb6df13;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2b8dffcb1ffe1da1aa7b6c3e2ef2aed8c603187bbc5cd958782eb15f5cc468ae795c7fb0778fc42d04976d49212dc0135d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a93fbf43bee33f90ad6b688e15b404b55ff745c830f5c46f67db8f7e9b94c3a13b67fa5711b6017edec69bff08fb20858d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heee5e809f2095b4d37314c81887d2e5886d6845451237b8c7e93cfc41b8a80be3c6427bc1bf2dd12fb07c6011449a0fd5964;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha8bf79a70f2d926b36309c6136c63823029a05a68f040368563b5566ad42b193daabbfa83423ecea9b3b9de50de5b143782d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee7085a8a14d3daed55ed85defd96ba1bdc81c54804693e62dd39f06198303a606f37ea1638d7e3225f734da9c6953f4eea6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e94b44e179c5a7e58b5b5b1fda9e08089e2ba3928dd62ff1c72f72d3dc36d04d20051878a6adb7fa0b49f0d9ad2aa0e1e78;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10acee3246cfaf98b2bc6b2b4b8a3a8128e6b3bd36f8a9ba27a61af804d8243bfe9bde5838bddeab09c6adb1adf389ad9ba3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd7299083a2666908ae791c002205907f7249b2b5467f9c0e2b5f3a0501ec50a8e9c0f14abc7e2660dc2fdeb2658396580a27;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b55c49bcc1d0430e970a7ebaa709e89af3bacb0ee721aaf0703ec55ac716e64d73536f9a5d88be8dd16c9e6d15ea37d5035;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9dfc5d87272bbcc9ce1480e8c3370b087bc0347840370b7ddeea5480acb21211a1692892bb919612beee01a032420d52958;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3546c3c31f67b71cd82ebe6d4cafe61bebb3800ce1179853708c27a92883e3cd8bbf25476bdde330b520f662b9fc920c96c6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h10a05f126bad268c325d775dfec2f7fcab541b9c12d1c215c23272d7d5b531f0383bd3e641f04668541af861eb88659a950f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h641f89d464e90ca6e3b8cb6dc7f19b9c4f5537ed1d02f63fae394b2a0be5686067fd7255ea7e1f8d962caa2996a17fc7507f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf021cff958e8b108fd22ac1e90754c5eff9b7943cef14a36af3056d4f2e948fa6569e94a25d311acfe2744b02b60e685d8b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ba09ffe6116a48a9be4b8a362ad396cd4ff39773615d2f2cc47dc919dd3aead24c9682935292708ee03091e5e99396d878f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33eb9ac31ae0c1a460c779f633508d92103ee9d076feb479a3907c83e8e21471e78cb21b9d0b840ac55e305912722a85f44e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf55f1007ae12b4ac94b1bfef13d62e632802c6dc340d4f660aa6c7de4f4c98a434e3d8196d25cd7a6663dab8dc4e904de0da;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h152bc62ec5bfd4148f4acd0949a145ae199af5e89f8a41f1c639efbe9f06153f27f3516374b58996e50e47003e20487b23e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5ad16dd8ce2cd62753367164fe9cddceb1e90eefb8c10d9e2753d71259b028c2658a047a1b449e5a365ffaab97f7daabab9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb11a731edf8ac70fa21cd74be8a267ff39cbed4fc3b272f697da91c92b75ac6b7b8fdb9ee725988ad2a125fbc4f2ba9d7d6f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h662bc21a765f86e5c0c5c0639ee05edc1936b89d544a473950174a0de29d29619cf87b11a12e8d074fd268cb67a990af1d74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2b9c9b936b5d20240032a720fe266bfe3e7b9bbea713d4d809664c3bb306a21decd7c615550d830650fe302c71c4b240286;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h669d9996fe7b049865c1e4f39ad6033e6efdcbae1a01307ccd66d47daeb85c2c40acf929b93510b3c1061d00723b94f4e223;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33ddfe7c42024493c48d43b33af2bf2d1d9a5d6e3723c2dce520c49ec6f8d4baaa616b753b6c1e28a8da3be91783b1c94a9e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb540cefe0fcf0fe216d4c58d26547141169eece508571aa6f66faa41dee33397b0a983f298a1548c340ed5c66d03bc0cecf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc180473f8bc37334acdfb36c44d94fcaefe922d6e04cf671f5500320a3b0b5815c39d4533b2cec9529dbbbd4106dcae4f47;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41442537def46b8e7925bde38d40b00755770228322bbcc582e44d5ae30ad271dfc71a6b351b29ee161a17a9b519bc737b5b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27039c7362f2fd9361c6a854fcdf4466886dc97fdbf0f71e53bbc76d851ea383622eaa1041a88d21c211039169b4353853c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5925f1b20519822cd4d3a72803fbd16b23cd82d7cdc2e69e1d9db35b2ee90ec2b788858f973658b8753d0a0c92c2cda303c1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he84e296990f8a803321f2e6ecdf3ec20ac81b6531e206c28c6cdd4ee28e435492d43c6467b17d0efada09679c204ba193c40;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea5ac675b5757d18c6c8b09fb59c18fd0baa176ae43850629398a0a73e95b956e13468ef3d0008e3e52d79a5535df29ee56b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb74db14aacfefa9e503cb8be64e63dbb88aaf18ff09d6cfc4bbee3a34fd7983290ca595fcd3130ea6e3163707a8f0431434f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha93cb491741d5a285c6ab33a446d3e73d25b79b619211c50efc3bf08f69dd9b57abd42311edea1dda57261e4d6e190bf3cab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9fc0c208fa270eeb525334e6fe4ea1e28a0ebea0028af9b9b8050901a6400aff6333d70126f1fd9f0ce515306623a6dd1b7d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb6d9c3661934351c79a25183fb0857757e7aef0ec55c073d8072b4b8932b5caee8b3e32e30fd769f8bad1aecd3298557d9c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5a92586d544c05145001fe42655332f5657f005fd5d57e187df585552c839742d6a6ea451e6ac2824abf97be6348972b470;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47b1f34ad641bd864ab12ef56b1a766f7905574de1eecd6d189b4948351695de3875c0662adf36cd8c4976e19dc95edee461;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h874b49b535006a54559fda0b480e554a8a9f520c141fd0928eb9882562ec960e269eb51548de1004d87f1bc955d5e0b5cd5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f22f89d00f2f946f60c1920b9bfc8628f72025b25a89610e6c147ac34b5e8e2f31e301947f61ca78fd998777599ee4c0809;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf996b78959d8a7eddb715116d1404026018dbc40dccaefedce7e928452cd9b530738099ecf4b569fa025ac320aac756026d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8273f33b912392892f3f970c1ab345ea7214b9a36fcaa3268d23844db12914c0b36279328cf5b644e110a948a2236f673961;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h728ddcd1d2a374550b837a78614862f65bc713deaae99e3d783de30b7e6b2f0b410cdd33aed31396705bf6eaf6c8f6268625;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bbe1b1f9472d5b8a64e6f71a5287db3b05877e3c33ab4f55820926f9e914f29befb1b6f6485cbef5515d1081580628638ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb31d1ed23ef44148064ee290bef7039e384b21ab887501dcc628c2f8a4518a4c002de665747e6083f4097226ea50aea69e8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76d35140c447579a4f1b519bb9814b624f11d1ddf7d008510260bf7f5f3d123c98e5b824221895899d8308ee36b5474cd8d3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'habbfec0179a5cd6083415331240d5bc7589653e2efe6b9efbf0a85ae2c271826110befb08804d065e689f4de5b5ef97a9faa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h698c3724e8e5db49add9013c77f64a18f305dfd6ae566234707e329c74989fb92b8b797ea5fed9601e3edbc3a1c25688cd2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4238edc0a4f4ca5391dc7c8a6340f1f2f867e3e482c24257b6630f3cfdf0e8cb00aeeae0f4ce6f0211136ca53a4b175d2a07;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ebad0da544960aeedc6a92d55aecccd37b9048e3c08ac423cebdfd2f49d6f48177276c4410aa0995c66cdb91c7142333bc1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32cd0ca0d19fa43216a8df8af4541bde6e303dc6381c6f9ed850047db30815af1dacd1a3205e932f087075a5ccc7bb76007c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c128881e0b098a54e4e64a532ba4d0176bd82551e617adc51e8084ee6c9fa2e6d5d2a1e22f433542566dd28a9c813f0cc9f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26e6cc3ced64bc05833344490c1f9c73abadcff103ed33e4167f21ec54dd2407a62e257ac3b4a4d51cd211c28db855caf82b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84983701fae9457298cf5505b6c28b791db8ccdc638f75ca25e0f26846ed1c01cab7e393f054323610c624c4adabce98eeb0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcbc37aaad83fb2510b8d6b371738d84edd2be3a835f6817f000459e78e4e6409fbc5ee29fd476240381d68eb3d2714d595a6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf62d6e9652e9358a6c395713290e0ef33287b8f881a4c5c44ab1a8b34631b7f2222318440b2274eb5d6906abe7c771fd56b6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6231b7e74e539732c7d99b69a017fdf17c0bd799f0dc7ac450c20e8b55b7d2508a9a03623ecf6a4a68d13af2643c2e5f19d5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he64f8274f54d878d4adf746790a3f07c9f02e325c64181f7ba3ad2ffde02312e33be786f47ff284a2452d86b8d339dff893a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3554bc5adacb7e7c5ad9e4c4820f3824e58c8657a1362b0ad827a5cfdec0014287308526cbb3bcbcb0f9485ea749785b0d77;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7671d44a5f708fc20c364edacff37b45cd006b6a5abdb4aa58a0fa39f2c4d5263ec759ff84f9c5f12e41fa02b7aca353b6e1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ed803ced8aabc0d44362d8ec019eeed396f382bc8110f66e428a61db81d47a17f1dbd62207b836b287a8c19994a93592713;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e6030cb423c95bd64602ae1e9ee2c83e81251ef72b8d51b6a997ba3bcf89a5e3fa6535f3e98cbe4486b4e6a6b2d4a010821;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h739cc1e1e1a8cccc9c3fb7c40e4b41d16a83b3e0754133f5e134c3e9478dc8da90b36f2cc7a2bd0d33fe51bd507b27136be3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h467a9a14bd00415c4f1787a1f1b6b2422e73127dba99c777c2285943828009f2608f3150307289d0f84af0c4b78a3826ecae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88e9ac4e52cfefb7334d7bd1840d4118c3acb1110d287bc63f1f24afa0e86163a8c2f99861ccbc00b220350c2456a028f275;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1421f73de40675c29234404dd740eeb2253abcdd563a229210a1ac91291b22320d583ba577419e033b6258ee0d4b8b22b687;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b3045965000a2d35b64c2bd5b7dc94bfeeeb6364e719b1d7ef99789659411548b82c4111ea4bef352328eaa0feada6e1b90;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf355d345e036a469fcfe80e1a4c0da8ade96386463a5508da5ebe6dd3f255b61c8f93162f33daf1ea65d5c94ac6748c7129;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80eacb04efd7da4af2ec96712895bf42f268a376d539c9ec38aac96d5efadb4b59975de4a573c8bd82240958de2016040894;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96dc857ea2ebce33e06a884048dc4d587dc02442d33aa9a33ccb07d07c7c635fda94f8483c45873b93b74201435a9ae26ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d1a7d8afbeab148240102253649088eb2d1d0fc6c5f0d87394744802b2bc20f498cb7c6dbcfc377c8e3be18eb3f932ab9b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a615701df2c55237a5db255c8c1f266fab6611eb4c80929fe89ceb87b9d6111115296d728190ed83f1354c2b161a25bfc2b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f6e10512353e9d0dd74fa85b96a0f8ce988c884f3178253b4d5e59613cc8ef89d6cf01cecd11be5a01c17652cbf782d4f9d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haac2fff9eb2a90ae1928a91a4122a0aece81ce1e455a4309c0ffa1bf7ee46916dd35a77688b525b5fb4a1d7f07ca5c0cf01e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ea42e14a7220c7339ed9994911e3f6b0ee6a018bed424852e03460c5f23205f735e62e5868914a7bf43fc0ed63013b882a2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc8d13db1d0486303d594ab751fc887835537af85617c3b67e1cf104e2e38fd57316274e5f26b8496e950963b010d2264ced;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce5735e4c8397b7330269b3ddf212bdfc846b5a723c82cce2a08e5a802d8305506b40513ae2d986c800b4949b2c15ca0db27;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41b0996cdb52dbfe7f10a05592f0ff90c47c0e9ea934f863d9a795532682979adb98a176a7eb0a5814e430f00e5ce8fe607e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b8e4bbf071a1b5580fa44a87dd264435f609ec0ec9b2656703a277fa5d36b632a91f46acf9b1164e12a3b7faee0219f97d2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44d0b6c41b0b4c19f780b5bd0c92921f6de37083767352b1581844ade0a962b5f4e4bb931c51b42063d4212acaadfd3d0a94;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h282561b02a572ff35d004693adfef984c6b31520aab400bc54ac6199a09548e0ae05c43711d0a9a224ad89c268e75b126dfe;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h574c71948d8e940e04eaae5b77e74e3423bcbca273004d1950f808b13881bdc3d58b5bec9af9978148b4d42996b1e4a8c7d1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d586d532ee2602a6558fbcbdb2d2c18c1aa7342c6796f5a7a4162993af075f56430d5e91ffc64092df2f18a33ca2d5ac6a2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44f65224020bc483b6a4a1125ff7cbc2789473020839afc6f57a16f631830c1663f39e4844349d43de1932e862ee06405056;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe016d0c11c261d88fcb66887badfbf8b10470fa2f30cd5a6b1359c6fd73429900eef855a57edfdebfb76cdc15060f6d3ce1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94c89b720c20cc0e658fd0690c0d15aab5547c8a1dbb9fb868f814e343b225f37d1f3900cdba6032f6be5b4d5441cd8fba89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84fdc1752b5c8f6e414dfc3ba63eb9ce455cc767930247382b13947066bbc62b614032210cefe13b891ce5da04f7bc767fb0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a140bc8bf88fb94eacca17bf6bffee379f081100a29df3509a76deaa04566adac61d735497d0895a1c39f71ba08f3d62295;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacb8b5c7fbd4b3791a102917c4f7f2d7df85626dc90bc23d7b75bad51a6a11bd40f2a238526c9e060c2c25fe9cd66851a0f5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b75b0b9a19396a1211183a3061c56344b54879155ca7b073281de552923c101f4f89279ed1f25e188c8ae57ffd0d72aba97;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53d8f17467438fdb83e42e1433750d4755e9a5e8e2b785c2f224aab6baeab60388ce9bb83d5c723ff4e5276952f126ad3c5d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24a313eaccb8547eb02444f7e971448117b38a5067eb7c81501a8d8ee542a4225d0ca4650b3c5525cf7e1641bca704721ecf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92542f192c889f6f7b498a5df55d7d9ab97a36b67ac764abfd82183588830eff6c127acc0d3fa866d3b5da1c4600b77ac41d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16486fc4fc8583544a75b3b02e1d97143fd879710d14926c14d58848e3fdd15a84d2c6516cba23b74c2088ea4c8f76eaef22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d1f402db724a28aafc367c22b4017949b88b00c820db78328c8f872968c00baef3c0da46cbc1fef40407cbc08158971e7dd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h922ef51f6bf319984779b261c4049bd2ec9ec3f5dbba81927d6895f1449787a696c51862192adfa6ccaefeab2b84f0a86d29;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7821d5f57caf6bae2e0a6098b3ce1794468cc7ee012885c94c7a0f4233e9e6147cf04d47dd55dd4e29570a0ffb18c4b8ba89;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b7039f14cfedfbc867fc74da4f7680ff255126c86eb3ae7d0860e39eb1fd2a3a29a602944163814a7ddf98bed6f1021a2e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdd7953d2466736b2fc67876e2e78c1f432314c329256dfdb6bf70df42e27e393250f7a5b127f33df464a52b6ec47c83ac45;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4f9a37665d23f8da15cae3b552c58b3a53b808a34c7bfacfd6fe57b5507d553a7d5a14012331d583d2fa31b750c8087a399;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3237cd0995783a1d38782df85705f5f205642f6a29e4e1ca203ae7fa4cc62305f889b946daa796675e1ad44c9d76b1fca6ca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde1cef6c47fc152d828463d811f0b2bb6c39e650b8d48d11fa2440c2da77bafa8a8f8930888289a44c86bda7a9d76c04cf0e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb52db844376fcd61834e98cc605be29f9aa010080a65ec9b534575d21bda257568323a833465f517c5654a5fe3d9bace846b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3596552ff1d723ae8bec4cc63491b25f261a4e4120e05e21c8fa353c4169a4d8cefe72c950f34dc9bdc832b28b9213d63b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92a1f06e9d3c4f88b5cdd0dc26e695727013dbd1a33bfa220d21f7df6f739dc6eb39c484871d361980f55633823e28c582c4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h75f7dd9dbabee0d1a8883235a1f3567fd8d6ab6d117c0614ae4b52cd17b55e48b114a431556b0cb10aeadbcf71b92a88e05d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c5eb3635052cf17a0af55fd1556d9e9934c53effa94ee36634a9763398bae99d77a76fe8c4ebb8e7769bbcd9f34e582cc83;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5403b8a38cc5a1e6642f1f09c41a2c361fc1233d32c7f78a65dfb2c5ad78c8aed26db4fc1032177f4a668ac550e7abc21d4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4bc02cc5f512c7a36d4c2e37e31c39f1a9f065ceac9964722da2513d2f1f563686d363dc8057828694d0a7e67f359ac1b858;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb091f4846f0c29aa7c9dc2cae9beb446c4af2fbcf2c179257f658865baf2d3941e4706a0fc1d11ab5e2be282757fbe49ef54;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h76442afc4f9ab6ed4a55d0543c8ddf5188463963a2271241499874793e2c606542630d8eb17415f91cea1e729f72445cbd3d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h306d7787cbcda2fb9166580b04115a4831d6fb17891427fc0987a6f5b4522e4f0b17fc20bf187d381ea23b8a8869a17fcb84;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f051b00145bd00ef26b3f7c2907106f7a4d3c7d9fccebc57d499ab59b2ab87b075ddc02f0995740bd04644f7577b3cad165;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31d94403cb36799731e7e0d7c7b011f573c8edd7fa1720c511170123e2ddc0cbdbb4e535ac8a9a4bdb0fb5a43c21f8bb1ed0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7e5d3f0e3bc01f73758e56ac0db2df7030a31096d6d70c36dfcccdc8263f634e43b83a5aa28d60779248808e8bfbc82328e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef2cdf2e0ab5c9fb816cc0a6b053af976350d5c8513a5203bd05f9e2238d3a2ee888a0dc7ca7a4a7d1fd5783ea55394fede7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69d0fb9b45f191e644bf62857cdbd0b420c5aa6ab1d92921756adb297f761e6167fc5958b6214cc065eff045a36f8a90d354;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5ae297430fbfe56028c808fa9f4ac52bd4c2414369c8a1ea75f8c26a57a74a73cf379d1697e12bc6564479afc52f8684b18;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2ebe8f5a35641b80301e5ac75933fb182965fe94e82ae32e56630aca655f7b9a1bc36be8223d5d06a089103552b0748ecf2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h921dc029b5a69b8352c83af92b317834bb931d464ed13223cef25d9d727c6103badb983273455167561f836d8f95b2eb6c69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a7363c90e62159bf3b85561547e736d73bbc23044e4812d140a6b680d39c572d2a480c0e6f18c502e10fd6c3ac0c0f4d164;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35a1d3919bacd41672c5bbff5bdfd21b3bea7263d8bbb65064002a2142d734f880f9620e9b6c5d4eb4d51ffcec310ffdea2e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc98be4ad23452e80591c1cfbd92cbea4a1122e5e98c8229d6ef44f5724aff918ac6d6c018e4b64abca36e3f4aaff9f11f039;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb9471b507dbba52f763dc53530e6e392d86178af30aeaef17840db853cefafdf5df233041ca4d5d384cb4b175cfc77e4b46;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2183a8cf8472bf26adc584a22c50b909071a947b0b21a8f571818132f7b49111aa88e6682d23d1ef7b9af24133cad3ac45a9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45a5480f72c7f0a44104994ef843a7ea3e2e0049232143509d5abe460b0a41ba395c122fcf1ca55c533b93fe9aa738ff03c8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2559c5a36d6068bf1300eba7ec11083346a7061b7e45ae20ec749762507083a927d7c6908ea457186136c5d918e429b8c2a3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf635c9e1896b21187675941c8a3063c41868020baa79a3da7aae0489da05c167df12b91e53b00aa13306371c76b8fd0a0a17;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6c20158d901e74b386b7d5dd604459cce983ea7916a2bacb39463920845d049ddddcce3d9afe2125078ea2edd09a139b12;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h157d5e8b584b1d9f4cb1cac2e2ed551df3f0557ceaf9e6f9760724e2d4f0b317bfc80d81d86fd0dbf944b4031f504002902;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc74a816865d8265ae071a7a9ccea9b25846ea9827ad508b89653182048547536da2ed4d547306bade305175e0d444b42001;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa2bd11dca03a750f2d09ae1fc5b74e57f32f1fd5555cdb89b99f73637cb79354121b8f461a890cbc7481258c71115db96c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e39417d53bb227abe9a9a630fe2039e370d861dd8f869f85d32ea9d8f1cd6a86f8b6ded03174389dc277eb683963e843abb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h91b9169389a094834a359528b8d8e4beb98d0e6a4b3c65c5db97e32b26dae4fb84c8bc9e7aa436a8102581a7c0146b152a69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc84d28f0988b0188f799c002d91a4425ebfd65a341418b959c3a910d526fd1dc85d7da7c8a0575a5899728d497abbfae850;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20c75eb0b8387d4b570fb80570ad76bc365f78d4b0c690009e89e3bdac87185b52a5c76f652823ee077926c01cddb51abbb6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d739b11e4b07c2cf14789e9125a926b02781396e1351bf022741e0151276a6ef654e537f596ad04cfd3b0c6b6e631bdef64;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8257da09ec38bd6179447500f6b2cbd47cde465573fefef36b245ec84abc2d125b6ad9485f0ed17331e44054cb626c8d516;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ebddb71746e54cc06734e96d1179df85017d46450a5c5464853cfec36c2451aac974dbed891292a4a730a1f5e7333fb358a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h390fc4ec3b88be92ae389cfc08ff891517760ded68699eb5fbcc1e494887eb1d8b6cb94ff0bac97c98753600dc06b3988abf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f2a1d0b0537281aaffacb72c78d74a435269fe044c51bce9e98b49e744c339d93f7fd1e6a762d2a50da734345e9a768827;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5642519c4f0422fee69ab4eae03c6541aba9d5d70536e576f75d601a650d0cf4dbcdd469f88adeba5f121fa6c1bc579eac7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8607c2f0e6d510aa864030ff15b066977bdd744b6614acd4f60796501a10eb05746b8060108cd7562d594f1169d77ef5ca10;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ea72f0b640286a57dc5c4bccb29f4b764c030bd66373aaeb0c20818229db005c555504a9332b74c2ae5ecb06ce3ca5fd032;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68dff86cb52bcecd6be10a30cee3252c785e6f21a1a1cffad764d67ef2915f189fb2c5a60f6d1617d82d8e577ee4754d2719;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47d0ee67f1192c40636a27e006905f8bf00f864a2ef1f45238f16139aff9c843a8fd4fb5c003ed41e1d9ddc7194803eaabac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcfc5d18ec445d0f14e112d8b7a26829531982195caad82195e66c6fb519055ef2b000c745c6331cb4ae937ca1641befe5062;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h47e2a0e5005169ecb74a4fcd0e3fe487363a004d0410986ff97f688798e88df84a21f70fd036052d5c31276129e29440763e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fae74cd7a657155b6f361102cfa952171ad5cc496931a7231c1f739109b6114e86219fca9c625bc44b30db843f57c118919;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35bb7d28422db63ab02a8d68a0db3c68b583f13c3f5f5e28ce1353d6bc614b088036ed56ece3bc878ed93b294f438be3f2ea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ccee1fae5578241661b98168b42e1367426f98d45c0bd916a709aca9614d9a61434d13ea72c66f0b276bf08d78709640a0b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd03f51ad99e921c1c296a8c3198ec8b49a3231e1776beff8a7cf0bdc744e2d681b3c48923af3fc6b37610ccfa76b656959e6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee769287bd41f78e49b83c080e5fc0d3008919038cc43a803095888857590a9dfbb87b265cf9d5a18b189350cc83ad1ca387;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6e7ccc2396b2c711a577f04112cacc7961ca3940bc2dd6a6670a9a6507c491d548be59969b74c5e24b767ab7d4e772322ed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9cf0e1a965d136f19b1f2628f7f14f09daeb4dd8a5056106891462fd43b3668840a35a112a5e4919fa5b1f908874f4ac7bf9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f20519c9b90b1acb683b46bafbcb78d93bb3a4cbc308cd9b4eb701185430ad69e25c40496d627845bdcbac6dc31e987cc3f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc5ef6e8ed8ce3cb02a0c0cf1770a8d79e9ba9024b85b63e32ce74eb62e5235955f78462472d9f8a612b0dff82b48b0846a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf22f13f569e76ec7171a25a0039db668684fca99ac8abffb2996f8ed55bb8b729d92721bdbb4041efed8c8ee070aad3a3ec1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99bff5fd514889cf912e68074fe344c0aa3e513073d76c71c7a92c4c2d8996eb5a269c8cd5e4367b531639ea876a1fb8e78e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33b8121812df82b1785b644c875abaafdcebd9e5a732eb3f37fca8e57782ba15e344f650922269842424320954dc94c28a3f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1518d9ec423b8826454b250e917c3327183dc0b14122290ff21b436907168074ba39f03cc462fac4a5aa8f90020bdd8c4c0a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec7268225b61c9229bd799c5dd4568ad4e620d1bd30a9e470b9638d3b6bd350abbde8a43abc94b5544e1842f0d9a992e52a3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83fbcf8744e9fee0d4ec8ee0b3426c638f21ca48675dc15d600d0e8bb701503237d7deef4ee7adc2b15f193c658b79964936;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc21a926a6a21e58add41409202f0444d4bab44b2d2f7d6fa31deaa0a72a97a1df1df68406c32e24fbbe4145955d3cccde5cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29e1b82f3271859ce8a2eaab1cc05cb79cf27c9506ff2b7db7bbc2d73bac518e077593c696e985269dc7e7830885c117783d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha18d6a98f49376ecbca013d0d1ae3fe90c6ac0321a369bd091325b5052189ee50add9740d89f33b1a9aed4d408ed6ee0f1b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9b324ef1a03f48c510597559025f65a1c2ac45fcc72119b7118a3d6ef1b54e868e9e6fbc682bcc7d36eae3e83f00e458ca;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h796c13a7b1495512aa41dc004ede5d8ef3fed16e3bdaf38eb9021dfcb6838958419503e0f7af263b66854af35bdd4767bcdd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66a2a7d62e30f49ed7bed7fe463283cbfddaa8d13a25696f892b806f46774d31e8d8127eecee88961596910ff5a3b82f53c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62c8e12c2c11e14b1ae0cd7c9ae0166be5347817ec2ecc3ad27484f367a738f676a174164be9e3cc5ffd6bc3094e8751507c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he965c3f09840fcac3642a13ac2463aad73ea28445777dcff4a81619b5ebd72c2f49976731603b3bc09bb6ff93324a934a5df;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85da6edd4cafe015dc3ebe3934aded7808bbb0436f2bc641028659f9a006b5171df240d1c55b3fa76eb4e4cf727c6fdcb068;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd7696b7d020da057495947bdf575c12a547241eaf7026291960deeaf853b8fe54c9e5f4e58bb66fb727e5c7538948668af2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12c667572bfd9dbfd6d441bb0681f03cd6b1003ab78e034c382c2f6f46eb88248fc8dc877b98573cbee0ad9df7b324417bbc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h753649840eec66b07b298922d14fa7727cf03e4b0e60274a4587a88b062f8ddfa18bb0a6df92dae83c8085d622f5d4301dce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ca53046a869d958635a31f3a1907fb8e13c149eec7fd9677acb67448fe14ecc8659db87a8d4d2c4bd25de0bbd308f65233;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h530842564623e1faeaf1ce5be5d01c0214732827bff8d1bdd15897dec797979c001769aa90ae14689a2ada8414fc8c5cc138;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf25a3355db13dbc03271aff61fcc4dd14a0b1f0fabf729e1e78ef69e54118a395b455515f0a5ae8ef33d791e8e3885bc3172;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc05b8816cbf98f3daeda3f627961c8547039b2ef446afbc68184cb2c1ba21bdf81af5b8e04dda235edf7b681ff7759edaa2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcbe73a7e9f920a80a3795550a312154a163fbe0be227dd03b43c244de21afb72a62ed2b7ea977bb26e95ee2adb0771e5c13a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h114b7578445e0d27cf25638a95aaae42ec39be987c4fde4ba278e5062822ec41afe1ceb7407bfbf16029d4aafe7358899291;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7452a42c392d3758b050c320ad90d2f08a60999643f45c80f6b0de677f1547804acfa9ac91bb307cd4e40e2b5a2fb53ec6a5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9af7609519c110e0b1bca230810eec83494f07b075712097141658dee94f22f06f4361eb1d192397870b1434ca5806c77872;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74b0f1b4b7740dba1e7dbaa4ebb90483496e752f324854710612d13e39615e3d082d523c45021ac7e2a29c6fa67c76b6feb6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96a82b1ec4d4f3be2e06a2983a88eec86110deaf547be55734c5e171b0c1c048670fa8189f478a376c6d73ac2460b9c4ab8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66e9a70e1d688427f3312b78bdc1ebca117bb6b81fab28dc75d2d02ca380b000b05a5212d63d8bffdf33352aacc57c8dad50;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h423ac626546680edfaa21c61eefd0710ff2b263d49e1175d1effc820cd00426bd37e3f990eb8655777d5bfef80e16162a523;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6cd99e00f125d6cfe42033876ae4faef373e75fddfd20e21dcf57ac016e883578381e9701a9093d919608b54ba16f803300;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd3677f6df722d16d863d3175b392b7bc465bc49d798de9b6e39d1c30cee72137206d2fbec7af8dc4a81ff3b029773837c74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h950afb9c3e41d21699d65e0b444a562ab292edc55fd7ddfe4351b9584bfb1f6c7e8839f018d5c02b5a8c1faa4c5b6177e7c5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe15ca02d2f2c10414ff6cc656ef17bd4056ab89cfac5c4ac99c45fe9ebc8088633cb5c6ac95205a90916ae5361c6da60922;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7c5c49040abff56649f28634809769de74d46ec4ff913ea28e2c26831368c41bf59a1eaab18cc1b5332f010dc4ed8d4bb53;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h988b3f043dfe9d04a5495e6c407b729ce96590721f4ab81886b06e5c79f6e94708471869e9203a873fb57692adff9437f7e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6e8a0b788109a61cbb35b4f51998134dac1e6702eb2821495b5a15200ee28cd4a2208ae6cdafdfcd8f1eacf131992516d43;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87cded374d1241fdbab024cbd8f6ac06b26dd06368e6aaadee30f287ce0b36fa5610e2271d974f0da29c6e8e5c75754b1d27;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he92c3f088b3cd289ef1e7c17f68e7fc8a4dcea900ce6edb789889c18243755162e02db02b548332fb4690e67b8eb8b7ffb02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e51961e0479c50ec42fefb6c10323e6d2504318a5f586874ba8c55aa42c41035ea008bd7184141166b40d8f5092d1786c54;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h252ef313ccdd20f21fc0b96b9610db6dba389770cb10019ae6b5966d183ef0cb056d32632275a51879465d1ad7035d5d61ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65ffe1e3c696f1de59ee94d1e78878f02cd422a9610e5a2018dcf00845adf06bb5a65379c061069e2db901a575afd071e9ff;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8699dee2834575a496d614e8ac8b9d1a7ddb3cf885b7528ab85d89e780984b9b521285d23727672b63b4e507c74325b183fa;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e10ed8dbf1905064345f6b2a40695999b16e4baca0fc966ea668e00693df5d7cd63012493cca8e2b9ba4a62523ddb11493b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28920190e55002c069f9bb7a1a9f6844663acab7543a9ee4b9f10fcd9d3e77e7de15c492dc8d9453a07b7bf217f418fc5f9a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7443ba09ffbfd9c0786d7729711aae4ea98dc451010ec5388207580870ccab907f2a511dac586c241912807d0c1c7340ba28;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he798eca608b57174865c8559b503f10e26df6acf13bbc9153b736c72d1039180959fe0a3b86b9b5381be407664946b744dc6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb767eed9919c4dd2dcb4d9fde1e7965f65390d7c27c77f41bb24edea38d2b63c83c9eeb80682ac770f6352015cdad6b1cdf2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf03a6d532ae36afdec6c66ffd2de6d5b0cdb43dc33162038974e9ddd4d02ce0870b59508dc676fa1b4b19058fe3a0999688d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49d00ce46a45d24a6f39d51e3cec1d4e15b35806e83b1a387126657b3e78d07c6b453598a2b04adf132607d37242b5324fa8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d4455eefd0576cd4e2fadf35a2f29c2958e4f1427dd7cff41107a6f6b362350007453aaf9eb4704dbf128fb64522cbd44a4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ad21bd0a4d5fe3ac55876926869774ad938eba472d0153fce68c9456dd9eec4ab9915de16e4684b69c99af67cd4269f4618;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h833560bae8941bfbfa19c98470e8c8615c4ca032b8ef977edb4436bda1271afbc071ea3062bac82c42d98f41258f4d522838;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6375fe8e003d35768f27b44e0329cdc56a5f63e6342e2aaadb78fac66c33ba98a18595f3b618663597415b4d100a6d974a28;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he859c5a43dacbd969c44b19b9335afe925a4f6b02e4bb5205808fa09edfa39e130b1d8364a1e9f5b79676a05f68e313f528c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5e90230b9d90bd8f913335b084361ea6df805d4815b998a5da3011aa90b1ff133b068ab1640700fedc9a845506a1389c96c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b34bb293b6727d62311f8c2994dabd7472eaa3c225bebbbda1b07e435b8485b9f79e0a206a1984d63344a76c97bb707e882;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5637af2fcc2580ec1eb4a1bc8368f3ef0eae533a1436e1a5bd7be587267749ba465f3d0117d9bc21fcedc30c7c68ddab6906;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a594732319f68ba9f75362cc381821dd2f83b02a999505bc455042b0f02b1cb28107d0e419a17ac57b4f201b141d2821beb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b02bf69e25a058f61eed2d1a53753f7704368f2291b8d2a552a29ad329eaa97f2c548004e578fce94af593e67eca75aa40f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1160592e95d2873d9565e8875ffda1236b9b033ae3101d8137eac0a2bb26fe0b674474c4c7bcf85a3a813c154db4a8454795;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9e91d888ec7443aed464e5d31873a77248e2b02385e6eb5153edc4eb322214e445901cd319c05689200085f36c10e1484b2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0ed171e7da1e9d8bb1b9fadc494ee1179ea7fd50adbfb4b50426c29bf98dcd1b5f6ac3adb6d5493bc28cef3de9d8db6e089;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9225474936d4af8a875cad3c8a0afe2979a3d8a82762294911951be05f3d91f17f5ae4ae676860bb395d07ba1491848626a7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97ce996008062fc5ca73df6dbe87f1fcd6edb59392c335ecac1b0f6864f89201c8b83e27ac925e9e2452954c0403f11dd5cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc78e45fba49ce35bd2277bb932867f84ca7edd385b4465e3106f64e8ee90e94d914ceab925e5a3e7a8367fade4b4ee74433f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h43a962b8924c052c5db2bc9c7fd60e04a9a8ff88709a83d1ff0c8670e1938d96d9fabdc5b52ad4f24e4721489c090e0957e2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17f2886e58307ad3d14507124482d8147e223dc28bf10973614d4baddc02a9b108805b1efcf712074049d2eb3714c0143af;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98ee1eb67d5cb4b28ba8d6d51807a4926cbe8297e7a4d236b01b3c2761a93d21200fc377afbebbc08d186efda813419ea126;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h33861d46b7e66498adac46831344252b33c0a142288b6bb8e9161669333bea3e3cd7c8fca1cbe14dd66b766a2bc09f9a9fc8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4615c767d9e716c99dd61f0de727f64b57010531434787f5147d5b1555f73a234b468eacda982a7a387007d57f765acdc78;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5017f800fdee0861f93bd8ebdcf0ebd0b0228e7a6324d4788e5dada4f0ee5d8d8c33165ef0af83ba2956bb498a544719033e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfea67a601b06974bf545d3267aaf5733523f5ab1a408ee3c59b1b7b6067e1adcc8f318ab4dc66928a3ae5843c50699679015;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h845f56dbcd44d3b6aae56b268e88e0a31db181a2332f15485fb404165f9de33b44c0bae3d8dd33e3df2e7eae47b381ec9829;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51c0e5be2cf9aa129baae7d111ccb7ab31625d149d7eaa0490da487e584ae527965e67994b8ae27afd1bb0aeb9c60c18c42;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5a62157b8d00e2e35cbfd513523c96ccaf16500bbafd60eee9a6112bee8497d3e2593dd65d2a827c817257a05a2be3c9c91;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he5d582544e85aa8e56b4f034270de0accd8ef1d3ef39ec8680a47ec21f9ac886d07e31109e2c5c2b791f9083bca5ed9c1ec5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc22920afb3be9520f9f7ccc9a919a8f913b720b14b8eae6d1a11870a898f3aee529f62e1c00c76c2db61941d8acf16e3eeac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8c3c4468ccd422557e70081b92d2448747a4aed5452064ee5761727717a7c8e6945c659ca6b4d09269e04c12eb009fe54f2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ea7ad258a84c6575b65b5603b447141a72454b5a01d03bbe0b3f6f546a0e67e01518fd6e98bea5612fe94684615eace697a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49719a2beb7fc6602371d8813e9b5515454f1418869435d7dc517c0ec46f866eb606ff0fe599a5acd84a24055830491522ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7944a6d3469ecb40fc29dec80804259f39a8236cabf9709ffdd7b7d809a1ceca44f99c67c8b628cab6bc43c4aa13d654aca8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he77be395b359e2639c4d72db51be775e8e40c3d40c6df3076d151a5ff60d78690245493bb7041d07c18f4f4dcb6a44f77078;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8649ffeca63f8e20d10cb7067f2e29104bf04a5b8c99c33cf0b7de9a151b060ab577c5b05df90fdb5168a4ce68e2018759ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha106fd85d521e64f30ce3b678aa2f06a74ce2986ee50ef43059d064cf71f8fb6c6d133fd10d4e8046fc770e49da3a83f4702;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e868d84442a824382df83e8f8011b632bc9e832bbfd906120c728588138d9b83a9fbe01d96ea52a2c17bfc59adc4b72a659;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heac40fce46d5d8f390fd2a5487a7393b76db78f8004d8cd56aee2876e45dd28b7932c8bebfd9ca5ebc2f1cd9b25c8797b931;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed81cd944f5285355059524e2517c8b055d2e367f6be14bfe8ed00f651ff6e51e8cfe561bf2b26474c3688a71e811a06ff8d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1efec9028aa9b04b4408b04195492e68ef77d06e0838eb2576995df8e526b0b5ac2faf7168ebef9c19844701b1a51a63c397;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b174a30ba0dfd7031a3656475c32da20e2caf9108036f3fc747b14a8b986db426bf7e2b08e65a09dce8f2b66ab9ae7ab6f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3174f99ee9f9b81766b0650a76f1e4c64baf57dee1cc42675736cbf6d11042cfc4605a8cb500e3e8540c2e51c0569fe2e98b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77eaf8db5393078f3f8672acdac0266f5c90488f8b290adff7663fc6734f170603a7332fdf9ebd8c102d170e70ee8367dfec;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e275894ea49f6327f8b12951b6fe564ccf875862316a712627c42732d94c183d735ba7633982d18092700542de9c3b3e12b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h883fb4d2a5639229dd6de3044ee69a331b5cf768f8aeecb9275ee62a06811c24e903dda11899a739c6b71818863e8a0ec19d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ddf2ade1e0f923c20617ff04a8b70c8a3d04d2483c8e46481cecbc732d0d59a489606df80eb8824f370e9c859788435dcc3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d10615ebdfe9492e2e10b606129af9fd643957b35abf5a0c4d2544d26ca95ab23825702ddbf21ff3338a9a15651c35d8184;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf160fd33b04b4f53ff41783be06ddeeac966c9c7bb4b4f7dcfd20ada8bdb9234ffe9967a9082bd392033afd3521e23bbab8c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4642d90cf05d84dc0df25c40ee01da163e3b227ac743ab4ddc76deda6989d68ef694f401d205699d179cc207db188cb6413;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb98a25a575a2056694421a3b8881477151105243abecf21169d251bb94c75d02437b6c41b02e3400f46f950bb93f3645960b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'habc680dbb3c08d30e87a0a98520e5d12307a8b49c7f2fb9e1a41c6085e5f3f26e4154e241422293718f49948eeb034411906;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc38e9de2366c6345245530aff55bd09da01e4ace933ceeba0dd85da16b4d4c03c2d4735db8658e9755d21338a72c7a3f319a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h517d639fd0860f1638621f1a4d72badf1d5c89ab165760fc9b2c628c2a97a38482956ef6e8176add54ffa579ff18c9e2e084;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc20bcf6efce489cc243b4e1d989d0ba0cf9a275db7c55e8de93e9a91271d8f23819c9178e8017c482a7685477b7999240760;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he47acea4c220f19dbba7ba3da1eb48aef6229c89d2b54219792bb3e245f505941bc7f27331b11e683cbb3b13aa1a231774d6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf50f8d77a87f5339b72d6b198256f507c08f5162584bbeb82eaffe300bee03f08ca69ca2c28aec42d19fb10ebcd1d716bd5e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h662c821269855cf151e8508a29b07cc616cc7ee546c318450a0a6daaa65c0f77237c2ace261215e09897d9b9c461c33eeea4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h426c5b94b0007ce88a61b55121031b5ee719a7f2d2650f7cc59ffbb5e9df04329545c1a98eb774748d794a33a393a22c4c1e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a1855f0791d583f2a7a91c6a3e2970f414a1a2e4a8f38de0c064bfa1f6a9a790164dd8363c83a32e24f56a968a0a75c2edd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba316607fa687775d2418abed6636784f2162509d8c05cf0f925a6df68ba00cef816f93463d3be85777924634c98731f71f3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82009a17c879f099e6d95712b7cae4b1c185ed35ac44825cb4f4d5a8ab9227141e9b5019ca99a6320110ad8a8d5172f3210;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe8ec1e1b4d8925d6c2a245038a70ba0968fb01c3550749b3d419add6bab55e0718363f1f02eb3b394b331cd20857d3df4bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9908fe880520b28fcd8a0fb8cd165fd2c7ebaadf2439f600f9a2ef9c88e85e2024cf4e0b70e058e442f2f9063f378a4c52bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab338f1285c41f533ad455d249fdb2d6de75fd53e72128d56d4e4ad407cfec2f5b62f5989e50270a526012d73dd85898a9c7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb95b45e64a67187d09b479b7e50128951132b98f78acbd6bf2e6e844d34119feb54e3c44013bbbcc7a9dc5ee808cf40e357;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha000bdf2845fb5fb757966b3d30f802dfd000f5b2d499c45ccd952ea4f94469500cc2316af844c9e18b4517e57ada985cdeb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78a1356fa6bc06cb4fc6cc5371cd3c188ce76f4be76a29dca397556da31021cffb3168a8de49368ccb0e7cadfbe46a6a5faf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7404b4ea25c3e4d24e9002efc44412bfb566b0dff4271a9d5d448a9e8da4994a0c10b881053462a5ccf15d0dbd932962a371;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d647a03fe3aa7af9f0cb05d3b8c45ca9947f92f5e6d2c1d6590eaf99fe6637390edc46119a0d0d42eb725005b9d26b1fe69;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1d037af437c49c41095aa194995be435759082fcb4b666cac277e3ef6b9e92de3aa323642e37d92f33b9d7c44589cd1e8c6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ac8e6bef8854b6f04b22b7c5a60b4a64867d078900ec67c0bd0e9f0caba2cd978c3de880485a7e02526261a4039074472d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41b484b19bc5cbf327e725f384a08d5120e4d8afc565bbd616dd641dd2eaece49392d99ec6996b146656e508adcd4b60605c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61ae93414472045908a0f6f52c4bc77db21671d500c391dd560b581a2e580c1d21605b7d99cbf8dea9308161c96d200194d2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa865d3f7da4f4b1314e74492268916644dc8fcb0faf7e09c88b4ef2b0ba544877596d74255361940d3fe0dd9acdda31032a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0f3c58014074a8c8492f37ef000b06ca8200a04ea22c3a9363a9314423fd94c554446aa9e0de97bf099cab5c7533c16e7bf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd97fa7d1ca2969aa70ef11518d584778fc8a2fefd96fb20349b4e49733de4d0b92e7f25d23f9cdd4c4dcfce26ffee9a2347a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h698f6a0827754235ebf297eb8eb4bda9af525fa20582e5eb34adcaa9c932c4562dd14def4b9273c99d4442124893e02a9f2d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haca58667a043522ff6125c9ed9b490743e2c5e668271600753096e62473d72fdf65367a8ee86306c2f2d2ee2a988d5b986b5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d4d54b80742472da8b981fcbd0bb424ea1321e218863b22c9251c8894d83c41ce3dc7fc387c7b4b12e2ea2d68aeb1475aa9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1de061ca40b25d9558a68b338e8625dab58cdb560ccb1bfaacf8d10a121602de08ac5b364d6560994ac993c1c8c8fd5a0399;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a2a3b77557259559ca6161c54f40be80ed951acbaafb122335b72a24a51233837eba44f9ce4ecf075f809bf1d72f526854;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h975306efcea8822a12ccac3f88eeafeaa775582a3c842f4818d364e9e1f7526e21b7d7114cc9ffff564e779a869d93a989d0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3fdde8aecff58719e00986deb285ee974617e29e335cf7bbc8b34c49c7a8869756d63f3fd88a407767b55a7fbd28a1d35420;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h712190af55ce76f0630a14b9ecaeac7870a7eab8200164461bd3fbaeb7adcd9faa49e1bbbb23b585b8ec6f7f6e0ef1cf1c79;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f26a6e4c8b2a1ca1a55517170c5e35875287dbbd97b243d790a6070f4b700ee7a74cdcd362bfe3429504632d474a972e0c9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5983d5c99fa4aee16c80e8a23a232e45fdee6be42a00aabb84364f558c437f21c793af67d45c7b905d25f11d33374a296a82;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa1b6c06d6464216575cc7aee7a1e96acf3268f3ffd5ddf8b5d3c042803384c54c70358f3e0a9c19a33f68ca042f06f34e96;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h783229379ce5cbe35785bfcba69e948ad972cf329d13613e1d37127a2fb4fc99f35b27eb9abf761e645561ce96b115075931;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf102a758f875b6242191c75c5818cccd8cd6ec4ad95504836c2c3bbf113f515c943a1ceb8d83f9280d30740499c9598dc8ae;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec82ede3b29a04619d911d461e113f3437a0d1390ce1e9c59d0550e2a7af0527ecce48c419b12d10efae3f08793ce7f76e3a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14ff3a5f42ddcad0236622a1411c4be4db8a55b759740af519ee050dbea22ad39f8ba38500ded22a718875efd1c4dd0ea3df;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89c73b333ee081387f28c4185537fb23b9b6b0f5e4adaf54d4c041363bff33d0ce4b889f5b745379eabad3d81307ee015122;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e0014fcffd2529b7903d287a50a82974799d46db3f507b6e3e128c0752dd0a61f25e75190edf9e1807e3dd9c3c5860deec5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37be1b8f968a080d6097177a9af34a8bad47a6107fb038b9168ac966c667404cb4490cf490e0c40883112c40664856403c3e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7beb7e95c261261e36a3a8f0934bac66678b1012a6309dc1b0b78f1f707f12524534bc030d3862458bf2f1bbfbf897d7377;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5352343fb7dd32ed65592091dc8ae33c82a35138c516978a659a44ba1afefcc019f43b37d1345b971b7fce87a2593af326a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h495c55f0832059ab4f9b0c3b667c58222249f1e0e195dae556663734bfce42b5bdf40f2cc5d0923c9a0e1c07c46e47ed0f5b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2fdebfd9afc6ad3ba13a4ea9d47b5faad825a88fd99e7cc37dc4dd5f7b4533cb23df108e96eb4ba4a742437a894ac2f7dc5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c8bc1bd090f6fa00df74e961963443ea6526df453a93b9cc19f6e8aeaaa1992465331d2cf6a9b10c3f9aee6b20aef9fee4c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52cf194008728ee23c395b92d4fdb85c651d8277260a3b0c0e493494aff92b53a84b01467eaf336e2009056ac748080de76f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha02429d09dec2fa8469c501b2a418e3a70e322a5369497bd0a0a679b321e98287c559063ce9a3dfbc559e45621cbda4ceebf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a43aca64fba0a482e566d97a93942380dce985e68aa1076f144773940fd57299ff0afaa00a2f1028b05726e7f7f3ffec4f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h282a6a20ba3f0d5675c27fd97307cbc04bd5852fa6494075cfee4217a2803ad9a123d62c20dbb1871471fd95e69450f24267;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3149888344cf6618b5c8c6fa3478c6b57fac859b482b7234ef952a635cb9c7f5177a0aaf80dc9af1318b60993db296882ac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hada0e9bbc5e2f0e3d19ae86b414550e00b81321ce60d4c0f4af66fc508069cbf72a56a9b97c06675859404a0d8eff7add1b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc7b13a047e94e4ac46e2da947c7d9dc18cb0fe4c41d7eed8f359b1f18b6f23d2dcb28689b1621f15d0c541775f983acf771a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd8b6316eb9ba1e0867e1ed409b82e0ba55b40d1daf21b23426b5540cbbaec8c3d903d43d0a0bf1928a414af1b4d3fb61dd35;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he73eb1c1ef36aab4cab7df9391fc88b1281eea0fab5814bf0b3f87554ee73be5231ba40079f2a2a93dd30cb2493b1207f62b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1e043b02c43f7c6861c8eeb0eaa58a548ce825459d703ec09095a3b688369f2710e2904d91492549b77fdff794526c612ab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7df3a251f9cbf0fad6c871fa5e2ab10742f6535e873da864cffbcb5b6b1e97c5fbc6c5baca0d95edcb013e3103328661042;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34babd8d1cea11d29de4ad485980b90b327f30c4b67adcabe1730a0e0f721bdffb552d3da6a6d49de134922115c4018d25c9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0d2daa5fb536b4d5c8673cce0473e8de614ca1e2eaa0ffa7d38e41ac41755520641c4345ed6e770f510f972f3c905b49822;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd079ef5a6c551c965454627e9af9f80eaa8d4aaaa4536b9a4b2259cf35347fe1f67e06f6ce0f049c486791bb15b394dc048e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h43cfc1bcdfc5fc06d1ca428ef72ce9fd9be4f6ac68592d0a3fdf461dbf1c24225b49f5fdcb9136ae1239e661cd1f759bb760;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69163415a13ea8f0bdd3254e08fa7dbd5dcf3aa810e9d38a382eb8a14616f267a563b6126db296f3b7fea21159603d8cb146;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb4492cfb72a87c14a63bf6bc170cdc011d6727f46355da3a54c82f301db50ce6b024e9219820f5d6dc3b2172d9a32193990b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h480afa438cec0db9b5afc2e5cfa683f8b2a149fc9500fa179d4aef38dffd71efab686872d880c09eafbc683656f27af1e464;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf5c640f98540b04bff7ee7fc3a20ef08169ec3f6cdceeb851d39599417a8ffe16632c39fa64f34184dfae2d3a7fd67fc7a6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6ea226a2de1479ba7d0e006d6457f252368a012dc5fa3c1248bb0504a628fab03b5bdac67849530c0c9f27cdbfe2954c35e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13e14669581614607038308b0f3f70b2c24fad309a1323bb81323a63bd781b7254be8a2fac975bf77ab835926340e8153137;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fd77db7bd15763aef45e360835058131d088cffae62aaae2ab03adaadf68d22fbbd28d7e3c17c3f975676196e106483ba63;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe955960740abcbf7836dce1b6edfd159c94a8d7036ec5a9e80383ec88197fbe75f5f5e56879d1a1deac9b854c26fdfac305;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heea8c891e4efa232ac52378c5578039b9670dfadd725323e7ecc4e1f6b46d31d43ecb67311e74c3d744c1b5305eda96f7c48;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bf39ee236960b2ebafa68f0c23e5cf4408f0bc5d61367ef4ba1bea20ac96dc4d36341eeaeda9fe62b3d2139d8ce0474e7ea;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h350c6f2909f0aacc524c4e9a8768295bd18090368fb3fc7445aba7b6057a74042c6a3530f436d9ff6dbe085140fa0065a529;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha382e37dd6ddd0fd2916e4e8e62bed956db9f2cfe10018c55be60525bba7ad95216d3c1cfe2116f5f64b041724cb5e3eaaab;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe8059d22e2d968b34e81876ad7712782ce27500802de390c1dd4deebac74311d35cf33816c4d9ac3040a78e02c3acbf3241;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h311ba1102ff68887c0a063c454a82bcb3dff2cca8fa9ca2497a3ffc7d75cd482fe0492a1cedd07efb06628851ccc803ca0bf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he46814ababcf4b413c09bf6bc68d19621c248454a3e779432067695eb2ad473784f4d47f2b8e4a01144820b518132e82f9c2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77fa9078dbd861dac2bf1f7e37a97432e29b069dd85d78f40434fbe56096ffcc83e35bfe1e2522c5fa45078dd7754e3b11f1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6e8c9f0eab0d9ed2148e6aad1438f0f2bcf25f85465df85b19cea57873ab97412e361112d0bf530b7aa40dd0d6e984ebd652;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd9d0a64378639d7fc796bd08a413bf6b9a5e45889e561c2e637fee68b5031193e22086974db8b512eb9ae642da4eb7c4cc7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c351fb31922f8063eb1adf24c00cece37ce9be49af7c509ebfd471a5dea2243a4d896b3a3c656acd3719cf1962ea8bf0b43;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba887bd4f3207850ef1f7de7af1187381313c51750786f891420803d98a6999709667a8fafa43d7407a969220c5450e6832c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b48101f3a2e370f36af69603a1d567f345cd382db9106b9ecbf237531cdd3fff0576786e0d69992a59e346bebbe3ef0e1a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0fdb921803a91425660eb5b4136c4017736d3b20c7aa096be060b79fad4ebeb1328d36af809cac67476704908e4a2f89d88;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda59cb559e392cc9bb203004c08d7b6624f5eed641d03c7cc57dcdf012a2b6b8617e71870e76ccd31357b9efc06951a776ed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31fb4987cb0dd8e93bc3e8b07cba24ddb8065484187b9b0b5f62da229836191a6b78c4de8db6d75f513a4d8b071a3febe1bd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf52c965485c90c2b5e72034518b97d3d1dc71ed263aacab49ff9bf02b24f9bf647da8cc9c5fedfeee629c3bad378efb23f9a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he447a3a6e10ca01e1eddd95f0169e9b1f452411bb5233dded59b045ec83ebfc9f8a90b1cc38ba681799099b48993ca56bab9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b5420694744c1c78372065c74896a9460159ea5b0bf67c29e3e8d1f6a7d9608dc3c41e1e9a5e4d287eb1138d4d018480712;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf106191665cb5e8e461ab70a943b2026ff7ebbbc3aa26e2c5815b7f06960fc600608b0e61d8af14ad9e569f518ba34ee470;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb87e4c8b7c4e1d9bead22e2875805bce8e977942e6f6de40d32a918b8a9b8a85c385c8e386d48b93b6d46808597f2f5c911;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc03405fcb557119ce089ada78e1fabf384b6c25435aca3a7fb785d7705b1684a143cef086a795d1afbc8d48de506b6e727a6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd78ca9e3e1d192d57c394130a4761912b9c428da49d04ee67396784daa230ecff0e987b9bb9d371386e26f1be0d889ce9775;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d98bda36c4742c3f31420b0838c38f2e33f568a32e011c85071615e38ef4a8fe741f6e471ff37bfc8f0c5ef710ecb522408;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c8fb6fcd4d0b95f8370abcdfdf1a9da8f192cc0b3555b8643e2b07d86de7614ec758235a3631bed987faece1de4c83cd061;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50292e7172d749c4010e14197622ba78725f79cdd18de4a45f9dc3e9e29705386dc0c728d90b5a2520b26ba19c017220be51;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6072e66550562138ad135fb9668dac69afa9324f34179313b9f05078a0fcf41eedd12084e808ed7ea84a7118824681590a06;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h225c00b11ba306fe47c6f9dcf44a08070b37dc88ceab21499893bc57d959acbd54ab095014a9de94f599a541a0d97c2889b0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb227e8aa96ffef920b3d7fd83321fae5368ac5e18b0684dcfbdcc8587be79118cffb8f8e2f72f7092e83db1289c0ba33115;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfef0e23d564158670e3ef4127620fd325a866f404dda1102561e84e971afce2d13ced3a561b5e2084d3f472ebc1ce57238af;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87916b71aee4718edd4fd0530d13c853d32727b7b4bb754985863bd461934af9cb3f9ca3a67856d78b11d08cd44d48d59578;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6390ec26ac36c193ac1326152bb5b406590ccc13ebeae40c549c50259c1d768a8f3dd4d27c4336f1b312a8b988059db1525;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96c18afd540a60f3934bf1ff878738231463720be1799201d0683a1427e969bb6517058d589f9ee468d6d6c61c9b94050b6e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h396297dd39706b8ef2c2a037315233d6d3f17d2df46bc2b8f851bdd91d3dc709811cc7b91e60cc61325e63625103bcabed5e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he33eb7d7262e46c9fde82d904e5939c18b0c08bc16ccc642dc39fa3989a0a3cda0e4b71d2f43dfa666775b756d2716ce5dd7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h382369d7042cf8572dd46be5df77d35792bd78614214bedf1c9e43da6145f39052f667da34e38156893ec8fefd6fefe7adc2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa88c2449f6e48ca8ebb0ee603fb483a46908319ceb3201a6ff1d382618aad210945eff9340e4cc3876228bfbf7fde510;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb394f826af4bdec23eae38261d073ca60cce90431254bd2c3f47016f8afb3cf2424eb19ff3363fd349ac4f6ed365971f5a33;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8b878e74cff595c1407741ad2fba8e63967141246c1fd56f4e40305a23f39556b4c9f1674d5857eb87a5471b5b9816514d45;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2bbbb32c48a4bd02d8cd4b67776fdd698a61dac1b2cc740a37efbf863a4466fb6ad9aebfcdbed2ebdc4b20a6a2122806138;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc18724200a1bfbe38cd045821a24c2af2673fb4d513f1fb18eb34efd679752586d7e39f4f43467b679308367572c692402e0;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b522dddf5808242882967de1ed680a03002c278757fd38c65f013b0bd14c21141800e04418d437d0be2f840c51323fd8a20;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h91c09b16f71dfcd4b21f5830e2ddd4d69e76871f5976c61a6188d3ee704b7f59643b68235af26134ea1b7a228747b0e3341;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde253e4daa2969c85a0b0e3c396176eebb4bcac708b5fe3206957117379cd640d8cd363daaf4432e9a8d8e9419b20bee2b78;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd49eb65a5cb720c92e270f45601457006387c94eb57819ca5096d1f59b2ed60f97dc7f9add2f9219aabab3d51e441efa703a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67861e1c493e28bb2109759a1733f7b9aaf050355d81edee3c642945fb829da39166283c2bdf646c5d939cdd09da56d6957d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4ec979bb2baf3b7032d538b53f286da051f0a4a136427c45f5e15bba6ab10568e5a5605e1f41e941663f45601575285957e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65dab8c81570aa7ddfa5fe1b1a5c8d86fa0c5e48723f981ab06f57dac487cb28d9cc9dd63546002a5be520eae828998eb1b1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ab94dea4a25c0e5473180209073672fe10c571678115b44cf72af7973db7e480fe4e88e90c6abf68394fdc59aadfb61402c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1436de2a8bea19bd66abe343b6e6d3a3a4a78361690d901a7399d8b570cad1ef0e4b432738768aafd1992407cc46377ccaac;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h90e8579330030a1c6ea884b2e690ab2881ffa14884e63d30db69d79228cc0bd0c36cb83f5874d2c4f0e7fbdf42c3f0dafd53;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46608a8611d123aec492ec4ce5cbdaaafc73678f8dd6031c4b71cd8ffdba4aac8597e2c6ede915a0ac98107a17c728ca095b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11463db34f9c9d31d6d4c372135c377b55943985217cbc5f87cfbeaa119616344200dd8374141dd0a6e18f3c886806bdcb98;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f08cd65302e09610c4d996135fca1111ab74fbd94f3341355e2bb971b7eb5dc04fc66628ca0326b2d34ca92ea817f5f5a59;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f2d6781196bd4b2b6e8a0bc157083390e9b0487963f1454730d85a694d0f8aa8bb364682529680e5020cd0367914c1415d8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfea81ef1d1b2b1c3b3e8a0245b838ed5326b09d8b0ac7cc528b96801125814573f9a1b8a2153aae2593edf453ab6d5217975;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff2fea70f4c6e41e57fdac55fb036ce865fddc36be38aca984c468b9e78949d265d763bd6e96757b6a229a1298613ae77ba4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1056dd71fc161b23ee9b95a81ecfe94749b4ec2747425025ddb93d52279f6c2ae26567d98ab6b376ff6517b5125ff27d44de;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4963d6f017ad45f6dc689e8c33710dde54894b53dd1d8402f6a954ea7b2f78c5cb775c1fe3f22938e4cfb3858cafe1e8db95;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf631e4a4ad12ea1e6981ae75faa9f23f971581cbc51dbfdd7dea409b5288fc727706a84b0e7cb1238d3189b0816baf739b4;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf202e05d4dcb60421e8f7179f12a8dd3ee434d35d4bf11703977d9e5ae827305a3e5973473d5cdb67ed6e75567cc26b20f47;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb7f0d0d6c95f56e7dbcc0dc70133d2ffdaf5a6064c3b92a7aec28a8c5a204e4046f2e7fd6c261d0882ded0bd1230e006f0d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf17e4f9eb94174210a97818ab10dfc9e9ce4bda20affba2a1e4b7287546c8265b087eb68306275f494b38cc797e2a48a8b63;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdea1a13ec1b68228d534178505ddf19fa9f0f9343ab782f98a80079e85353fe9417ce2070bc3b66060fdce8b51299fbcaad;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h657b71e3c87e826f9f879cd98c17e6c403317ce036bf78160576688499d4c8656f5849fcf9a3afafe94aa6b3812e545e5bd2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4badd3347c484314aea9a89488adcedd8efcea8c34448480ea3479cde6b1a1d260a051b7258d37a4f025542d0c8b19667d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf919b37f0606550defc0c7429ebf643c112843dc51c1e01d115fe17d163d1bc7a64be73f5b69b9c8506c092941d512b3e0be;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3b5b0ddfd93414a87b856fd1968524cc97dccca05d366596383de86a35e41705411275bec40f1d83fd14311af02a35f2899;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f1fb11a892e0444fb0ddce8c84b1cc9ca12990bf717b6ac0dc45168bc4d63b0897e662a0cc559ac3bad66b38f3df5dac88;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7970acef449d5e2be58f54e92076f9d840e9983d6de00a38aaba383554a466fabdde1bd85fafc7d72f00c00f819ae4267e15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc175b5b2ee14a0b96ae05ea322822bef557b3d500a5ce09f05abbf645baf0a88d4966d42eb72f6f80306ca7f6ff2fe4ec428;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56360bc8f463879273fb242f0172656611c135b088ec140563d4a4ad963cdd184683319f5b6582bba6ac13be572f103a42c6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4375e7fd89018e6292fac74a76844395802c94e7ccff0b805399460df4cd41bdf669413fb687580e5fd62495581689e87b4f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha909f9be6b9df0e17ac84aa5263748fc72b69ac1da2e95d7098abb74f2ae9138b0b10c758771e67c58a4ccbf9d26c142b2cb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd1798e9c04237fbc77153c7dc9fea047f9c364e392c4bdaa5ceb0c11d2b669bfa76a2799c8078062efc6f8c01d14c935cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h135d164fe6df324befde2916c8aa855fa94859851cfb719204720825ce8f352774cbf3f33012b4801e490287ad3e4c6fb853;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h847b1c6b2a819cf19cda97931cd95dbb54366a14790192eb40b2908875840ff6b4317124c6304a7b456c19290955bc0f6b7c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6860e4ac0bd5133cfabe727f35ec449d5336de9ff716d1290a5231ef2d837f29c599f8451a86c51772736beb3081ea5d9ed7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c359c784159aefccc542a3aada2f78b5ee5f7353ba0428b46c0d48168fa9e1831261728252e4c5d36d0f7fe860a27352e96;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haea718e2e9734034ca6811e3d5367023792d0c85435abcbbfba18377057183efc096d5685fd38fa1c97ea4e1ad2b1b5fdc34;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b48f3b1a4ed47d95308054804dc389d6153e9f62aca2e172b2db306cb94cbe1cee7c3f3b15c53d755564d6d167d9d24107e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c3c633ffbc081558a647892dde0b960164d9277a14f99c15e8460149bbed51b67416fb977cdd4c8998ea7a9ae30b9c8b490;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb7deb03306ce230a37b6db44279863e3d0f607fbee0955ffd460e6217baf6447e9da14a816eef7cd738ad7aec3f1218e0ab9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d6e658ccaca4689406fe9c733697ff9c54c8e415f6d40f6ddb8987499474931f84bbedc96e9fda969edb08747540205524e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa44aa65bc190dcb58e01a4e3f2a4fd6776df3c1b61ec6793f40a8c9a47ae524064922a0fc2a892878f56c122b52d601c07e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5646126c98bf25aaf9eaaeb76faf042723ddc39881a22826ddea8ed8a5b59a3e1bbafba371a69b96fb3d6d727545b36198f1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f51102da7b2610472325855f8fed9f6f7847e71a548830950927d856f8baacb7823fcfcd9883b62dbbe6dabb95527a7d2b8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62c739e4f904534d29a4590b3dbb0cb74e9817b9bbdbde9bc0237bc503a7a0f85e56cf9bac79793fd5f99a50a13132f6968d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3dcaebe823500fb619f5605d7513e215e4a214933280c3e34de2331e7e534d036302eebe9805a9497e2e265e720c17f7bd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcab6ec2e8cdd65c1a213626654664c992837ee93bfcc6042f4dc72501318ccbe8fa8fae3f5c087f91b77df46ef874a671ca1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h931cd27989dfb5c1fccdaa73afad9f4551c438a0364effb02d3651ad1afbe1e5e589be5b6b86813ecb1ef07ccb91db31b60b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d7d8d804c3aea8982e4ed3bb05efdb268b47c080265e7661ad097749698a986be1647ef0e72267cc51584f08fbc552c764c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7457135ae5ea670e08fedcf870ec335487d2f74c3073ce18d5f828626fa5eb93f932732b6c887d50b3ae4a140db2e0948e15;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h671d13887135f67e8d98d81d59570fdaceaf42ec1e4da78b4173754fecfe0d8c9ec1d2a1bdb00d74fd259f12f996cac3a9ee;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d3c95c8b0d0404f28bb267f51bb3c1d8caf28f9d090f37a5dd5da729a0861eec966afb3db3630c8d16b9e9f03305895229d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hecfc20dfcee0fca4b6ebb16662d784d1f402c4e72a8d3b38ef347a6aa464be9de73bfc81a114847f3891b5bf5cd5f1bcaf8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e1667f9232004d8b60d71961e3d74c3d88f737ea951ead2098e3027f30603ad04efd78d48ed7f673a3430ddcee709855a0c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c2c0889d39e1ffb0af7457f24aac201373b1a8fa53db3a121719d0d936229f45d9e61f629c62107b3401c294330a6940512;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70eae5e61db1c60824c1f3ecd3d45435ba22d488f3d19b3c6fb364a08ec113a76d8d4bd8234eafb1a915c6c915b7f126915e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heb9cb5c3c3c52d75e7c20bd4265e126f840e4222dce140a1f045433c1d931f115433c99d6081a52fa99edb6d1cb5d19d269;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e77197acae115712aca0fa2ef55188dc99edada16722d1d6da56483434d1383fc715e580ef33d9adb9c77898535c2c50b56;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52999e74706aa80d5eff652e7e62a77a8c632b95cbf528bf94ac7994066a884e0a5ee812b7ef94efe7c085ada207b7cf5c88;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a6f3e3497fc3870fefdf4b06c845667cb525d3c6343ded255c5e88fbf5bea68b8231495077dbc5385cfcb48702283b8c02;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdf52a077e7aae507393f4a555ead15e664e7ac8d89e4710c9a1129052141921af686e7ce719b2cea46ed7a6bf31bb61fafb7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f787fb67a00020e76c082267b094e554cf5a9bf9f8ec1e1278325110c01d1f0390705fbe44f09c3e46814c30a07e08fdc3b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1cebcc1bd5619c321b9f05415f66cc6aa35e214ddd2d237c00ddbf213760df8e478a2480f3b21427670a8177ea41e432c67;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h248202cc6deff150ace2cc7a8ca323cbad3cb9fba41f2fcb2919fb8a8ba136ed1b44081199e94d8a6446293f35b24efe13d9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32dceb0f77e16722cdf45fd6406795db8d0a7309280f7114e9ce9b683bca179ac3ca0779e01890eb614479c1845dda9d91ef;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f1290dab0c7edd8643f282b984385f3f37d6d8166d86908ec3da0b2439a701930ed90bfd07405d89a9aadadf1a1d048cbbd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf26ea356bca4b082e2dfe0b58021725ba7bf0c24e83aa67965c79275797430d1eb1303e01da70c4978d7f7072397c517761f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd89291af476f4663732c6b25b0f35c5dfb1088584aa709248e288a2ddfe7bae63b467e4ea12ab690ddc0cc7ccf9f0fa45502;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e17ec1889e7e1d98c3cba960bcfa06e4a770645bac9577b1da6131423740cd34f484fcd9772a2ecc55261940f5c600b9d87;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7339d2541132eab4aef308e9ab69fb14d5f2a558ee351b9d4180c97807ec285c606065e0077bdaf76b71618fe94347dc4c4b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c19090145c463574bace7ff70905a74a91b57b18005a80fb61ffc3b3c313a06a745e54f9bf0fc26bd4ff4020beac0cc794e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8dc0777049471d651db358cb81aae15c9f99bf22f04c4f051d59660234b3b94f3c605b62e571f3018ab17eee4aabab3aebc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9596821b2a90df17b127bc05aa522161d5680e7ab0530f7ed0ab5b009c5c02371d6f6fd12272a13893c4a4e71d801c5abc3e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb964f07dcc11cb9f189f6b3af4ca81a7a6c99a097d585dc8512f884c41c6befbb770b8fb413426a310d2b31bbd0df1df980e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd809d9dd1ffd5b579b81624bff49879075bb0af3e12081f64d6aeae83c36abfb9916bac5d78048ab01373bc26131b0c9ff17;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8a55b08f5ebadd614e50a3161b390702254901883e1d644de29709476c53c75d9c2f2c4f5ecda1d5b546b40e20680bc826f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he162c8f85b79377b7ca7ba9a22354138ea17401ca29223b520c4c16d3daabf01e92dd14206669bc952f33a7046c5615db8b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h985aa46e64ebd22a3ec00a9f093a47038148d2d85d3b19d3be35cc66996401da6b2da4b2d3c5f61df5d5cf4602f77434aaed;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4560b8c15d32685b0ae0c2dc5d4b0d4cb211fd9546ac3083b3cb9eb73ea8d45b62b2d60423c27ebf1c80b2b3cc245f3918a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hefcd5e49a960f63db334c46470ccdc44a0c8c242d1fa99a29905866329e56060f845ea07f36584b3d4353550a052f952ef2e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hda277a94752fa1a32d80cf6ac1910783e2b715ef8bac069337ec8f1f53823f1e00fb57c4600f4c99501e2e0a2377970fdc19;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h649bf30b163a2c3f3e4d09b01c9d29127801bf97f5e9d1c3262534a58c9974c16353eb89596d3ddd43470661738cd7917e88;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3d8a6cccd23e42ea4ea632cec3f51a9ea085416a74e8e201bfb2b9d14e83d3a9ea3d2a79c0d621f59a5c8d9e09ce64fc1cf3;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h63bf7dba6f9a7384b2588384db21494e505d0b5c23ed5ac84a5c527b2d3107968eb5124de099f74dd576ae2371a8280bc183;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4435daffed94ee2db6d2760ff6a8b8998b81c6cd9f562fbe53f7aa55b8d7f0985e1ecc21aba948ae18428974c461feb483b9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7adbdbf07b7cf8c2445b677dc08e904b9f0263dfdddb1622c8e0e4b1ebddab8b769ad61ad3708338a4b861d721761b6555fb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55a4fe1d3d839c8aeeef9ee0ae716d4a045f850c5baf45da6894ac902dd027f7ef54a4ccfc74204052618a2454efd9de0af8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h191a9b20c50fe67f799f5a1b2762ea3f41b9542f82c2273ced5d025db9a880c8a6cd2d28783a502fc4cbbcc887961ac0bd8b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2563d068d2974d862e4a9d95226f52ed93a70f944947319ef5fd4652c422076b3ef8be3fe928067bc4351e7d36905c1eecb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9867673546149494062dd73ab283f32d7c97634d039048b02794bcfdcd66b54d85198c35a40360f0d51d4be17dff2d7ea6ba;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f824833659cf1bbfa9eeec8ef25e5015fbf3e402a7d13e1ea2cad5203b4f88077fd109d3436ae4c3fef9350008d174bdd6b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbef1cb219ba940c43dcd4a3a0240fa0386faa2042acdc00f453e44e60a2766f86bf2133da84143796a90e58a9a57ebd32866;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9c653b204f7533e8b5bb52b22d3efabc59df3722bfd4537f08b0b1ef23b1b6c08ad3b15bca738f1cfdabf5a64ce1503951;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f14be1665d7791c73b4506764ad1aaedf1672186de0b6962525740aa6a5d2ec72e664e96b4f88c5008bc2e08c455bac62bb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcbeb231df6443ebe6773502b51077708baae0bd5acce4527d58a513572a7c23a6639a92390e0b448af05297ffc51dbd56b95;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85d2a66aadc1ef98416e110750cdbb0baa79292334cd53c50ab6a53419b94c0711423030ee22f8b1875ba2d9a95df54d4410;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h489521de569d3dc3a8833e2cef512e41a934dcda5534e43416f83a79969708582254eae75280933be8969015028f2d5f161b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd63ba62b939705db3f70a6782ac499c18dca7b18d1fa03f3c38f9d6b4fe381aee5c148202c3f2bb8d5daf8cb7e90907a978a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7aff50ba6895b67819dd52ab082cce10ba19db69ccc7529e8e9a8867afb723a42132470a2d49682ccfc879fca1f1546bdb74;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31ca547f29d39232eda08242fe262af77735bc4a5abe95486e4360f5d9ab687e75a5b4892080a0a47f8a1f51b3ec31eaafc9;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc5298fcdddb71328c078dcc4bedf72ba56c57c6a51ed7abb08070961baa23add2d2944b79622056811c73757d3e38ddd4e78;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc2a5d911f047787cd5781b542e52a866f2265fb3f95e7944ceab811f5eff764e9f2f9d628215389fda1f587b4aec87d4da7d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70822fb1a26e12df64b03fe4ab85d3d8160251ce28986793b9f8bbe80706db2f10aece091b1fcfefdebd9bc4b4c915d36311;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e6adcd16c2a237299a01048e6776846e5dfb83b0401830f8f271e9652db1908d73c6708457676e846434a32e9dc5622fb5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he769c9167604db9b394b75fdb3f0b3c0624acd05ec2869eb44dab1b708e2e29f92b7d19ad45ee81dc23c5522bad19f73f199;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9720168327ec8b7c25c74b4fb4134fbcc860cfcd07b282a9e12b60f160da32b3b767edd133185d38f8ad34430f99bec1edd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8cfc01c23ff535a498df520898592d5549349cc6fc8077176063161af0b0ebad098072ae4ff87b15570f62e04813aefa96f8;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd88bfa2201a57b0a3d6b82fed4a1e5caa1272d408455204a6e80c1ce75f1ac04398545f9ad41e0cdf0f17f2456d79ce0736a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41c4dbef13f098889a9dffaba337beebfb56e886c5e52fb6536d00742e8a7c8791e77eb4fc51260a945f0b2569b64fc63757;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba2a2d3c325e8934e89941133c78931f9fa41e4fc04f5f99d41e4df44776cfd38a9854d5d7b132e46d998c491ba4eebf161b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha36208c581ea899703705c314228c414b81e4c028b3a40cf0aa817d99d5bdf537565212b461040ebaf257269fa5fc58d2f3b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27c33e91267765c667a3ea5964c0f9fac8c9cee4e6c40e6df9a3e13e9d066b03436757899f03238ce37d698464b4d2631223;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd049525bef764b9e0f6914e407ee81a68e0c476bf45f9d91b20ab4a2b18ba097aceffeb19ad786135a7de4ed379cff4a9c97;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h338a340263b23a315247b3e5a571ad453784877e215210cabf1bd72241237491afa64d08fa258c0c5dc8e6730e6b9f0a6e7f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae034c496bafd8f4bd09313696cce1b5d585542d9a133b7d16d78ca3cc88bb20710aa91a4a900aa3d81a04348bea6a992209;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ae834b6ca22e7804be663b15dacf525f2a8480eac06cb91c07b00f37011ed8c51405f958eb6aee2f4fc58c00bea3cbc4a32;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1aa2e8ca39f8c5f852f4755f43239ab625f430853bea0ee05ee5d2db33541b523da801b967e36345d60ac081adc330ca0a5b;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h879760b84378fed1b105d88de75f8458d6ef418d50b3e5d199db7fa59a0a22dc8da549e90b311be1a5d20a0e9fc67e6d5af2;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5769a864fbfe8a8c5921661d7e22f6b2862cd3256f370e533e0eda7446165b3b8ec216974b1e7084362282e91984275bc3a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a15b1d5bd919a21480b54cb6bad06f5e85a921a8808062299f3e9e27b6a3fbf65df46d0c0f1cab1be78f8875f6e0a56b140;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3b7aea25f28dc2851ae91acc6b30ca74c66840627a905adc3dfaab302d30261f67b866fd63314d9d7314e83643078b65ab22;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f50ca67275e3d645e1c4199e30d0e71b4f3c5cd10d5e4a7b58cd34167d4189a3d8bed1acfd46cc22f30da5dc54a02bef0d7;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97f106dbc7aeb09f7312a695bf8686c515942f8f6ff817e644704daae8bc84a83394fe017e64cab4a03cba40433adc175ebf;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa31852bb6f52852a33fae5c161c375b4e1bc2934cfde9e9600cd49931412cf09b710686666ac62613e1b7defe73da05c78f;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7433b071297f5000b98e21eec95d1d114157b71b760fb919a9779c86c221c511cc6a38112ce24587077635218de75f933c07;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd65bb01a79f29f2618d0d2ae9d2d8eb10fce0c0134bec834114bbace36c3cdf75bb9242277c5e936d32c3cc141c674d95973;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1ba9077f1972fb1061d71eebee9c030175a9d9225cc26ced06717b51f021782705aba42352963881d4984b17365bff3f8d5;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c76c0049835bb5d0655a2d6527290a8f86e585a4ee4eb23c6ffbd6401ee5d8a153b42a4a531ceff77fd5c2dd6f25584a21d;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31fe9aed99623031db5a61443d2e1615d5e3bbe319489f7978f2e5f487940a8588a21cee90d88fe23b856d06892e3320abdc;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab0e0bc4eed642d880a56db31c5fd987f28770f0079b6340d1183a238a5f909a644ab819bcb2fd105e37a9b1fb2e296769eb;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd49df57d541f1e971152e86010fc1b0428e5834bfca9b8cf3126aa79ae70e22e11177dc7282726043b2aadedeb8f4c706cb1;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1aab056e04334a2b3c4735882750d6b1bb0780e270378be9c57c5da7fd0c1423164c7c2c2f48b95835368741c87013da7fd6;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fb29b6f6573a04497acff9dc90e111e2f38e4b34801bbd9f6c206b349cd16d9a5cf13aaa357119437b954ee307452962b3c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he80ba56b9007d1980d15e9ff5e55de5933687499c4dc0b46c8c2fb93d2cb0faf07464efa231c2432c59c0bc2270a0445e48a;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he2d6b31d7c411f10aae81071bdc8eb35587f1278d5aed71fa68530ed1820146f925dfc844e66ad14ee2bcd17994a488b355e;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6da2d824bd6f8ed2747eb4b31d5f8833ba280a2f4cb8d00f2191749dfa663a16f9bab1360d34e2019761fdd3e2ce32d91d6c;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h977b719aa06e375c6771f5893df27bd072841ad09fed8ffb475612c41cdc20770daaee2f5a42c471316711b5405af4ca59cd;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacb1bd582bb4c0f69ca627a13830ba69d7f79661a23e155bd6d4346ae59f971d0b481eb5cd2aa6f8b4a82ad7e471856ab9ce;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h43b50816d7e8003ef73fb5148285036d7804398acc3527305b47b92f3d310f9f92c3800982b93f30f7ea33e83e24e2d8cc50;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6df6b38c785ffa0e9fc2bc5c9f424c021400425c2cbcb3947c6329e8241fe2b2b8e38a67e255386bd83e19e60b1b3369472;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h206c91eea8e2e0ef023e73e44da48fc86bcee534cddfef55d6863fa66f8f30e09e09a5b17f25c78de98175f8c0f7a0deb734;
        #1
        {src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cb169344ff53ad86468b7fa7963b34ca662c2ab5cc97e545c333284de590e4b6c5e6ece102ccc7fd51f18cbf1dc9418234f;
        #1
        $finish();
    end
endmodule
