module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17);
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    compressor2_1_54_12 compressor2_1_54_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17));
    initial begin
        src0 <= 54'h0;
        src1 <= 54'h0;
        src2 <= 54'h0;
        src3 <= 54'h0;
        src4 <= 54'h0;
        src5 <= 54'h0;
        src6 <= 54'h0;
        src7 <= 54'h0;
        src8 <= 54'h0;
        src9 <= 54'h0;
        src10 <= 54'h0;
        src11 <= 54'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor2_1_54_12(
    input [53:0]src0,
    input [53:0]src1,
    input [53:0]src2,
    input [53:0]src3,
    input [53:0]src4,
    input [53:0]src5,
    input [53:0]src6,
    input [53:0]src7,
    input [53:0]src8,
    input [53:0]src9,
    input [53:0]src10,
    input [53:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16)
    );
    rowadder2_1_17 rowadder2_1inst(
        .src0({comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0({dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [17:0] stage1_0;
   wire [17:0] stage1_1;
   wire [17:0] stage1_2;
   wire [17:0] stage1_3;
   wire [25:0] stage1_4;
   wire [29:0] stage1_5;
   wire [18:0] stage1_6;
   wire [17:0] stage1_7;
   wire [26:0] stage1_8;
   wire [25:0] stage1_9;
   wire [19:0] stage1_10;
   wire [24:0] stage1_11;
   wire [16:0] stage1_12;
   wire [6:0] stage1_13;
   wire [7:0] stage2_0;
   wire [8:0] stage2_1;
   wire [5:0] stage2_2;
   wire [7:0] stage2_3;
   wire [11:0] stage2_4;
   wire [7:0] stage2_5;
   wire [12:0] stage2_6;
   wire [10:0] stage2_7;
   wire [7:0] stage2_8;
   wire [11:0] stage2_9;
   wire [10:0] stage2_10;
   wire [7:0] stage2_11;
   wire [12:0] stage2_12;
   wire [6:0] stage2_13;
   wire [2:0] stage2_14;
   wire [0:0] stage2_15;
   wire [3:0] stage3_0;
   wire [6:0] stage3_1;
   wire [5:0] stage3_2;
   wire [1:0] stage3_3;
   wire [5:0] stage3_4;
   wire [2:0] stage3_5;
   wire [3:0] stage3_6;
   wire [5:0] stage3_7;
   wire [4:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [2:0] stage3_14;
   wire [1:0] stage3_15;
   wire [0:0] stage3_16;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc615_5 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_1[0]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc615_5 gpc5 (
      {stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33]},
      {stage0_1[1]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc615_5 gpc6 (
      {stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_1[2]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc615_5 gpc7 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43]},
      {stage0_1[3]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39]},
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35]},
      {stage1_5[5],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45]},
      {stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage1_5[6],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[7],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc615_5 gpc16 (
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52]},
      {stage0_3[48]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[8],stage1_4[16],stage1_3[16],stage1_2[16]}
   );
   gpc615_5 gpc17 (
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage0_4[6]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[1],stage1_5[9],stage1_4[17],stage1_3[17]}
   );
   gpc606_5 gpc18 (
      {stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[2],stage1_5[10],stage1_4[18]}
   );
   gpc606_5 gpc19 (
      {stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[3],stage1_5[11],stage1_4[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[4],stage1_5[12],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[5],stage1_5[13],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[6],stage1_5[14],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[7],stage1_5[15],stage1_4[23]}
   );
   gpc606_5 gpc24 (
      {stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[8],stage1_5[16],stage1_4[24]}
   );
   gpc615_5 gpc25 (
      {stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_5[6]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[8],stage1_6[9],stage1_5[17],stage1_4[25]}
   );
   gpc606_5 gpc26 (
      {stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[8],stage1_7[9],stage1_6[10],stage1_5[18]}
   );
   gpc606_5 gpc27 (
      {stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[9],stage1_7[10],stage1_6[11],stage1_5[19]}
   );
   gpc606_5 gpc28 (
      {stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[10],stage1_7[11],stage1_6[12],stage1_5[20]}
   );
   gpc615_5 gpc29 (
      {stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_6[48]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[11],stage1_7[12],stage1_6[13],stage1_5[21]}
   );
   gpc615_5 gpc30 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34]},
      {stage0_6[49]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[12],stage1_7[13],stage1_6[14],stage1_5[22]}
   );
   gpc615_5 gpc31 (
      {stage0_5[35], stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39]},
      {stage0_6[50]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[13],stage1_7[14],stage1_6[15],stage1_5[23]}
   );
   gpc615_5 gpc32 (
      {stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43], stage0_5[44]},
      {stage0_6[51]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[14],stage1_7[15],stage1_6[16],stage1_5[24]}
   );
   gpc615_5 gpc33 (
      {stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49]},
      {stage0_6[52]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[15],stage1_7[16],stage1_6[17],stage1_5[25]}
   );
   gpc606_5 gpc34 (
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[0],stage1_9[8],stage1_8[16],stage1_7[17]}
   );
   gpc2135_5 gpc35 (
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4]},
      {stage0_9[6], stage0_9[7], stage0_9[8]},
      {stage0_10[0]},
      {stage0_11[0], stage0_11[1]},
      {stage1_12[0],stage1_11[1],stage1_10[1],stage1_9[9],stage1_8[17]}
   );
   gpc2135_5 gpc36 (
      {stage0_8[5], stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9]},
      {stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_10[1]},
      {stage0_11[2], stage0_11[3]},
      {stage1_12[1],stage1_11[2],stage1_10[2],stage1_9[10],stage1_8[18]}
   );
   gpc1406_5 gpc37 (
      {stage0_8[10], stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage0_11[4]},
      {stage1_12[2],stage1_11[3],stage1_10[3],stage1_9[11],stage1_8[19]}
   );
   gpc606_5 gpc38 (
      {stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[3],stage1_11[4],stage1_10[4],stage1_9[12],stage1_8[20]}
   );
   gpc606_5 gpc39 (
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[4],stage1_11[5],stage1_10[5],stage1_9[13],stage1_8[21]}
   );
   gpc606_5 gpc40 (
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[5],stage1_11[6],stage1_10[6],stage1_9[14],stage1_8[22]}
   );
   gpc615_5 gpc41 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38]},
      {stage0_9[12]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[6],stage1_11[7],stage1_10[7],stage1_9[15],stage1_8[23]}
   );
   gpc615_5 gpc42 (
      {stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_9[13]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[7],stage1_11[8],stage1_10[8],stage1_9[16],stage1_8[24]}
   );
   gpc615_5 gpc43 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_9[14]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[8],stage1_11[9],stage1_10[9],stage1_9[17],stage1_8[25]}
   );
   gpc615_5 gpc44 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_9[15]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[9],stage1_11[10],stage1_10[10],stage1_9[18],stage1_8[26]}
   );
   gpc606_5 gpc45 (
      {stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_11[5], stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10]},
      {stage1_13[0],stage1_12[10],stage1_11[11],stage1_10[11],stage1_9[19]}
   );
   gpc606_5 gpc46 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27]},
      {stage0_11[11], stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16]},
      {stage1_13[1],stage1_12[11],stage1_11[12],stage1_10[12],stage1_9[20]}
   );
   gpc606_5 gpc47 (
      {stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33]},
      {stage0_11[17], stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22]},
      {stage1_13[2],stage1_12[12],stage1_11[13],stage1_10[13],stage1_9[21]}
   );
   gpc615_5 gpc48 (
      {stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38]},
      {stage0_10[48]},
      {stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28]},
      {stage1_13[3],stage1_12[13],stage1_11[14],stage1_10[14],stage1_9[22]}
   );
   gpc615_5 gpc49 (
      {stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_10[49]},
      {stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34]},
      {stage1_13[4],stage1_12[14],stage1_11[15],stage1_10[15],stage1_9[23]}
   );
   gpc615_5 gpc50 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48]},
      {stage0_10[50]},
      {stage0_11[35], stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40]},
      {stage1_13[5],stage1_12[15],stage1_11[16],stage1_10[16],stage1_9[24]}
   );
   gpc615_5 gpc51 (
      {stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_10[51]},
      {stage0_11[41], stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46]},
      {stage1_13[6],stage1_12[16],stage1_11[17],stage1_10[17],stage1_9[25]}
   );
   gpc1_1 gpc52 (
      {stage0_0[44]},
      {stage1_0[8]}
   );
   gpc1_1 gpc53 (
      {stage0_0[45]},
      {stage1_0[9]}
   );
   gpc1_1 gpc54 (
      {stage0_0[46]},
      {stage1_0[10]}
   );
   gpc1_1 gpc55 (
      {stage0_0[47]},
      {stage1_0[11]}
   );
   gpc1_1 gpc56 (
      {stage0_0[48]},
      {stage1_0[12]}
   );
   gpc1_1 gpc57 (
      {stage0_0[49]},
      {stage1_0[13]}
   );
   gpc1_1 gpc58 (
      {stage0_0[50]},
      {stage1_0[14]}
   );
   gpc1_1 gpc59 (
      {stage0_0[51]},
      {stage1_0[15]}
   );
   gpc1_1 gpc60 (
      {stage0_0[52]},
      {stage1_0[16]}
   );
   gpc1_1 gpc61 (
      {stage0_0[53]},
      {stage1_0[17]}
   );
   gpc1_1 gpc62 (
      {stage0_1[52]},
      {stage1_1[16]}
   );
   gpc1_1 gpc63 (
      {stage0_1[53]},
      {stage1_1[17]}
   );
   gpc1_1 gpc64 (
      {stage0_2[53]},
      {stage1_2[17]}
   );
   gpc1_1 gpc65 (
      {stage0_5[50]},
      {stage1_5[26]}
   );
   gpc1_1 gpc66 (
      {stage0_5[51]},
      {stage1_5[27]}
   );
   gpc1_1 gpc67 (
      {stage0_5[52]},
      {stage1_5[28]}
   );
   gpc1_1 gpc68 (
      {stage0_5[53]},
      {stage1_5[29]}
   );
   gpc1_1 gpc69 (
      {stage0_6[53]},
      {stage1_6[18]}
   );
   gpc1_1 gpc70 (
      {stage0_10[52]},
      {stage1_10[18]}
   );
   gpc1_1 gpc71 (
      {stage0_10[53]},
      {stage1_10[19]}
   );
   gpc1_1 gpc72 (
      {stage0_11[47]},
      {stage1_11[18]}
   );
   gpc1_1 gpc73 (
      {stage0_11[48]},
      {stage1_11[19]}
   );
   gpc1_1 gpc74 (
      {stage0_11[49]},
      {stage1_11[20]}
   );
   gpc1_1 gpc75 (
      {stage0_11[50]},
      {stage1_11[21]}
   );
   gpc1_1 gpc76 (
      {stage0_11[51]},
      {stage1_11[22]}
   );
   gpc1_1 gpc77 (
      {stage0_11[52]},
      {stage1_11[23]}
   );
   gpc1_1 gpc78 (
      {stage0_11[53]},
      {stage1_11[24]}
   );
   gpc2135_5 gpc79 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc80 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc81 (
      {stage1_0[10], stage1_0[11], stage1_0[12]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[2]},
      {stage1_3[4]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc615_5 gpc82 (
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7]},
      {stage1_3[5]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3]}
   );
   gpc615_5 gpc83 (
      {stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage1_3[6]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc615_5 gpc84 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_3[7]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc85 (
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage1_4[18]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[3],stage2_5[3],stage2_4[6],stage2_3[6]}
   );
   gpc615_5 gpc86 (
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage1_4[19]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[4],stage2_5[4],stage2_4[7],stage2_3[7]}
   );
   gpc1163_5 gpc87 (
      {stage1_4[20], stage1_4[21], stage1_4[22]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[2],stage2_6[5],stage2_5[5],stage2_4[8]}
   );
   gpc606_5 gpc88 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[1],stage2_7[3],stage2_6[6],stage2_5[6]}
   );
   gpc606_5 gpc89 (
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage2_9[1],stage2_8[2],stage2_7[4],stage2_6[7],stage2_5[7]}
   );
   gpc606_5 gpc90 (
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[2],stage2_8[3],stage2_7[5],stage2_6[8]}
   );
   gpc615_5 gpc91 (
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage1_7[13]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[3],stage2_8[4],stage2_7[6],stage2_6[9]}
   );
   gpc615_5 gpc92 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[14]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[4],stage2_8[5],stage2_7[7],stage2_6[10]}
   );
   gpc1163_5 gpc93 (
      {stage1_8[18], stage1_8[19], stage1_8[20]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_10[0]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[0],stage2_10[3],stage2_9[5],stage2_8[6]}
   );
   gpc606_5 gpc94 (
      {stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26]},
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage2_12[1],stage2_11[1],stage2_10[4],stage2_9[6],stage2_8[7]}
   );
   gpc606_5 gpc95 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6]},
      {stage2_13[0],stage2_12[2],stage2_11[2],stage2_10[5],stage2_9[7]}
   );
   gpc606_5 gpc96 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[1],stage2_12[3],stage2_11[3],stage2_10[6],stage2_9[8]}
   );
   gpc606_5 gpc97 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[2],stage2_12[4],stage2_11[4],stage2_10[7],stage2_9[9]}
   );
   gpc606_5 gpc98 (
      {stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[3],stage2_12[5],stage2_11[5],stage2_10[8]}
   );
   gpc606_5 gpc99 (
      {stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17], stage1_10[18]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[4],stage2_12[6],stage2_11[6],stage2_10[9]}
   );
   gpc606_5 gpc100 (
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[2],stage2_13[5],stage2_12[7],stage2_11[7]}
   );
   gpc1_1 gpc101 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc102 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc103 (
      {stage1_0[15]},
      {stage2_0[5]}
   );
   gpc1_1 gpc104 (
      {stage1_0[16]},
      {stage2_0[6]}
   );
   gpc1_1 gpc105 (
      {stage1_0[17]},
      {stage2_0[7]}
   );
   gpc1_1 gpc106 (
      {stage1_1[12]},
      {stage2_1[3]}
   );
   gpc1_1 gpc107 (
      {stage1_1[13]},
      {stage2_1[4]}
   );
   gpc1_1 gpc108 (
      {stage1_1[14]},
      {stage2_1[5]}
   );
   gpc1_1 gpc109 (
      {stage1_1[15]},
      {stage2_1[6]}
   );
   gpc1_1 gpc110 (
      {stage1_1[16]},
      {stage2_1[7]}
   );
   gpc1_1 gpc111 (
      {stage1_1[17]},
      {stage2_1[8]}
   );
   gpc1_1 gpc112 (
      {stage1_4[23]},
      {stage2_4[9]}
   );
   gpc1_1 gpc113 (
      {stage1_4[24]},
      {stage2_4[10]}
   );
   gpc1_1 gpc114 (
      {stage1_4[25]},
      {stage2_4[11]}
   );
   gpc1_1 gpc115 (
      {stage1_6[17]},
      {stage2_6[11]}
   );
   gpc1_1 gpc116 (
      {stage1_6[18]},
      {stage2_6[12]}
   );
   gpc1_1 gpc117 (
      {stage1_7[15]},
      {stage2_7[8]}
   );
   gpc1_1 gpc118 (
      {stage1_7[16]},
      {stage2_7[9]}
   );
   gpc1_1 gpc119 (
      {stage1_7[17]},
      {stage2_7[10]}
   );
   gpc1_1 gpc120 (
      {stage1_9[24]},
      {stage2_9[10]}
   );
   gpc1_1 gpc121 (
      {stage1_9[25]},
      {stage2_9[11]}
   );
   gpc1_1 gpc122 (
      {stage1_10[19]},
      {stage2_10[10]}
   );
   gpc1_1 gpc123 (
      {stage1_12[12]},
      {stage2_12[8]}
   );
   gpc1_1 gpc124 (
      {stage1_12[13]},
      {stage2_12[9]}
   );
   gpc1_1 gpc125 (
      {stage1_12[14]},
      {stage2_12[10]}
   );
   gpc1_1 gpc126 (
      {stage1_12[15]},
      {stage2_12[11]}
   );
   gpc1_1 gpc127 (
      {stage1_12[16]},
      {stage2_12[12]}
   );
   gpc1_1 gpc128 (
      {stage1_13[6]},
      {stage2_13[6]}
   );
   gpc2135_5 gpc129 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc130 (
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1]}
   );
   gpc615_5 gpc131 (
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4]},
      {stage2_5[6]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[2]}
   );
   gpc615_5 gpc132 (
      {stage2_4[5], stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9]},
      {stage2_5[7]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[2],stage3_6[2],stage3_5[2],stage3_4[3]}
   );
   gpc615_5 gpc133 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[3]}
   );
   gpc615_5 gpc134 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[4]}
   );
   gpc606_5 gpc135 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[2],stage3_9[2],stage3_8[4]}
   );
   gpc615_5 gpc136 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10]},
      {stage2_11[0]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[1],stage3_11[3],stage3_10[3]}
   );
   gpc606_5 gpc137 (
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[1],stage3_12[2],stage3_11[4]}
   );
   gpc1325_5 gpc138 (
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10]},
      {stage2_13[6], 1'b0},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[1],stage3_14[2],stage3_13[2],stage3_12[3]}
   );
   gpc1_1 gpc139 (
      {stage2_0[5]},
      {stage3_0[1]}
   );
   gpc1_1 gpc140 (
      {stage2_0[6]},
      {stage3_0[2]}
   );
   gpc1_1 gpc141 (
      {stage2_0[7]},
      {stage3_0[3]}
   );
   gpc1_1 gpc142 (
      {stage2_1[3]},
      {stage3_1[1]}
   );
   gpc1_1 gpc143 (
      {stage2_1[4]},
      {stage3_1[2]}
   );
   gpc1_1 gpc144 (
      {stage2_1[5]},
      {stage3_1[3]}
   );
   gpc1_1 gpc145 (
      {stage2_1[6]},
      {stage3_1[4]}
   );
   gpc1_1 gpc146 (
      {stage2_1[7]},
      {stage3_1[5]}
   );
   gpc1_1 gpc147 (
      {stage2_1[8]},
      {stage3_1[6]}
   );
   gpc1_1 gpc148 (
      {stage2_2[1]},
      {stage3_2[1]}
   );
   gpc1_1 gpc149 (
      {stage2_2[2]},
      {stage3_2[2]}
   );
   gpc1_1 gpc150 (
      {stage2_2[3]},
      {stage3_2[3]}
   );
   gpc1_1 gpc151 (
      {stage2_2[4]},
      {stage3_2[4]}
   );
   gpc1_1 gpc152 (
      {stage2_2[5]},
      {stage3_2[5]}
   );
   gpc1_1 gpc153 (
      {stage2_4[10]},
      {stage3_4[4]}
   );
   gpc1_1 gpc154 (
      {stage2_4[11]},
      {stage3_4[5]}
   );
   gpc1_1 gpc155 (
      {stage2_6[12]},
      {stage3_6[3]}
   );
   gpc1_1 gpc156 (
      {stage2_7[10]},
      {stage3_7[5]}
   );
   gpc1_1 gpc157 (
      {stage2_11[7]},
      {stage3_11[5]}
   );
   gpc1_1 gpc158 (
      {stage2_12[11]},
      {stage3_12[4]}
   );
   gpc1_1 gpc159 (
      {stage2_12[12]},
      {stage3_12[5]}
   );
   gpc1163_5 gpc160 (
      {stage3_0[0], stage3_0[1], stage3_0[2]},
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_2[0]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc161 (
      {stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage3_3[1]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc1343_5 gpc162 (
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[0], stage3_7[1], stage3_7[2]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1]}
   );
   gpc1343_5 gpc163 (
      {stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc164 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc165 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], stage3_14[2]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc1_1 gpc166 (
      {stage3_0[3]},
      {stage4_0[1]}
   );
   gpc1_1 gpc167 (
      {stage3_1[6]},
      {stage4_1[1]}
   );
   gpc1_1 gpc168 (
      {stage3_15[1]},
      {stage4_15[1]}
   );
   gpc1_1 gpc169 (
      {stage3_16[0]},
      {stage4_16[1]}
   );
endmodule
module rowadder2_1_17(input [16:0] src0, input [16:0] src1, output [17:0] dst0);
    wire [16:0] gene;
    wire [16:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[16:16]}),
        .S({3'h0, prop[16:16]})
    );
    assign dst0 = {carryout[16], out[16:0]};
endmodule


module testbench();
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor2_1_54_12 compressor2_1_54_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h6854f6759e3047d555cfd716c7d00af99b98bf22da96ba80c5b4b823e981b74d314b7c19fc69f3e7031628eea6dd1b85094e655618fecab5ca1e663ba3e1bbdfeee6cc20a91cf83a69de7bd12617f9f4e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h55f62448d9eb69c5a3a539b4efd50c1f8f2cb3d0bcc6af4029a230d2a6b3a935c6f88debdf483e67166b25916c5a76d62f9e1aed11e8d0b8728554302620c02a066be871fb35d7cc85055b40198598e1a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'he4f54cc1b3c56ce33bdb59627a4be29275610504b4e4040a2193539a3d5715fb534946b026875471db021a6ee94e21a6f14ff177c39ef850ec902b77b58f85205e52a9393b8acdb0fddffab00391891e3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hee078d1cd3f13ea77b76b7cc4d0a2a3f2ec8fe353d8b43c26225a2c7156d8a6ecd023ea2459715612b791389d8b5083974cbe15625096bd854d52285af96651c9ca5c380fb70c32e8e981fe9c36b1a8fba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'ha5688dd8329d71c5c97bb77907876ebc9e2b55a1194c88997d0e639eeb10b5ffcd1322aace40e74ae6b4fff1a431e65e54f3936190b79ffadc35c2299b32d612854de4ef8e41361e3b29b95a0fdbe62692;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h4fc561d18cbeb3c4972d71c91205ff4594e2cac91ca7c55005a2b417fd8110fbb229467b5d5efcd750151c696b9eb0886cd0cdf4c1c52b6eb95e8c448728e426aca3bdd9303dbcc4eb9841d21b60ccc32d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hae2cd90813905f1b925fdcf24cead613c48d2a3776d0686635b47f1ba5b07cf620c586c50cd1ca7f3079d157f7accce191f6e083f70186157070fc8de6c9729cc807def08e53c64d38c4ef131090634d34;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hdda3c8b15a2e01e2eeca30cbb4a5ce44721a4315dd4a39e533053e2b3ca04ba097b86eef41217f00013d81684d3c022eec74a580388caa0385bfa52cd684de213ffe60877d3ef3c7c8190e88f008cb8255;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h4fb70355e1f72c5e6028f47eeffc80c8769179214f4c0f7e48276de923db2f4e860d62137a485f33bbaf8f3b2508d3cae330ef0dbe744f665cf90f491ef786988c1da87fbbd94765863fb1897f592ffa37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h46217187eadbb1336e11eec9e037982253bc95f41dc054bb257f171aef02bcec7c018fecfceaea94c4c559a297f6bbdf70e6c77ca2c65223d3bd40d80fcf65e3e62a06c37791e86df0fee8b2e59c04c3ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h69f86162107df8db18b75a4f4ae2ac93964eba26ba6634c8e9c017154371343a01b680c2347b551f4402905379cf635d62cbac7599e26c302043add913f967948d38551516664fb79403fedfd090884c96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hf5a009ea4e5a83d49537333216059a7631b97254ae94924bd5afcbaf646d29b0fda83e4a781245fc5d05dee6afda6fd4049a18d31dfde32444b50cc766d897829355f4e73cfc32e6aa102bfb29f344ba61;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9741154b521a2acd5c5c24bbcfe069660147b2b691e93b30a199bd1d0d27f9e85980e0da9b1d39985bdddbae47d723060a3c3119d3bc697e4ed62228dea2c1d8efc2f318c1ec2098c09f431ea8e54c58d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hf01c1fe8b38848d5b66aa3e6198be0a1f764c12180c1e138bbaa8f8f4ce8bfae5b68bb3c9dc1aaff04c56461ed0718b38cc074e755b1ff4a55d098aa34a3ef599e99ac1f419e2dcbe632cc8a09e9d3528c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb5906330158e534bbff68faf117ae0a6d0932b4c5c163607cba5f8bb33bd394ad9c602fc813e7281346c95a67e42bb2ed632522920bab6b16f578b5b4a93185edf2f70d2e91dbd2268e7ea12fad1499245;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hef66caec607f9957c497c5753737aebc0c3124c522762e6a49eff97e7e4c2f08799b6cb853e220fe4efa6ff33505d0aaf736041d60c566e57a3f1f9bb1581daea32b8b8716dd0b94a5c1bec7bebb0409da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hf9cc55e236770d693178256226b9239883319f130ef94ab56208d50c0b638368557c1fae34055771be0ebef79604105d38345c57299e3de1991087e6ede5c94b352e72a4e5dcaa608b3acadd87acbad763;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h604b9157fa963fdd72c419c82fefb9af5fa5b15f9f827ced44236c0a87381df6c2533266a6f6579ec1ef74a27b7c593036b1c09d5846c6cf4697423d2a7aabea01f60a3f91f78f0ebab1b9e1e585ee0793;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb8ecb02c5b4e283a47d1bd44e7ec96f034b311ef443c72400e03715a4921153a26ccdc97ca8700eed6618a2fad564264020a25932d505d3d94f26c2d8fd95f34d605dbbe047ae34f0788fc64c52dc697e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h677bd78f78278c6de8e695279fe88de40804120a7ecfe6078ebdc00b0abafc88b2bd4b8ceb6a552582dc8b8f77fabeac219cf03974e1dfcdacaa047f2b1133680a9f6126be1c281387a8ccb852f1505c33;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9354a929997e27f841b01de130c6ad0909da5692af47b87f2d84a51486ed96ad79c7cd338063bc382f59d4e0b30bdbdffb0d9688b1f5d6f2cd396b1b1998049ddf031d2c6afe756a2b57441880c09fa3f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hfaa7d506b2d7f654adee505074149896d512e3a3fd8cb4a3e9f1558deafb1c268d78af11c783e61fdb3e4964edb4d78cac296571212c4d0290b1cd87aa448024314462f7d2d0d158bcb2ac2824eb3a88a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9fc8420f26d06e3c4f3c2a3099b8b22a20f1c90b77fd5f2900a7e3898bbb200c53a2794ee238548bcc46e831af9f23b1b529d27d2284e59daef6aa44f52cfe82db3ccaacdaee9c911b0f3910a964807fac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h6f4a7e1bca0fe317fbec126f3a482c3a574ee0cc3edebdf23a65178c6f20c9e3910286415aff55d003391883c9abfea6ef03367b3f2b14638410e32a7e4bd61b13925adf01b6f5bfa3d3453d8dae041963;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h1aefe5fe75695ba9ec6bbfa0cc908584eacbb65e61eda1884bdc89428bbdd2b55b805be3b11603ab2074ef35a3916c3eac304a972d784e1e888e040e4cca3327939ccb6b46018c2aef38168665bc6dc00b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h5739010a73d137e36a7b89f1cf078c5e15db4fb6f576965b30532f33ec12b461b83b0363bafe7264c01910640f68cd77dac6ffa4f002ca0c87191933afe2055bd92a3c8aea3c285a27b7a4726983dd5d4f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h3263733eb0fd837d52a13247f413d4a21c654b2be18f99ec6235ffab06cff0e5a456146b73ff1743d43ea1531132092f20a9b9513b86f539a1e08dfd00cbfc879797c7b13d2d322da3b2126445f4b6f7de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h923759b72ade9ac203ae5fa6e2b3d2908f50eea5f00bd93ab0e130354e0bd582fcf79474d703539a571c17957cc3609de7721e58605417fd5fcf1120753fa90a18b8f24b76612e2debf684f71cfdb3ecfb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h5d908827801fceeb6f192cf1973bc308a7415d49701d92c61889195ca3dfe26f0d9be1a92d3ef6f94e4e0d8a1cd4f7ac042f41595e875b73d4df94a5355f197b4cfb665d0d798838991a5057e08d4ca3a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hdcf6af1306ad33f07ac25b5ab0ead76f59dc539352217e46d660a3071b9393bcd7356e7a6e933a9c89ca078c110e14c331c4392069b4e9dbf34651249e1c7055ca19654c9af1279418aae21b6c2d1fab1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'he6d501a2605bc6287467ab770f2d5779a338337e89d95c5a8ce19a7b0f7135f48dbb1fa39f856ffe51997221efea22f8b57d338941a7d5d414fc9e0e75c4f24f8d2edec8016594e094d9115bc2605ba1d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hec52dd30695b3cc8476ff1014772965e5fd110b8fe10a87862a6f5e9ca311b8fb53807d14f65fcde596a9546e2ed3054d200f079ac8bba16599d6d08f99e9f92afa13657697b0f93de4c71725d7fd69a7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h68865d882c259858eb7eb601cdb4f6579775764ceee1ee199732490e76cd034bfd01cda23425d5aabe27e549ec86352d7f08e63c52e29a6752f8ed6e4fbb92a2ae94513a3ca3207dfed8325ae7a1e2a3c6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h1f95d0b717123f43addac743b07df4a92e7e007676615e2570984f24048c7c2eb0d6374ea21f9df8f3d8add4664f8a5471d0c65a6474da19414840b9a2a0aa0d488a8de3eb11c1b601ffc1aca6ba60e42a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h6207b5678ade3b6909ac6cf92894948418019edc9d1dbaecc835ffba22040a43003940f9a85bb5777a9c9785c67bfdcdaa3d9d60e0b7a02497f1d03d782e3112e21c274f3f30b97068cef0fbec318c6f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9f58ce88a50e26862d159c58dd5282f547425fbcfd7d86bc2bc1a6caa79e5d1d8276224a6856e2d62b3b5e3fe67818664cfbddf9dc8333e8fa4bfdd5436bc766d4c0d974ba116d4ee8a320b3688c782e37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'ha910f587fc92dc2406ad9da7ddc1fcd9de460bfaf25fc9688f78e4f7ef3686d26bf84edc722df40b7467f708e5a147718fa88eb0c56d39d69fc7c300710eb826d14cc4badfff492b8b7545cec919523209;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h4387458e86256f4ddfc3d0f1152a926ce4f2363bad289801c7a65b72ba4a8fd8541b6582ae648f09fe701630c6b1c59824050a7cc8695587bef6e9f2de2e9e2f6beef145b520aa309b038cb31fab5da140;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7708188f085a4e1fd6de832c5ec92b9407a9c49507068a5bbeeced393b3d51cbcda52e216c0368f22162e04b442518a40c7d7be75ef36149c24d41afa5e97e511d4bcdb649120e9e3f6cba991f9351ffae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'ha0062465abc2d09e4d223c9ac0cb98bf6c9b5f6bb6b6054cc67c8ab3cf9571477d9b2e3ffc06a3573399ac1c00b22d01d8d21d077fd39605e28fd3a35bb273298c2b4e32a88e6d8ea88b24f5cef982b753;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h117bc9b661953b9c1b1427133d0535b558a3187633a5a8e00d6d67d2a02e23d2abea4794842bac56195ae3b5cd97a67f93f465f4736afe536444b32a8718bf413a4a41771da72c9721934f743b7c1b8cc0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h35c4f87a7fdc0c33665c28d8314b4409fd26d162ce1b3f13767a31c1180e57585989fa64796cd0c3a074910946439a91a296f8b15168c972bf5b6bb91a7ab3f008b14b62828c48b204aeb26fbcf1149897;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb811d9127bd465c385c3ce418c44e4f4189de5794ea7e6208a946bd69ebc387bb6a595055e3d2e315cbc82815985210c286706236132a7d5653b2b89c560ac79e8edc4d92ef53011d6b2d1573a3e46365d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hbf26c3cc8c11527156c77f759e9bb4e9b739f06db428240fc30e2fa83a02447368fcbce82f2827f5acc2599d6ec2858e933ef405eda4de4be939c3a8a4a67e67222a4d0e15cba0999a00aecd4096f90dc8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hed9fe6d97845c28d222cac550827a8ddbb724cf0691909fb46829c1510cc57f0dcfe519deaeb3a1f2370a63837c5c23c0ea836cc11e7a979d32335e9c70624e4c1adede2f5eeedb9ee28546e982f4a6823;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7ad9629b9879fb850fe120b516353cf94be75b33515a7d9b9ddaf046f05134d7953a3b0283cae8d856ce9580190269dfafcbe9217094428eb097d31c0a813bd556ff198deb99aded209510f81a3c0cd8f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hd1289c33e0adbf0946bdd26bacbafdee6a618d064b471d281bb81f36b2b7fdcbdb68f0cfbb4a3b64f432e8dc534334ef6898f5c2ce3a048eebeec4030da088636f13ef0f9b615fe20d309dd05358599a10;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9185b23bac359bfa6a5b4825d86895fc1e554a5b951ea0be0609b6cfafc762e928adc0ce4d86ad500165aa085ed90763723091f9d37f978a6875164da1818b02dcc3b910acd2373f6d4ba794ec23dad93;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h70068ea6697b8e322c7a215f2cdc3a74bb2b5614ba516cc155126dab4ec75c38e1111fda86035e29493f4b002ffb36e5e211a6cd041b5cf9de0954df603ce876e0b82b0c298542b7ecc6b9c06f731189bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'heefe6dd7b1b1549048fb544b64f00a155f66e2986e4a61818c575e1a5079ed7826d8c9a27b7f9afda736ddc7dbd184aece5f6930e45597f56f1b3de8da38b86d099ac1750ca37dbfebf52523139ec6c27e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'heb1188dc6a86e49635aecf6a96e9ea97f1c36b5dc2b44eced9e66fdc88200e525de932d4dc7137d66253b5cc3d4e127df17dff430fab3883a54ca4694883afbe315a06a1159f62383c3c986ee97f4fb7e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hc5b59220bf818b68a66191f5e6d10513f75a83eea818bc7ed15c6d2ef09d6f7837243df5c45e2a834dafe1422689b2cbb5f10b76012eb8a06a3c0662eb298f0d2c2b8d50e2b4101a39a5a50fc9bc8c8ac2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h1501b9e1dcd597a485c79ee0712571f67cedbd7c6b8b28e2500545c6646a2c2fb8a45d5719f072345c7656e104171a61d679736e0dda4cc4cd186906711f2d1e9741d354b92f07aa7e4a59abc51ef42db2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7e5d877327802ad212924101ecc680422d3c659d8a28ab1d8a0aa8fd9385c7c8825969d67bd446a560db3f83ca317e52fb80ad53da31e2bd241ae4da5120aa69d8c1e6c3df41a3841d5259d25a53d1587e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h90e4fab544a7b45c401533b00fed0ebe0f4b56f240c619f6ab604edc6c1cbf65801026ffb90fd21b5e2f9e9ef817c15d773aa9b0c8202e026d627e050c00c6dd7556419a9e161367855a3f759389bb0f49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h394516e8cb381045d5ed1030b6a93b2e50e471b25cbffbf978fbbdc59f34bd9dece921b8ee59aa611aba6a41eab8f6c0c9a73c367b0e584903b5df690e0deef38c8c320ac945003db62fd662a268157a02;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h19a8db13de03fd890c50213bfe33895d4f7e75049c8fdda13fadecc8115c59d5470d39af4dd0038bd5f0468c9cb9fbf97efe0604b7fc45aa43debb721a417cb389947ca4e31c5cf39bf6088d5069a5920b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h92f8f4a5aceeabeca66303bd8412a861d72aa273a4d0536066a41a80c5cbb78d313e539b815df179eea691302cd43c383e70840904ac1deb93c7b17769310c1bd005c2ec8e12430a294b189cf70e3e3f30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h141d661de11235cb4644a1a12dd1b81cd769aa7d699f120caebf7a0c008a1b03b47bc1f8bf93e4d2adb514e74c9993d1711bf9edec68f6ec24d103c4241400058a887d7f752b9cc05c9a7b34071e25ee9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb74621eea22cb33e51a686df5bb12cc0fa3896417e5ce4461cd3d6e3644ca7ece1fef32f443f9815b1efb3476db5931f985db52bcf14dd28605c2fe43517591d829c62d8e8b98152bc3851180409a8d9bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h13828a0bb8f9c1085354a21d5477e539f358950f011281008b39b8ede031020cfec561be528297c88aadf2885fbfa34f4ae37159044dc56657fbb86073539afcd90ce7f1cc8e865dac0b7837ecdc8bec3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h7f01a04cf8eb2d0b6c963c2e7a6037d40fcc2df1e034484bac8d2f6585de4577b08ce9be9dffbf6c9f01e8fd34561e6acf5dda66e2d1422b7b692965625db373cd4b5e8875ba93c4f23843df74d91fb883;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hffd9dff982752d5f09eb87c6c7fc90ec16bf91eba431ff9e65de4ad93fa4ecb0d3d1a8e361685aedb5b888e60f161b8f3191d9e9a054bd3dbeda6aa97c6560ee0de376b9d1fe48033084a7f6725b6a0a1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h380b32f7b69fc03295b4b3e04564e16edef5464d4bce6b1b05d049547c6bdf526a6d8f78097daa1669df68d14255aaafe855c55bb7a6a18685033ba81f12dae7bc61ac4d85aecbc36bab9de317945ffdd9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'haa977104014674cd275b791c090a98ffee8bf9c8264f9852ac4858c1bf0c9444487daef3fe21d941e495bfb2f3b48829a1a8aa97a4cba9e11bd9af796d0948cd5fdea0b31a8c5898c0045844658f31b6fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h5759c94759c97b9ea2e6a6baa7724f61d72147df55efe7fcdee880a27b9ff15efc6bc9e33c9998a5a1b9c308df81b4ff0e52fc44a156a7ccf46af8e80bd43c2f6ce1ee5fbc8033878d38e035e2d6e0ba78;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h8269996ccd6a7ff266c029aac85ae74fcb56783de3bc9cd35fe9920dae1df9f5baa430c9ce8c75bdc28101d2f78b81b5e61752e1ce129ea4aeff097c7d2952128c3a954ca5b7e20b8900f2990cdbcd47b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h6df98a8f409662116f91698a8b0c70c2d296647e4e22f10e74866f4c6a9403ac8f4072a7caa301c5f20664fc92e04501baf912b6d0d6989dfafa2e4e31b086b74e285d365ddf10e55386f113d985c1c4dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h3effdaca7d4e8970a1c1cdbfa8e24b4272c18048920de994298c8c12a10c80adb78dd058b4f0d031db529790a4d6292d6feb282faf620358e066adf455897c3581c2f0245b079c331d68b8efc602d08fc8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9dcac4f6f43409fc1fba49c2d02b6c556991bb37bbce34207f33b77279c9c4b7ca9ee1c346c4625cd548d1448a92f762b74a709887b2d471765cd4cb6b0cb95241a4e798de607696d0e76f8441e4e63ec0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h8659d78a67085fb9decf40c248a52c1e071017f6bac9f317ccc81f7de43cd867dbdcc147158c6c735c7dfdefc514d7312decf02d9dce9a874f0414e700d2e620203829b108ba061c9e0ac7e9f8cd0162fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hc61ca5d576a9da4f7715a68753f098b39ca109cfef843aa839ba17a3cf1ce0d07c7647a19b93fd0d2a1b5841ba4d35d488c8e9f9abb8e965fbe618d33576750a6af4eaa28bd13fb8c55c7240f079d624e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h899e507ff3f6c57a77111ed988c09a0bbc26ccdb5053c5f2fb2c139d6d09262fa136aa28eb431a38f0b9e7b6146da0f956da687d14ce7c58585174901202691487872e7cd2a0a01023657ffe354d8d9f5b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hb6d8526b4873ffb5c12db6ce4d49b055f2fdbdca838b3efdbc279236f414e2ec14c2bb49e7cffa35284fe0cf9994b2130a33db5b2284dc148e6385ab6a5b77e266d57ea38cfbba99ddc7d6d364f2016f79;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h45823052f1f30aad09ea9189be9f685d9f511ef2d7fa93e6cd1c1d7ad90bdd4fd5f83518b13f896071eeffee67bc117707b15840821f7900337f2476ccafc70e83f4289fde3e5f1fd05b1fcd831e63e1ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'ha1a7201a6d6316df2c6ead08332d3aff6c9d9f0989658c94da33efa8000ce4156018e8856c39ec6400965ecbfc743b7f55a01969a54ad0a42c8589a31b4e713ec23ee4ae118ee1ccea661447d22395e5a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h8c117e82ba781372c6c1f069b16a045f5dcb31d9af4737c9dbfbd4c47d7fea2a2108bb3b95340f27c00a02a224608117a7d3ae1b415d419e0d69ad3b791cccfc7fcb420127d938db56b4d5160c500c3e65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h43d4b92ff8451e4c3dd06708b91378406f96aa930e5fc684921a30f6ab8c893766ca5fdbc718b8d942541b55caa3f5abd3a27f5c94876379bff1bd1a14f41ffb14fb75c22dfd6756271bd4a281e1f29079;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hbb43c354f9d143d82bc984b5574b17540a91b7dbe62588a4610e3e9f47919c09341a9e2a060799966e56d30dee818b2326871c867322fbd51d71e14ab81e8665d3e0198e895399497b480cf488cbcd6e36;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h5bda3f13a2cc5e387d59fa4910f6e9dff0b486f0e3864bbe2bd0dee00db57e4ca6e6e46874177031035f66bf54404ee9cb33a3e172e0e1d06720653e4b624a6e779163ba73c68eece328ef31bc2675e6d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hccb1d43a4280a63187a1137cc7d00f177a274a1135d1f349c71812c04e4df53c9860acc26166e230988edbcbe0736ea332387b784e87266fb12ab6b534fa7f1af2018be1fc777e0a4c973c0a2e8d57d35a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h3baa49bf782a169671952c830a917dca776d615662339c1777ac663fc5df72adff4e2c9d016fc00135e4a72aa03a781b10069b5f690f483523d54d0c91ce9cb985a0acd1b46cd53aa471226901c981733a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hecfea114aeb685776d74308b01b37d198bc22493860ed8efa119af7a69a9ec1a12b1d634d0eafcd549896d5e6748e46b1323082b61ac5137da1d6290a07a200eb4caad20887f03671c766eea5894c83fc8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hba0f60b25a2a84010f0797fc2047c57c126db20c68fc6a97048fc8c7b7e72c4106c47ebca9c8179c63e1b7587be2f1f395bffce093ddf36bee6811b9ac1d6b8167030d1c4a1ad0c40304c4489db71a663a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h24c3d7898e30609636512f2877724ca38a14a2e1531625872d65790793b4abd870b71e3a7058c646d309936e951228d5ee6b718108fe3f162bcc2ee33369448cbd8c695e01ac2602319248f851244cc8a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h187cea8a3cdddf52d37efa6f8a758ceb7f4b8ba2ba7d9ccabb4a9e52f859e7cf015e6bf917d3d93ebe112adb032c24e3ed59811ea129f0270fb971f9a8df09b0d006d3b2bde8f382e18371029dab42d23b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h5f3c818655a6030e2d796f8e2abf32ffa5df558683c88d50600a3b2e7389f6ee47149c5750786c1bc8507527a82177737906dfcd246f66361c34463981f3381e359fedcb0a78e2f8401ed2666e81bb0d67;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h3e1d4990275c7445c1a384d23ef08b3da2d10276ad0b9e7378488f49c133cb420804343b1d6bbbdc69e48dd6270fac653d4ca718f5aa244bbee9af7bc15933a3824c0006487c1c80f0dffab2955968d88c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h9c33196b037a0edbeca15430473c70cd325c3c8ae126b24a7845bf5d5019fde9f48fb1fc232dd0b1556d1c771b2b9751488c49eb70396a454c93fd776258ae062dca5675f5ce6d8083dd60b7c4593068b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h3f557ff6e50fba9a0e0edd3f2c9c86c2210c481420cc3fe53f5a57d9a072df4738ddc45c6c4f7da690c1548bb2254967902847257777becee7bcb1ba440bad20a6bf7cfb27bcc201bf01c321c2e2825d87;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h4801f8220ee59a52664d719b3eaaaeb91277b035edf292fba7b27e4a9b4d8ca15e6284b542285fb25d1ea879f0363242129da8b2811566618f3095e2233b49f2943494bb7770d30d0660b4b92ae6015a7f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'ha0872b8b604f69079b1bcf152ec69c6cf470e79bb29ed3fe42aaf12df4e239197b94432f9b865d4c58fd1fb4d46939db72a6201340b41cb9bd625ec001ae18de3610666c18986d6a689e32ffe9ce9977ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hea0d351e439c688ebcb978d1b93f4ffd0d5bb1a42027c38e5a1773ba6081c8ccbc2c8e9a5f8b37012b54ab1f0752e16d948f502f6fb2a9d3a3805280877b3f2eec9663151c3f31579e6677a5c71e9f0a8d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h35eeaad6fcc413cffbf892b5f0b0763743aadc5421b347855ba709510a794dbde2a381d045ea37143c88151728bb3810b88a6493389c0ee86a894645538a34cdb46a7563ad1ecada8fd1049b0ee35579c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h6dc189b990704a2bb2c389f37b41ba2aadb408f1376e3cc7ec3eef62a3005a1c132156b2a3aae28ba280d5e4c8b247682c1c7c845ea055bd2f706b57463b8708c206ddf8fdc5197fce197ffffcbc6ffcb5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hbe76c389b63ebbc4f54dd2e3b63b707dda627c4ea255fc24e6a5b298fe704b6ddabfcf57ee998d5186d278d643935c1967b36e0cbe901a4a3b3fedabe3ead806df8628888d94e78ef45b9700550d85fb19;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h83dfa81d909d6883785bdf33a1e0816e9121071593b33751994931a93b8e3e16661913bdf057a4432a2cb7d7c046a61e1736384bd9fdd6af0308478ab86da377e8f0bebdbd7d592f1e672d910e1312885e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'hf8b8c423e8e4188210711d4a2180dc91f9509dc49abea5cae72ee3b69dc8c3a60c369f1ecc5b238ccd07b02773c39347cfab01607dc7d58f782a20438f3ed92cd44e04eb5957b9a410898736ae34c9c2cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h36cfeaaf9f4bfbeaf1519a1b275786648fcd3b576b58bab46169554737883069287719759c86c05262efd501746590adc8e517fc916612641551ae74db3b7db641a09da7fccb29cc10f87a6a1fec8ee989;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 648'h4f1e6773a1f2818bd77308613c06cf7826bd448d69c57ebbba4ceda1baba8759b395eb08be74ebd8537c1850a0f3bfff886aaeffb0143c402a64bc1292cfc5374839c4409ea963c65faeff4c352ce5ceea;
        #1
        $finish();
    end
endmodule
